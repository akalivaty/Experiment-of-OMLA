

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U554 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U555 ( .A1(n715), .A2(n951), .ZN(n721) );
  BUF_X1 U556 ( .A(n627), .Z(n628) );
  NOR2_X2 U557 ( .A1(G651), .A2(G543), .ZN(n671) );
  NAND2_X2 U558 ( .A1(n709), .A2(n814), .ZN(n758) );
  INV_X1 U559 ( .A(KEYINPUT105), .ZN(n780) );
  INV_X1 U560 ( .A(KEYINPUT17), .ZN(n525) );
  NOR2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  INV_X1 U562 ( .A(KEYINPUT23), .ZN(n527) );
  OR2_X1 U563 ( .A1(n741), .A2(n740), .ZN(n522) );
  OR2_X1 U564 ( .A1(n790), .A2(n777), .ZN(n523) );
  XOR2_X1 U565 ( .A(n748), .B(KEYINPUT31), .Z(n524) );
  INV_X1 U566 ( .A(KEYINPUT26), .ZN(n711) );
  INV_X1 U567 ( .A(KEYINPUT100), .ZN(n724) );
  INV_X1 U568 ( .A(KEYINPUT102), .ZN(n755) );
  NAND2_X1 U569 ( .A1(n930), .A2(n523), .ZN(n778) );
  XNOR2_X1 U570 ( .A(G543), .B(KEYINPUT0), .ZN(n555) );
  NAND2_X1 U571 ( .A1(G160), .A2(G40), .ZN(n813) );
  NOR2_X2 U572 ( .A1(G2104), .A2(n531), .ZN(n907) );
  XNOR2_X1 U573 ( .A(n528), .B(n527), .ZN(n529) );
  INV_X1 U574 ( .A(KEYINPUT72), .ZN(n569) );
  NAND2_X1 U575 ( .A1(n903), .A2(G138), .ZN(n541) );
  AND2_X1 U576 ( .A1(n541), .A2(n540), .ZN(G164) );
  XNOR2_X2 U577 ( .A(n526), .B(n525), .ZN(n903) );
  NAND2_X1 U578 ( .A1(n903), .A2(G137), .ZN(n530) );
  INV_X1 U579 ( .A(G2105), .ZN(n531) );
  AND2_X1 U580 ( .A1(n531), .A2(G2104), .ZN(n627) );
  NAND2_X1 U581 ( .A1(n627), .A2(G101), .ZN(n528) );
  NAND2_X1 U582 ( .A1(n530), .A2(n529), .ZN(n535) );
  NAND2_X1 U583 ( .A1(G125), .A2(n907), .ZN(n533) );
  AND2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n910) );
  NAND2_X1 U585 ( .A1(G113), .A2(n910), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X2 U587 ( .A1(n535), .A2(n534), .ZN(G160) );
  AND2_X1 U588 ( .A1(G102), .A2(n627), .ZN(n539) );
  NAND2_X1 U589 ( .A1(G126), .A2(n907), .ZN(n537) );
  NAND2_X1 U590 ( .A1(G114), .A2(n910), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U593 ( .A(G2451), .B(G2446), .ZN(n551) );
  XOR2_X1 U594 ( .A(G2430), .B(KEYINPUT109), .Z(n543) );
  XNOR2_X1 U595 ( .A(G2454), .B(G2435), .ZN(n542) );
  XNOR2_X1 U596 ( .A(n543), .B(n542), .ZN(n547) );
  XOR2_X1 U597 ( .A(G2438), .B(KEYINPUT108), .Z(n545) );
  XNOR2_X1 U598 ( .A(G1341), .B(G1348), .ZN(n544) );
  XNOR2_X1 U599 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U600 ( .A(n547), .B(n546), .Z(n549) );
  XNOR2_X1 U601 ( .A(G2443), .B(G2427), .ZN(n548) );
  XNOR2_X1 U602 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U603 ( .A(n551), .B(n550), .ZN(n552) );
  AND2_X1 U604 ( .A1(n552), .A2(G14), .ZN(G401) );
  AND2_X1 U605 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U606 ( .A(G860), .ZN(n615) );
  NAND2_X1 U607 ( .A1(G81), .A2(n671), .ZN(n553) );
  XNOR2_X1 U608 ( .A(n553), .B(KEYINPUT70), .ZN(n554) );
  XNOR2_X1 U609 ( .A(n554), .B(KEYINPUT12), .ZN(n559) );
  NAND2_X1 U610 ( .A1(n555), .A2(G651), .ZN(n556) );
  XNOR2_X1 U611 ( .A(n556), .B(KEYINPUT65), .ZN(n576) );
  NAND2_X1 U612 ( .A1(n576), .A2(G68), .ZN(n557) );
  XOR2_X1 U613 ( .A(n557), .B(KEYINPUT71), .Z(n558) );
  NAND2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U615 ( .A(n560), .B(KEYINPUT13), .ZN(n568) );
  XOR2_X1 U616 ( .A(G543), .B(KEYINPUT0), .Z(n665) );
  NOR2_X1 U617 ( .A1(n665), .A2(G651), .ZN(n561) );
  XNOR2_X2 U618 ( .A(n561), .B(KEYINPUT64), .ZN(n674) );
  AND2_X1 U619 ( .A1(G43), .A2(n674), .ZN(n566) );
  INV_X1 U620 ( .A(G651), .ZN(n562) );
  NOR2_X1 U621 ( .A1(G543), .A2(n562), .ZN(n563) );
  XOR2_X1 U622 ( .A(KEYINPUT1), .B(n563), .Z(n573) );
  NAND2_X1 U623 ( .A1(n573), .A2(G56), .ZN(n564) );
  XOR2_X1 U624 ( .A(KEYINPUT14), .B(n564), .Z(n565) );
  NOR2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n570) );
  XNOR2_X2 U627 ( .A(n570), .B(n569), .ZN(n951) );
  OR2_X1 U628 ( .A1(n615), .A2(n951), .ZN(G153) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  INV_X1 U631 ( .A(G120), .ZN(G236) );
  INV_X1 U632 ( .A(G69), .ZN(G235) );
  INV_X1 U633 ( .A(G108), .ZN(G238) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n571), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U636 ( .A(G223), .ZN(n847) );
  NAND2_X1 U637 ( .A1(n847), .A2(G567), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT11), .B(n572), .Z(G234) );
  BUF_X1 U639 ( .A(n573), .Z(n669) );
  NAND2_X1 U640 ( .A1(G64), .A2(n669), .ZN(n575) );
  NAND2_X1 U641 ( .A1(G52), .A2(n674), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n583) );
  NAND2_X1 U643 ( .A1(G90), .A2(n671), .ZN(n579) );
  INV_X1 U644 ( .A(n576), .ZN(n577) );
  INV_X1 U645 ( .A(n577), .ZN(n678) );
  NAND2_X1 U646 ( .A1(G77), .A2(n678), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U648 ( .A(KEYINPUT9), .B(n580), .Z(n581) );
  XNOR2_X1 U649 ( .A(KEYINPUT68), .B(n581), .ZN(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U651 ( .A(KEYINPUT69), .B(n584), .Z(G171) );
  INV_X1 U652 ( .A(G868), .ZN(n691) );
  NOR2_X1 U653 ( .A1(n691), .A2(G171), .ZN(n585) );
  XNOR2_X1 U654 ( .A(n585), .B(KEYINPUT73), .ZN(n595) );
  NAND2_X1 U655 ( .A1(n678), .A2(G79), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G54), .A2(n674), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U658 ( .A(KEYINPUT74), .B(n588), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G66), .A2(n669), .ZN(n590) );
  NAND2_X1 U660 ( .A1(G92), .A2(n671), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X2 U662 ( .A(KEYINPUT15), .B(n593), .Z(n938) );
  OR2_X1 U663 ( .A1(G868), .A2(n938), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U665 ( .A1(G63), .A2(n669), .ZN(n597) );
  NAND2_X1 U666 ( .A1(G51), .A2(n674), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U668 ( .A(KEYINPUT6), .B(n598), .ZN(n604) );
  NAND2_X1 U669 ( .A1(n671), .A2(G89), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n599), .B(KEYINPUT4), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G76), .A2(n678), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U673 ( .A(n602), .B(KEYINPUT5), .Z(n603) );
  NOR2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U675 ( .A(KEYINPUT7), .B(n605), .Z(n606) );
  XOR2_X1 U676 ( .A(KEYINPUT75), .B(n606), .Z(G168) );
  XOR2_X1 U677 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U678 ( .A1(G65), .A2(n669), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G53), .A2(n674), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G91), .A2(n671), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G78), .A2(n678), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n933) );
  INV_X1 U685 ( .A(n933), .ZN(G299) );
  NOR2_X1 U686 ( .A1(G286), .A2(n691), .ZN(n614) );
  NOR2_X1 U687 ( .A1(G868), .A2(G299), .ZN(n613) );
  NOR2_X1 U688 ( .A1(n614), .A2(n613), .ZN(G297) );
  NAND2_X1 U689 ( .A1(n615), .A2(G559), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n616), .A2(n938), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n617), .B(KEYINPUT76), .ZN(n618) );
  XNOR2_X1 U692 ( .A(KEYINPUT16), .B(n618), .ZN(G148) );
  NAND2_X1 U693 ( .A1(n938), .A2(G868), .ZN(n619) );
  XOR2_X1 U694 ( .A(KEYINPUT77), .B(n619), .Z(n620) );
  NOR2_X1 U695 ( .A1(G559), .A2(n620), .ZN(n622) );
  NOR2_X1 U696 ( .A1(n951), .A2(G868), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U698 ( .A1(n907), .A2(G123), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT18), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G135), .A2(n903), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U702 ( .A(KEYINPUT78), .B(n626), .ZN(n632) );
  NAND2_X1 U703 ( .A1(G99), .A2(n628), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G111), .A2(n910), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U707 ( .A(KEYINPUT79), .B(n633), .Z(n992) );
  XNOR2_X1 U708 ( .A(n992), .B(G2096), .ZN(n635) );
  INV_X1 U709 ( .A(G2100), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(G156) );
  NAND2_X1 U711 ( .A1(G559), .A2(n938), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n636), .B(n951), .ZN(n688) );
  NOR2_X1 U713 ( .A1(G860), .A2(n688), .ZN(n644) );
  NAND2_X1 U714 ( .A1(G93), .A2(n671), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G80), .A2(n678), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U717 ( .A(KEYINPUT80), .B(n639), .ZN(n643) );
  NAND2_X1 U718 ( .A1(G67), .A2(n669), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G55), .A2(n674), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  OR2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n690) );
  XOR2_X1 U722 ( .A(n644), .B(n690), .Z(G145) );
  NAND2_X1 U723 ( .A1(n671), .A2(G86), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n645), .B(KEYINPUT82), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G61), .A2(n669), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U727 ( .A1(G73), .A2(n678), .ZN(n648) );
  XNOR2_X1 U728 ( .A(n648), .B(KEYINPUT83), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n649), .B(KEYINPUT2), .ZN(n650) );
  NOR2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n652), .B(KEYINPUT84), .ZN(n654) );
  NAND2_X1 U732 ( .A1(G48), .A2(n674), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U734 ( .A(KEYINPUT85), .B(n655), .Z(G305) );
  NAND2_X1 U735 ( .A1(G88), .A2(n671), .ZN(n657) );
  NAND2_X1 U736 ( .A1(G75), .A2(n678), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n661) );
  NAND2_X1 U738 ( .A1(G62), .A2(n669), .ZN(n659) );
  NAND2_X1 U739 ( .A1(G50), .A2(n674), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U741 ( .A1(n661), .A2(n660), .ZN(G166) );
  NAND2_X1 U742 ( .A1(G651), .A2(G74), .ZN(n663) );
  NAND2_X1 U743 ( .A1(G49), .A2(n674), .ZN(n662) );
  NAND2_X1 U744 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U745 ( .A1(n669), .A2(n664), .ZN(n668) );
  NAND2_X1 U746 ( .A1(G87), .A2(n665), .ZN(n666) );
  XOR2_X1 U747 ( .A(KEYINPUT81), .B(n666), .Z(n667) );
  NAND2_X1 U748 ( .A1(n668), .A2(n667), .ZN(G288) );
  NAND2_X1 U749 ( .A1(n669), .A2(G60), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n670), .B(KEYINPUT66), .ZN(n673) );
  NAND2_X1 U751 ( .A1(G85), .A2(n671), .ZN(n672) );
  NAND2_X1 U752 ( .A1(n673), .A2(n672), .ZN(n677) );
  NAND2_X1 U753 ( .A1(G47), .A2(n674), .ZN(n675) );
  XNOR2_X1 U754 ( .A(KEYINPUT67), .B(n675), .ZN(n676) );
  NOR2_X1 U755 ( .A1(n677), .A2(n676), .ZN(n680) );
  NAND2_X1 U756 ( .A1(n678), .A2(G72), .ZN(n679) );
  NAND2_X1 U757 ( .A1(n680), .A2(n679), .ZN(G290) );
  XNOR2_X1 U758 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n682) );
  XNOR2_X1 U759 ( .A(G288), .B(KEYINPUT19), .ZN(n681) );
  XNOR2_X1 U760 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U761 ( .A(G166), .B(n683), .ZN(n685) );
  XNOR2_X1 U762 ( .A(G290), .B(n933), .ZN(n684) );
  XNOR2_X1 U763 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U764 ( .A(n690), .B(n686), .ZN(n687) );
  XNOR2_X1 U765 ( .A(G305), .B(n687), .ZN(n855) );
  XNOR2_X1 U766 ( .A(n688), .B(n855), .ZN(n689) );
  NAND2_X1 U767 ( .A1(n689), .A2(G868), .ZN(n693) );
  NAND2_X1 U768 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U769 ( .A1(n693), .A2(n692), .ZN(G295) );
  NAND2_X1 U770 ( .A1(G2084), .A2(G2078), .ZN(n694) );
  XOR2_X1 U771 ( .A(KEYINPUT20), .B(n694), .Z(n695) );
  NAND2_X1 U772 ( .A1(G2090), .A2(n695), .ZN(n696) );
  XNOR2_X1 U773 ( .A(KEYINPUT21), .B(n696), .ZN(n697) );
  NAND2_X1 U774 ( .A1(n697), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U775 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U776 ( .A1(G235), .A2(G236), .ZN(n698) );
  XNOR2_X1 U777 ( .A(n698), .B(KEYINPUT89), .ZN(n699) );
  NOR2_X1 U778 ( .A1(G238), .A2(n699), .ZN(n700) );
  NAND2_X1 U779 ( .A1(G57), .A2(n700), .ZN(n853) );
  NAND2_X1 U780 ( .A1(n853), .A2(G567), .ZN(n706) );
  NOR2_X1 U781 ( .A1(G220), .A2(G219), .ZN(n701) );
  XNOR2_X1 U782 ( .A(KEYINPUT22), .B(n701), .ZN(n702) );
  NAND2_X1 U783 ( .A1(n702), .A2(G96), .ZN(n703) );
  NOR2_X1 U784 ( .A1(G218), .A2(n703), .ZN(n704) );
  XOR2_X1 U785 ( .A(KEYINPUT88), .B(n704), .Z(n854) );
  NAND2_X1 U786 ( .A1(n854), .A2(G2106), .ZN(n705) );
  NAND2_X1 U787 ( .A1(n706), .A2(n705), .ZN(n929) );
  NAND2_X1 U788 ( .A1(G483), .A2(G661), .ZN(n707) );
  NOR2_X1 U789 ( .A1(n929), .A2(n707), .ZN(n850) );
  NAND2_X1 U790 ( .A1(n850), .A2(G36), .ZN(G176) );
  INV_X1 U791 ( .A(G171), .ZN(G301) );
  XOR2_X1 U792 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  INV_X1 U793 ( .A(n813), .ZN(n709) );
  NOR2_X2 U794 ( .A1(G164), .A2(G1384), .ZN(n814) );
  INV_X1 U795 ( .A(n758), .ZN(n710) );
  AND2_X1 U796 ( .A1(n710), .A2(G1996), .ZN(n712) );
  XNOR2_X1 U797 ( .A(n712), .B(n711), .ZN(n714) );
  NAND2_X1 U798 ( .A1(n758), .A2(G1341), .ZN(n713) );
  NAND2_X1 U799 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U800 ( .A1(n721), .A2(n938), .ZN(n719) );
  INV_X1 U801 ( .A(n758), .ZN(n737) );
  NOR2_X1 U802 ( .A1(n737), .A2(G1348), .ZN(n717) );
  NOR2_X1 U803 ( .A1(G2067), .A2(n758), .ZN(n716) );
  NOR2_X1 U804 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U805 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U806 ( .A(n720), .B(KEYINPUT99), .ZN(n723) );
  NOR2_X1 U807 ( .A1(n938), .A2(n721), .ZN(n722) );
  NOR2_X1 U808 ( .A1(n723), .A2(n722), .ZN(n725) );
  XNOR2_X1 U809 ( .A(n725), .B(n724), .ZN(n731) );
  NAND2_X1 U810 ( .A1(G2072), .A2(n737), .ZN(n726) );
  XNOR2_X1 U811 ( .A(n726), .B(KEYINPUT98), .ZN(n727) );
  XNOR2_X1 U812 ( .A(KEYINPUT27), .B(n727), .ZN(n729) );
  INV_X1 U813 ( .A(G1956), .ZN(n959) );
  NOR2_X1 U814 ( .A1(n737), .A2(n959), .ZN(n728) );
  NOR2_X1 U815 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U816 ( .A1(n732), .A2(n933), .ZN(n730) );
  NAND2_X1 U817 ( .A1(n731), .A2(n730), .ZN(n735) );
  NOR2_X1 U818 ( .A1(n732), .A2(n933), .ZN(n733) );
  XOR2_X1 U819 ( .A(n733), .B(KEYINPUT28), .Z(n734) );
  NAND2_X1 U820 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U821 ( .A(n736), .B(KEYINPUT29), .ZN(n741) );
  XOR2_X1 U822 ( .A(G2078), .B(KEYINPUT25), .Z(n1020) );
  NOR2_X1 U823 ( .A1(n1020), .A2(n758), .ZN(n739) );
  NOR2_X1 U824 ( .A1(n737), .A2(G1961), .ZN(n738) );
  NOR2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n745) );
  NOR2_X1 U826 ( .A1(G301), .A2(n745), .ZN(n740) );
  NAND2_X1 U827 ( .A1(G8), .A2(n758), .ZN(n790) );
  NOR2_X1 U828 ( .A1(G1966), .A2(n790), .ZN(n750) );
  NOR2_X1 U829 ( .A1(G2084), .A2(n758), .ZN(n749) );
  NOR2_X1 U830 ( .A1(n750), .A2(n749), .ZN(n742) );
  NAND2_X1 U831 ( .A1(G8), .A2(n742), .ZN(n743) );
  XNOR2_X1 U832 ( .A(KEYINPUT30), .B(n743), .ZN(n744) );
  NOR2_X1 U833 ( .A1(G168), .A2(n744), .ZN(n747) );
  AND2_X1 U834 ( .A1(G301), .A2(n745), .ZN(n746) );
  NOR2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n522), .A2(n524), .ZN(n757) );
  XNOR2_X1 U837 ( .A(n757), .B(KEYINPUT101), .ZN(n754) );
  NAND2_X1 U838 ( .A1(n749), .A2(G8), .ZN(n752) );
  INV_X1 U839 ( .A(n750), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n756) );
  XNOR2_X1 U842 ( .A(n756), .B(n755), .ZN(n768) );
  NAND2_X1 U843 ( .A1(n757), .A2(G286), .ZN(n764) );
  NOR2_X1 U844 ( .A1(G1971), .A2(n790), .ZN(n760) );
  NOR2_X1 U845 ( .A1(G2090), .A2(n758), .ZN(n759) );
  NOR2_X1 U846 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U847 ( .A1(G303), .A2(n761), .ZN(n762) );
  XOR2_X1 U848 ( .A(KEYINPUT103), .B(n762), .Z(n763) );
  NAND2_X1 U849 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U850 ( .A1(n765), .A2(G8), .ZN(n766) );
  XNOR2_X1 U851 ( .A(KEYINPUT32), .B(n766), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n768), .A2(n767), .ZN(n787) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n945) );
  NOR2_X1 U854 ( .A1(G303), .A2(G1971), .ZN(n935) );
  NOR2_X1 U855 ( .A1(n945), .A2(n935), .ZN(n770) );
  INV_X1 U856 ( .A(KEYINPUT33), .ZN(n769) );
  AND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n787), .A2(n771), .ZN(n775) );
  INV_X1 U859 ( .A(n790), .ZN(n772) );
  NAND2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n944) );
  AND2_X1 U861 ( .A1(n772), .A2(n944), .ZN(n773) );
  OR2_X1 U862 ( .A1(KEYINPUT33), .A2(n773), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U864 ( .A(n776), .B(KEYINPUT104), .ZN(n779) );
  XOR2_X1 U865 ( .A(G1981), .B(G305), .Z(n930) );
  NAND2_X1 U866 ( .A1(n945), .A2(KEYINPUT33), .ZN(n777) );
  NOR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n781) );
  XNOR2_X1 U868 ( .A(n781), .B(n780), .ZN(n786) );
  NOR2_X1 U869 ( .A1(G1981), .A2(G305), .ZN(n782) );
  XNOR2_X1 U870 ( .A(n782), .B(KEYINPUT24), .ZN(n783) );
  XNOR2_X1 U871 ( .A(n783), .B(KEYINPUT97), .ZN(n784) );
  NOR2_X1 U872 ( .A1(n790), .A2(n784), .ZN(n785) );
  NOR2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n793) );
  NOR2_X1 U874 ( .A1(G2090), .A2(G303), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G8), .A2(n788), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n787), .A2(n789), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U878 ( .A1(n793), .A2(n792), .ZN(n830) );
  NAND2_X1 U879 ( .A1(G141), .A2(n903), .ZN(n795) );
  NAND2_X1 U880 ( .A1(G129), .A2(n907), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n798) );
  NAND2_X1 U882 ( .A1(n628), .A2(G105), .ZN(n796) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(n796), .Z(n797) );
  NOR2_X1 U884 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n910), .A2(G117), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n888) );
  NAND2_X1 U887 ( .A1(G1996), .A2(n888), .ZN(n801) );
  XOR2_X1 U888 ( .A(KEYINPUT95), .B(n801), .Z(n812) );
  NAND2_X1 U889 ( .A1(n907), .A2(G119), .ZN(n802) );
  XNOR2_X1 U890 ( .A(n802), .B(KEYINPUT92), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G107), .A2(n910), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U893 ( .A(KEYINPUT93), .B(n805), .ZN(n810) );
  NAND2_X1 U894 ( .A1(G131), .A2(n903), .ZN(n807) );
  NAND2_X1 U895 ( .A1(G95), .A2(n628), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U897 ( .A(KEYINPUT94), .B(n808), .Z(n809) );
  NAND2_X1 U898 ( .A1(n810), .A2(n809), .ZN(n889) );
  NAND2_X1 U899 ( .A1(G1991), .A2(n889), .ZN(n811) );
  NAND2_X1 U900 ( .A1(n812), .A2(n811), .ZN(n991) );
  NOR2_X1 U901 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U902 ( .A(KEYINPUT91), .B(n815), .Z(n842) );
  NAND2_X1 U903 ( .A1(n991), .A2(n842), .ZN(n816) );
  XOR2_X1 U904 ( .A(KEYINPUT96), .B(n816), .Z(n834) );
  INV_X1 U905 ( .A(n842), .ZN(n827) );
  NAND2_X1 U906 ( .A1(G140), .A2(n903), .ZN(n818) );
  NAND2_X1 U907 ( .A1(G104), .A2(n628), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U909 ( .A(KEYINPUT34), .B(n819), .ZN(n824) );
  NAND2_X1 U910 ( .A1(G128), .A2(n907), .ZN(n821) );
  NAND2_X1 U911 ( .A1(G116), .A2(n910), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n822) );
  XOR2_X1 U913 ( .A(KEYINPUT35), .B(n822), .Z(n823) );
  NOR2_X1 U914 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U915 ( .A(KEYINPUT36), .B(n825), .ZN(n921) );
  XNOR2_X1 U916 ( .A(G2067), .B(KEYINPUT37), .ZN(n839) );
  NOR2_X1 U917 ( .A1(n921), .A2(n839), .ZN(n837) );
  XNOR2_X1 U918 ( .A(G1986), .B(G290), .ZN(n934) );
  NOR2_X1 U919 ( .A1(n837), .A2(n934), .ZN(n826) );
  NOR2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U921 ( .A1(n834), .A2(n828), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U923 ( .A(n831), .B(KEYINPUT106), .ZN(n844) );
  NOR2_X1 U924 ( .A1(G1996), .A2(n888), .ZN(n998) );
  NOR2_X1 U925 ( .A1(G1986), .A2(G290), .ZN(n832) );
  NOR2_X1 U926 ( .A1(G1991), .A2(n889), .ZN(n1002) );
  NOR2_X1 U927 ( .A1(n832), .A2(n1002), .ZN(n833) );
  NOR2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n835) );
  NOR2_X1 U929 ( .A1(n998), .A2(n835), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n836), .B(KEYINPUT39), .ZN(n838) );
  INV_X1 U931 ( .A(n837), .ZN(n985) );
  NAND2_X1 U932 ( .A1(n838), .A2(n985), .ZN(n840) );
  NAND2_X1 U933 ( .A1(n921), .A2(n839), .ZN(n986) );
  NAND2_X1 U934 ( .A1(n840), .A2(n986), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n842), .A2(n841), .ZN(n843) );
  NAND2_X1 U936 ( .A1(n844), .A2(n843), .ZN(n846) );
  XOR2_X1 U937 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n845) );
  XNOR2_X1 U938 ( .A(n846), .B(n845), .ZN(G329) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n847), .ZN(G217) );
  NAND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n848) );
  XOR2_X1 U941 ( .A(KEYINPUT110), .B(n848), .Z(n849) );
  NAND2_X1 U942 ( .A1(G661), .A2(n849), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n851) );
  NAND2_X1 U944 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U945 ( .A(KEYINPUT111), .B(n852), .Z(G188) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  NOR2_X1 U948 ( .A1(n854), .A2(n853), .ZN(G325) );
  INV_X1 U949 ( .A(G325), .ZN(G261) );
  XOR2_X1 U950 ( .A(n855), .B(G286), .Z(n857) );
  XNOR2_X1 U951 ( .A(G171), .B(n938), .ZN(n856) );
  XNOR2_X1 U952 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U953 ( .A(n858), .B(n951), .ZN(n859) );
  NOR2_X1 U954 ( .A1(G37), .A2(n859), .ZN(G397) );
  XNOR2_X1 U955 ( .A(G1991), .B(KEYINPUT41), .ZN(n869) );
  XOR2_X1 U956 ( .A(G1956), .B(G1961), .Z(n861) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1986), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U959 ( .A(G1976), .B(G1981), .Z(n863) );
  XNOR2_X1 U960 ( .A(G1966), .B(G1971), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U962 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U963 ( .A(KEYINPUT114), .B(G2474), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n869), .B(n868), .ZN(G229) );
  XOR2_X1 U966 ( .A(KEYINPUT43), .B(G2678), .Z(n871) );
  XNOR2_X1 U967 ( .A(KEYINPUT113), .B(KEYINPUT112), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U969 ( .A(KEYINPUT42), .B(G2090), .Z(n873) );
  XNOR2_X1 U970 ( .A(G2067), .B(G2072), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U972 ( .A(n875), .B(n874), .Z(n877) );
  XNOR2_X1 U973 ( .A(G2096), .B(G2100), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n879) );
  XOR2_X1 U975 ( .A(G2084), .B(G2078), .Z(n878) );
  XNOR2_X1 U976 ( .A(n879), .B(n878), .ZN(G227) );
  NAND2_X1 U977 ( .A1(G124), .A2(n907), .ZN(n880) );
  XOR2_X1 U978 ( .A(KEYINPUT44), .B(n880), .Z(n881) );
  XNOR2_X1 U979 ( .A(n881), .B(KEYINPUT115), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G112), .A2(n910), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G136), .A2(n903), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G100), .A2(n628), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n886) );
  NOR2_X1 U985 ( .A1(n887), .A2(n886), .ZN(G162) );
  XNOR2_X1 U986 ( .A(G162), .B(n888), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n894) );
  XOR2_X1 U988 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n892) );
  XNOR2_X1 U989 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U991 ( .A(n894), .B(n893), .Z(n918) );
  NAND2_X1 U992 ( .A1(G139), .A2(n903), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G103), .A2(n628), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n902) );
  NAND2_X1 U995 ( .A1(G127), .A2(n907), .ZN(n898) );
  NAND2_X1 U996 ( .A1(G115), .A2(n910), .ZN(n897) );
  NAND2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U998 ( .A(KEYINPUT47), .B(n899), .ZN(n900) );
  XNOR2_X1 U999 ( .A(KEYINPUT117), .B(n900), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n987) );
  XNOR2_X1 U1001 ( .A(G160), .B(n987), .ZN(n915) );
  NAND2_X1 U1002 ( .A1(G142), .A2(n903), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(G106), .A2(n628), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n906), .B(KEYINPUT45), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(G130), .A2(n907), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(n910), .A2(G118), .ZN(n911) );
  XOR2_X1 U1009 ( .A(KEYINPUT116), .B(n911), .Z(n912) );
  NOR2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(G164), .B(n916), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1014 ( .A(n992), .B(n919), .Z(n920) );
  XNOR2_X1 U1015 ( .A(n921), .B(n920), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n922), .ZN(G395) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n929), .ZN(n926) );
  NOR2_X1 U1018 ( .A1(G229), .A2(G227), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n923), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G397), .A2(n924), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(n927), .A2(G395), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(n928), .B(KEYINPUT120), .ZN(G308) );
  INV_X1 U1024 ( .A(G308), .ZN(G225) );
  INV_X1 U1025 ( .A(n929), .ZN(G319) );
  INV_X1 U1026 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1027 ( .A(G16), .B(KEYINPUT56), .ZN(n957) );
  XNOR2_X1 U1028 ( .A(G1966), .B(G168), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(KEYINPUT57), .B(n932), .ZN(n955) );
  XNOR2_X1 U1031 ( .A(n933), .B(G1956), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(n938), .B(G1348), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G171), .B(G1961), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n949) );
  NAND2_X1 U1038 ( .A1(G303), .A2(G1971), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n947) );
  XOR2_X1 U1040 ( .A(n945), .B(KEYINPUT123), .Z(n946) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(n950), .B(KEYINPUT124), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(n951), .B(G1341), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1047 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1048 ( .A(n958), .B(KEYINPUT125), .ZN(n984) );
  XNOR2_X1 U1049 ( .A(G20), .B(n959), .ZN(n963) );
  XNOR2_X1 U1050 ( .A(G1341), .B(G19), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G6), .B(G1981), .ZN(n960) );
  NOR2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1054 ( .A(KEYINPUT59), .B(G1348), .Z(n964) );
  XNOR2_X1 U1055 ( .A(G4), .B(n964), .ZN(n965) );
  NOR2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(KEYINPUT126), .B(n967), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(n968), .B(KEYINPUT60), .ZN(n972) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G21), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(G1961), .B(G5), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n980) );
  XNOR2_X1 U1063 ( .A(G1986), .B(G24), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(G1971), .B(G22), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(G1976), .B(KEYINPUT127), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n975), .B(G23), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(KEYINPUT58), .B(n978), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1071 ( .A(KEYINPUT61), .B(n981), .Z(n982) );
  NOR2_X1 U1072 ( .A1(G16), .A2(n982), .ZN(n983) );
  NOR2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n1011) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n996) );
  XOR2_X1 U1075 ( .A(G2072), .B(n987), .Z(n989) );
  XOR2_X1 U1076 ( .A(G164), .B(G2078), .Z(n988) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(KEYINPUT50), .B(n990), .ZN(n994) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1081 ( .A1(n996), .A2(n995), .ZN(n1005) );
  XNOR2_X1 U1082 ( .A(G160), .B(G2084), .ZN(n1001) );
  XOR2_X1 U1083 ( .A(G2090), .B(G162), .Z(n997) );
  NOR2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1085 ( .A(KEYINPUT51), .B(n999), .Z(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  NOR2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1088 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(KEYINPUT52), .B(n1006), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(KEYINPUT121), .B(n1007), .ZN(n1008) );
  INV_X1 U1091 ( .A(KEYINPUT55), .ZN(n1030) );
  NAND2_X1 U1092 ( .A1(n1008), .A2(n1030), .ZN(n1009) );
  NAND2_X1 U1093 ( .A1(n1009), .A2(G29), .ZN(n1010) );
  NAND2_X1 U1094 ( .A1(n1011), .A2(n1010), .ZN(n1035) );
  XNOR2_X1 U1095 ( .A(G2090), .B(G35), .ZN(n1025) );
  XNOR2_X1 U1096 ( .A(G1996), .B(G32), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G33), .B(G2072), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1019) );
  XOR2_X1 U1099 ( .A(G2067), .B(G26), .Z(n1014) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(G28), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(G25), .B(G1991), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(KEYINPUT122), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(G27), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(KEYINPUT53), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1028) );
  XOR2_X1 U1109 ( .A(G2084), .B(G34), .Z(n1026) );
  XNOR2_X1 U1110 ( .A(KEYINPUT54), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(n1030), .B(n1029), .ZN(n1032) );
  INV_X1 U1113 ( .A(G29), .ZN(n1031) );
  NAND2_X1 U1114 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1115 ( .A1(G11), .A2(n1033), .ZN(n1034) );
  NOR2_X1 U1116 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1117 ( .A(n1036), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

