//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959;
  NAND2_X1  g000(.A1(G211gat), .A2(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT72), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(KEYINPUT72), .A3(new_n208), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(KEYINPUT22), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n205), .A2(new_n202), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G226gat), .ZN(new_n215));
  INV_X1    g014(.A(G233gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  AND2_X1   g019(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT67), .B1(new_n223), .B2(KEYINPUT66), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT28), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n219), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT27), .B(G183gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(new_n220), .ZN(new_n230));
  OAI211_X1 g029(.A(KEYINPUT28), .B(new_n227), .C1(new_n230), .C2(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT26), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT68), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n234), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n238), .B(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n226), .A2(new_n231), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n218), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(G183gat), .A2(G190gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n242), .B1(new_n219), .B2(KEYINPUT65), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n218), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n245), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n233), .A2(KEYINPUT23), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT23), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(G169gat), .B2(G176gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n252), .A3(new_n232), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n249), .A2(KEYINPUT25), .A3(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n243), .A2(new_n257), .A3(new_n244), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n258), .B2(new_n253), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT29), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n217), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n217), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n241), .B2(new_n260), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n214), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n217), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n212), .A2(new_n202), .A3(new_n205), .ZN(new_n268));
  INV_X1    g067(.A(new_n211), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n268), .B1(new_n269), .B2(new_n209), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT29), .B1(new_n241), .B2(new_n260), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n267), .B(new_n270), .C1(new_n217), .C2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G64gat), .B(G92gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n266), .A2(KEYINPUT30), .A3(new_n272), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n266), .A2(new_n272), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n275), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n266), .A2(new_n276), .A3(new_n272), .ZN(new_n280));
  XOR2_X1   g079(.A(KEYINPUT73), .B(KEYINPUT30), .Z(new_n281));
  AND3_X1   g080(.A1(new_n280), .A2(KEYINPUT74), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT74), .B1(new_n280), .B2(new_n281), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n277), .B(new_n279), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G113gat), .ZN(new_n287));
  INV_X1    g086(.A(G113gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G120gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n291));
  INV_X1    g090(.A(G134gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G127gat), .ZN(new_n293));
  INV_X1    g092(.A(G127gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G134gat), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n290), .A2(new_n291), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n295), .ZN(new_n297));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n297), .B1(new_n298), .B2(KEYINPUT1), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G141gat), .B(G148gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n305), .B1(G155gat), .B2(G162gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G141gat), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G148gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G155gat), .B(G162gat), .ZN(new_n313));
  INV_X1    g112(.A(G155gat), .ZN(new_n314));
  INV_X1    g113(.A(G162gat), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT2), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n318), .A3(KEYINPUT4), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n296), .A2(new_n299), .A3(new_n307), .A4(new_n317), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT76), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n317), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n296), .A2(new_n299), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n307), .A2(new_n317), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  OR3_X1    g129(.A1(new_n320), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n331));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(KEYINPUT5), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n324), .A2(new_n330), .A3(new_n331), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n333), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n330), .A2(new_n319), .A3(new_n322), .A4(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n327), .A2(new_n325), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n320), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n340), .B2(new_n333), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n337), .A2(new_n341), .A3(KEYINPUT75), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT75), .B1(new_n337), .B2(new_n341), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n335), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(G85gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT0), .B(G57gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n346), .B(new_n347), .Z(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT6), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n335), .B(new_n348), .C1(new_n342), .C2(new_n343), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT77), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n344), .A2(KEYINPUT6), .A3(new_n349), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n350), .A2(new_n356), .A3(new_n351), .A4(new_n352), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n285), .A2(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n241), .A2(new_n300), .A3(new_n260), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n300), .B1(new_n241), .B2(new_n260), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G227gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(new_n216), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT33), .ZN(new_n369));
  XNOR2_X1  g168(.A(G15gat), .B(G43gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(G99gat), .ZN(new_n371));
  XOR2_X1   g170(.A(KEYINPUT69), .B(G71gat), .Z(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT70), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n369), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n374), .B2(new_n373), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n364), .B1(new_n360), .B2(new_n361), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT32), .ZN(new_n378));
  INV_X1    g177(.A(new_n373), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n261), .A2(new_n327), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n241), .A2(new_n300), .A3(new_n260), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n365), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT32), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n382), .A2(KEYINPUT33), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n368), .B(new_n378), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n377), .A2(KEYINPUT32), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n377), .A2(new_n369), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n379), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n368), .B1(new_n390), .B2(new_n378), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n366), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT31), .B(G50gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(G78gat), .B(G106gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n328), .B1(new_n214), .B2(KEYINPUT29), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n325), .ZN(new_n398));
  INV_X1    g197(.A(G22gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT78), .ZN(new_n400));
  INV_X1    g199(.A(G228gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n401), .B2(new_n216), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n329), .A2(new_n262), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n214), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n398), .A2(new_n399), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT3), .B1(new_n270), .B2(new_n262), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n402), .B(new_n404), .C1(new_n406), .C2(new_n318), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(G22gat), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n400), .A2(new_n401), .A3(new_n216), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n405), .B2(new_n408), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n396), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n405), .A2(new_n408), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n409), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(new_n411), .A3(new_n395), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n378), .B1(new_n384), .B2(new_n385), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n367), .ZN(new_n420));
  INV_X1    g219(.A(new_n366), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n386), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n392), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT35), .B1(new_n359), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT82), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n426), .B(KEYINPUT35), .C1(new_n359), .C2(new_n423), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n423), .A2(new_n284), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n353), .A2(new_n355), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(KEYINPUT35), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n324), .A2(new_n330), .A3(new_n331), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n333), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n333), .B2(new_n340), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT39), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT40), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n348), .B1(new_n435), .B2(KEYINPUT39), .ZN(new_n440));
  OR3_X1    g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n438), .B2(new_n440), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n441), .A2(new_n284), .A3(new_n350), .A4(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT37), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n266), .A2(new_n444), .A3(new_n272), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT79), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n266), .A2(KEYINPUT79), .A3(new_n272), .A4(new_n444), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n444), .B1(new_n266), .B2(new_n272), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n450), .A2(KEYINPUT38), .A3(new_n276), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT80), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n449), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n453), .A2(new_n280), .A3(new_n430), .A4(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT38), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n450), .A2(new_n276), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n458), .A2(KEYINPUT81), .B1(new_n447), .B2(new_n448), .ZN(new_n459));
  OR3_X1    g258(.A1(new_n450), .A2(KEYINPUT81), .A3(new_n276), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n418), .B(new_n443), .C1(new_n456), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n387), .A2(new_n391), .A3(new_n366), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n421), .B1(new_n420), .B2(new_n386), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n392), .A2(KEYINPUT36), .A3(new_n422), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n418), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n359), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n462), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n433), .A2(new_n471), .A3(KEYINPUT83), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT83), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n425), .A2(new_n427), .B1(new_n431), .B2(new_n429), .ZN(new_n474));
  INV_X1    g273(.A(new_n471), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n477));
  XOR2_X1   g276(.A(G15gat), .B(G22gat), .Z(new_n478));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G15gat), .B(G22gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT85), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT16), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(G1gat), .ZN(new_n485));
  INV_X1    g284(.A(G1gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n486), .A3(new_n482), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n480), .A2(new_n482), .B1(KEYINPUT16), .B2(new_n486), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n490));
  OAI21_X1  g289(.A(G8gat), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n488), .B(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT14), .ZN(new_n493));
  INV_X1    g292(.A(G29gat), .ZN(new_n494));
  INV_X1    g293(.A(G36gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n496), .A2(new_n497), .B1(G29gat), .B2(G36gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT15), .ZN(new_n499));
  XOR2_X1   g298(.A(G43gat), .B(G50gat), .Z(new_n500));
  OR3_X1    g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n499), .ZN(new_n502));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n504), .A3(new_n498), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n477), .B1(new_n492), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n501), .A2(KEYINPUT17), .A3(new_n505), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n506), .B2(KEYINPUT17), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n501), .A2(new_n505), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(KEYINPUT84), .A3(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n492), .A2(new_n510), .A3(new_n512), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n507), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n512), .A2(new_n515), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(new_n477), .A3(new_n510), .A4(new_n492), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT18), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n517), .A2(KEYINPUT89), .A3(new_n518), .A4(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n517), .A2(KEYINPUT18), .A3(new_n518), .A4(new_n520), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n492), .B(new_n506), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n518), .B(KEYINPUT13), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G113gat), .B(G141gat), .Z(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G197gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT11), .B(G169gat), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n534), .B(new_n535), .Z(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT12), .Z(new_n537));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n531), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n532), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n526), .A2(new_n530), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(new_n523), .B2(new_n524), .ZN(new_n542));
  INV_X1    g341(.A(new_n537), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n541), .B2(KEYINPUT90), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G230gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(new_n216), .ZN(new_n548));
  NAND2_X1  g347(.A1(G85gat), .A2(G92gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT7), .ZN(new_n550));
  INV_X1    g349(.A(G99gat), .ZN(new_n551));
  INV_X1    g350(.A(G106gat), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT8), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n550), .B(new_n553), .C1(G85gat), .C2(G92gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(G99gat), .B(G106gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G57gat), .B(G64gat), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n558));
  XOR2_X1   g357(.A(G71gat), .B(G78gat), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n559), .A2(KEYINPUT91), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  INV_X1    g362(.A(G78gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(KEYINPUT91), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n561), .A2(new_n557), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n556), .A2(new_n560), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT10), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n554), .B(new_n555), .Z(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n560), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(new_n569), .A3(new_n568), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n548), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  AOI211_X1 g374(.A(new_n547), .B(new_n216), .C1(new_n573), .C2(new_n568), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G120gat), .B(G148gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  OR3_X1    g380(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT97), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT97), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n577), .A2(new_n584), .A3(new_n580), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n546), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n472), .A2(new_n476), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT21), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n492), .B1(new_n589), .B2(new_n572), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(G183gat), .ZN(new_n591));
  AND2_X1   g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G211gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n572), .A2(new_n589), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT92), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n597), .A2(new_n603), .A3(new_n598), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n510), .A2(new_n512), .A3(new_n571), .A4(new_n515), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n519), .A2(KEYINPUT93), .A3(new_n571), .A4(new_n510), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n556), .A2(new_n513), .ZN(new_n615));
  NAND3_X1  g414(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT94), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n619), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n610), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n617), .A2(KEYINPUT95), .A3(new_n619), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n624), .A2(new_n620), .A3(new_n610), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT96), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n617), .A2(new_n619), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n628), .B1(new_n623), .B2(new_n621), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n625), .A2(new_n610), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n622), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n607), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n588), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(new_n358), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(new_n486), .ZN(G1324gat));
  XOR2_X1   g437(.A(KEYINPUT16), .B(G8gat), .Z(new_n639));
  NAND4_X1  g438(.A1(new_n588), .A2(new_n635), .A3(new_n284), .A4(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n642), .A2(KEYINPUT42), .ZN(new_n643));
  OAI21_X1  g442(.A(G8gat), .B1(new_n636), .B2(new_n285), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(KEYINPUT42), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(G1325gat));
  INV_X1    g445(.A(G15gat), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n392), .A2(KEYINPUT36), .A3(new_n422), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT36), .B1(new_n392), .B2(new_n422), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT99), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n651), .B1(new_n466), .B2(new_n467), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n636), .A2(new_n647), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n392), .A2(new_n422), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n636), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n647), .B2(new_n657), .ZN(G1326gat));
  OAI21_X1  g457(.A(G22gat), .B1(new_n636), .B2(new_n418), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n588), .A2(new_n399), .A3(new_n635), .A4(new_n469), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n633), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n472), .A2(new_n476), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n626), .A2(KEYINPUT96), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n620), .A2(new_n621), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n667), .A2(new_n668), .B1(new_n669), .B2(new_n610), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n462), .A2(new_n470), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n653), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n672), .B2(new_n474), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n664), .ZN(new_n674));
  INV_X1    g473(.A(new_n607), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n666), .A2(new_n674), .A3(new_n675), .A4(new_n587), .ZN(new_n676));
  OAI21_X1  g475(.A(G29gat), .B1(new_n676), .B2(new_n358), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n588), .A2(new_n670), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n607), .ZN(new_n679));
  INV_X1    g478(.A(new_n358), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n494), .A3(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n681), .A2(KEYINPUT45), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(KEYINPUT45), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n677), .B1(new_n682), .B2(new_n683), .ZN(G1328gat));
  NAND3_X1  g483(.A1(new_n679), .A2(new_n495), .A3(new_n284), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n685), .A2(KEYINPUT46), .ZN(new_n686));
  OAI21_X1  g485(.A(G36gat), .B1(new_n676), .B2(new_n285), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(KEYINPUT46), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(G1329gat));
  NOR3_X1   g488(.A1(new_n678), .A2(new_n607), .A3(new_n656), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n653), .A2(G43gat), .ZN(new_n691));
  OAI22_X1  g490(.A1(new_n690), .A2(G43gat), .B1(new_n676), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g492(.A(G50gat), .B1(new_n676), .B2(new_n418), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT101), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT48), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n418), .A2(G50gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n694), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n696), .B(new_n699), .ZN(G1331gat));
  OAI21_X1  g499(.A(new_n433), .B1(new_n671), .B2(new_n653), .ZN(new_n701));
  INV_X1    g500(.A(new_n546), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n634), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n703), .A3(new_n586), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT102), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n701), .A2(new_n703), .A3(new_n706), .A4(new_n586), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n358), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT103), .B(G57gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1332gat));
  NAND2_X1  g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n284), .B(KEYINPUT104), .Z(new_n713));
  NAND4_X1  g512(.A1(new_n705), .A2(new_n707), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(KEYINPUT105), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(KEYINPUT105), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT106), .Z(new_n718));
  AND3_X1   g517(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n715), .B2(new_n716), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(G1333gat));
  OAI21_X1  g520(.A(new_n563), .B1(new_n708), .B2(new_n656), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n653), .A2(G71gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n708), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1334gat));
  NOR2_X1   g525(.A1(new_n708), .A2(new_n418), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(new_n564), .ZN(G1335gat));
  NOR2_X1   g527(.A1(new_n607), .A2(new_n702), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n666), .A2(new_n674), .A3(new_n586), .A4(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(G85gat), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n730), .A2(new_n731), .A3(new_n358), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n673), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(KEYINPUT108), .B(new_n670), .C1(new_n672), .C2(new_n474), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n729), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n736), .A2(KEYINPUT51), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(KEYINPUT51), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n737), .A2(new_n680), .A3(new_n586), .A4(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n732), .B1(new_n739), .B2(new_n731), .ZN(G1336gat));
  INV_X1    g539(.A(new_n713), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(G92gat), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n737), .A2(new_n586), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744));
  OAI21_X1  g543(.A(G92gat), .B1(new_n730), .B2(new_n741), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(KEYINPUT51), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n736), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n734), .A2(new_n729), .A3(new_n735), .A4(new_n749), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n751), .A2(new_n586), .A3(new_n742), .A4(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G92gat), .B1(new_n730), .B2(new_n285), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n747), .B1(new_n755), .B2(KEYINPUT52), .ZN(new_n756));
  AOI211_X1 g555(.A(KEYINPUT110), .B(new_n744), .C1(new_n753), .C2(new_n754), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n746), .B1(new_n756), .B2(new_n757), .ZN(G1337gat));
  XNOR2_X1  g557(.A(KEYINPUT111), .B(G99gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n730), .B2(new_n654), .ZN(new_n760));
  INV_X1    g559(.A(new_n759), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n737), .A2(new_n586), .A3(new_n738), .A4(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n762), .B2(new_n656), .ZN(G1338gat));
  NOR2_X1   g562(.A1(new_n418), .A2(G106gat), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n737), .A2(new_n586), .A3(new_n738), .A4(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n552), .A2(KEYINPUT112), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n552), .A2(KEYINPUT112), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n767), .B(new_n768), .C1(new_n730), .C2(new_n418), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n751), .A2(new_n586), .A3(new_n752), .A4(new_n764), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(new_n769), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n766), .B2(new_n772), .ZN(G1339gat));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n517), .A2(new_n520), .ZN(new_n775));
  INV_X1    g574(.A(new_n518), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT114), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n778), .B(new_n518), .C1(new_n517), .C2(new_n520), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n527), .A2(new_n529), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n774), .B1(new_n781), .B2(new_n536), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n575), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n570), .A2(new_n574), .A3(new_n548), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT54), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n784), .B(new_n580), .C1(new_n786), .C2(new_n575), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n582), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n787), .A2(new_n792), .A3(new_n788), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n789), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n542), .A2(new_n537), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n775), .A2(new_n776), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n778), .ZN(new_n797));
  INV_X1    g596(.A(new_n780), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n775), .A2(KEYINPUT114), .A3(new_n776), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n536), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(KEYINPUT115), .A3(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n782), .A2(new_n794), .A3(new_n795), .A4(new_n802), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n803), .A2(new_n633), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n794), .B1(new_n540), .B2(new_n545), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n782), .A2(new_n586), .A3(new_n795), .A4(new_n802), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n804), .B(KEYINPUT116), .C1(new_n807), .C2(new_n670), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n670), .B1(new_n805), .B2(new_n806), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n803), .A2(new_n633), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n808), .A2(new_n812), .A3(new_n675), .ZN(new_n813));
  INV_X1    g612(.A(new_n586), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n607), .A2(new_n633), .A3(new_n546), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n358), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n423), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n702), .A3(new_n741), .ZN(new_n819));
  NAND2_X1  g618(.A1(KEYINPUT117), .A2(G113gat), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g620(.A(KEYINPUT117), .B(G113gat), .Z(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n819), .B2(new_n822), .ZN(G1340gat));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n586), .A3(new_n741), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(G120gat), .ZN(G1341gat));
  NAND3_X1  g624(.A1(new_n818), .A2(new_n607), .A3(new_n741), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(G127gat), .ZN(G1342gat));
  NAND4_X1  g626(.A1(new_n818), .A2(new_n292), .A3(new_n670), .A4(new_n285), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(KEYINPUT56), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n818), .A2(new_n670), .A3(new_n741), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G134gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(KEYINPUT56), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(G1343gat));
  NOR3_X1   g632(.A1(new_n653), .A2(new_n358), .A3(new_n713), .ZN(new_n834));
  INV_X1    g633(.A(new_n789), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n835), .B(new_n790), .C1(new_n540), .C2(new_n545), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n670), .B1(new_n836), .B2(new_n806), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n675), .B1(new_n837), .B2(new_n811), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n418), .B1(new_n838), .B2(new_n815), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n834), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n418), .B1(new_n813), .B2(new_n815), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n310), .B1(new_n843), .B2(new_n702), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n813), .A2(new_n815), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n654), .A2(new_n469), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT118), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n846), .A2(KEYINPUT118), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n845), .A2(new_n680), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  NOR4_X1   g648(.A1(new_n849), .A2(G141gat), .A3(new_n546), .A4(new_n713), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT58), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n546), .A2(G141gat), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n816), .A2(KEYINPUT119), .A3(new_n847), .A4(new_n848), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n853), .A2(new_n741), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n845), .A2(new_n840), .A3(new_n469), .ZN(new_n857));
  INV_X1    g656(.A(new_n834), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n838), .A2(new_n815), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n469), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n858), .B1(new_n860), .B2(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G141gat), .B1(new_n862), .B2(new_n546), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n856), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n851), .A2(new_n865), .ZN(G1344gat));
  NOR2_X1   g665(.A1(new_n814), .A2(G148gat), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n853), .A2(new_n741), .A3(new_n855), .A4(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n845), .A2(new_n469), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT57), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n838), .A2(KEYINPUT121), .A3(new_n815), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT121), .B1(new_n838), .B2(new_n815), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n840), .B(new_n469), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n871), .A2(new_n586), .A3(new_n834), .A4(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n869), .B1(new_n876), .B2(G148gat), .ZN(new_n877));
  AOI211_X1 g676(.A(KEYINPUT59), .B(new_n308), .C1(new_n843), .C2(new_n586), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n868), .B1(new_n877), .B2(new_n878), .ZN(G1345gat));
  NOR3_X1   g678(.A1(new_n862), .A2(new_n314), .A3(new_n675), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n853), .A2(new_n607), .A3(new_n741), .A4(new_n855), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n314), .B2(new_n881), .ZN(G1346gat));
  NOR3_X1   g681(.A1(new_n633), .A2(G162gat), .A3(new_n284), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n853), .A2(new_n855), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n857), .A2(new_n861), .A3(new_n670), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G162gat), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT122), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1347gat));
  AOI21_X1  g690(.A(new_n680), .B1(new_n813), .B2(new_n815), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(new_n285), .A3(new_n423), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n702), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G169gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n893), .A2(new_n423), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n713), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n546), .A2(G169gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(G1348gat));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n586), .A3(new_n713), .ZN(new_n901));
  INV_X1    g700(.A(G176gat), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n814), .A2(new_n902), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n901), .A2(new_n902), .B1(new_n894), .B2(new_n903), .ZN(G1349gat));
  NAND4_X1  g703(.A1(new_n892), .A2(new_n607), .A3(new_n284), .A4(new_n817), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G183gat), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n607), .A2(new_n229), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n892), .A2(new_n817), .A3(new_n713), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g709(.A1(new_n892), .A2(new_n670), .A3(new_n284), .A4(new_n817), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n911), .A2(new_n912), .A3(G190gat), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n911), .B2(G190gat), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n670), .A2(new_n220), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n913), .A2(new_n914), .B1(new_n898), .B2(new_n915), .ZN(G1351gat));
  NOR2_X1   g715(.A1(new_n842), .A2(new_n840), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n469), .A2(new_n840), .ZN(new_n918));
  INV_X1    g717(.A(new_n874), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n872), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT124), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n875), .B(new_n922), .C1(new_n840), .C2(new_n842), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n653), .A2(new_n680), .A3(new_n285), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n921), .A2(new_n923), .A3(new_n702), .A4(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(KEYINPUT123), .B(G197gat), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n846), .A2(new_n741), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n546), .A2(new_n926), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n892), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n927), .A2(new_n930), .ZN(G1352gat));
  NAND4_X1  g730(.A1(new_n921), .A2(new_n923), .A3(new_n586), .A4(new_n924), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G204gat), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n892), .A2(new_n586), .A3(new_n928), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936));
  INV_X1    g735(.A(G204gat), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n936), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n892), .A2(new_n937), .A3(new_n586), .A4(new_n928), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n935), .A2(new_n936), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n933), .A2(new_n943), .ZN(G1353gat));
  NAND2_X1  g743(.A1(new_n871), .A2(new_n875), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n924), .A2(new_n607), .ZN(new_n946));
  OAI21_X1  g745(.A(G211gat), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT63), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n949), .B(G211gat), .C1(new_n945), .C2(new_n946), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n892), .A2(new_n203), .A3(new_n607), .A4(new_n928), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT126), .Z(new_n952));
  NAND3_X1  g751(.A1(new_n948), .A2(new_n950), .A3(new_n952), .ZN(G1354gat));
  NOR2_X1   g752(.A1(new_n633), .A2(new_n204), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n921), .A2(new_n923), .A3(new_n924), .A4(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n892), .A2(new_n670), .A3(new_n928), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n204), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n957), .A2(KEYINPUT127), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(KEYINPUT127), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(G1355gat));
endmodule


