//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  OAI221_X1 g004(.A(new_n204), .B1(KEYINPUT94), .B2(new_n205), .C1(G1gat), .C2(new_n202), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT94), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G50gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT91), .B1(new_n210), .B2(G43gat), .ZN(new_n211));
  INV_X1    g010(.A(G43gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT90), .B1(new_n212), .B2(G50gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT91), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(new_n212), .A3(G50gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT90), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(new_n210), .A3(G43gat), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n211), .A2(new_n213), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT92), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT92), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n218), .A2(new_n222), .A3(new_n219), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n210), .A2(G43gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n212), .A2(G50gat), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n224), .A2(new_n225), .A3(new_n219), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n221), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT89), .B(G29gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G36gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(G29gat), .A2(G36gat), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n231), .A2(KEYINPUT14), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(KEYINPUT14), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n228), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n226), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n209), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(new_n235), .B2(new_n237), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n218), .A2(new_n222), .A3(new_n219), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n222), .B1(new_n218), .B2(new_n219), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n242), .A2(new_n243), .A3(new_n226), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n237), .B(new_n240), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT93), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n236), .B1(new_n228), .B2(new_n234), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(KEYINPUT93), .A3(new_n240), .ZN(new_n250));
  AOI211_X1 g049(.A(new_n208), .B(new_n241), .C1(new_n248), .C2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT95), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n239), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G229gat), .A2(G233gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n238), .A2(KEYINPUT17), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT93), .B1(new_n249), .B2(new_n240), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n226), .B1(new_n220), .B2(KEYINPUT92), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n245), .B1(new_n257), .B2(new_n223), .ZN(new_n258));
  NOR4_X1   g057(.A1(new_n258), .A2(new_n247), .A3(KEYINPUT17), .A4(new_n236), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n209), .B(new_n255), .C1(new_n256), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT95), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n253), .A2(KEYINPUT18), .A3(new_n254), .A4(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n208), .B(new_n249), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n254), .B(KEYINPUT13), .Z(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n250), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(new_n252), .A3(new_n209), .A4(new_n255), .ZN(new_n268));
  INV_X1    g067(.A(new_n239), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n261), .A2(new_n254), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT18), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G113gat), .B(G141gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT11), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G197gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT12), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n266), .A2(KEYINPUT96), .A3(new_n272), .A4(new_n278), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n262), .A2(new_n272), .A3(new_n265), .A4(new_n278), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT96), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n272), .ZN(new_n284));
  INV_X1    g083(.A(new_n278), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n289));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290));
  INV_X1    g089(.A(G211gat), .ZN(new_n291));
  INV_X1    g090(.A(G218gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n290), .B1(KEYINPUT22), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G211gat), .B(G218gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n289), .B1(new_n296), .B2(KEYINPUT29), .ZN(new_n297));
  XNOR2_X1  g096(.A(G155gat), .B(G162gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT77), .ZN(new_n300));
  INV_X1    g099(.A(G155gat), .ZN(new_n301));
  INV_X1    g100(.A(G162gat), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n300), .B(KEYINPUT2), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  OR2_X1    g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(G155gat), .B2(G162gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(new_n300), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n299), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT78), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT2), .B1(new_n301), .B2(new_n302), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT78), .ZN(new_n314));
  XOR2_X1   g113(.A(G141gat), .B(G148gat), .Z(new_n315));
  NAND4_X1  g114(.A1(new_n312), .A2(new_n314), .A3(new_n298), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n296), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n314), .A2(new_n298), .A3(new_n315), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n315), .A3(new_n303), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n321), .A2(new_n312), .B1(new_n323), .B2(new_n299), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n289), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G228gat), .ZN(new_n328));
  INV_X1    g127(.A(G233gat), .ZN(new_n329));
  OAI22_X1  g128(.A1(new_n319), .A2(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n326), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT84), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT84), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n325), .A2(new_n333), .A3(new_n326), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n320), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n318), .A2(G228gat), .A3(G233gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n330), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G22gat), .ZN(new_n338));
  INV_X1    g137(.A(G22gat), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n330), .B(new_n339), .C1(new_n335), .C2(new_n336), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G78gat), .B(G106gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(G50gat), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT85), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n345), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n338), .B(new_n340), .C1(new_n346), .C2(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G1gat), .B(G29gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT0), .ZN(new_n352));
  XNOR2_X1  g151(.A(G57gat), .B(G85gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  XOR2_X1   g153(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT70), .B(G120gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G113gat), .ZN(new_n358));
  INV_X1    g157(.A(G113gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G120gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G127gat), .B(G134gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT1), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G113gat), .B(G120gat), .Z(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n363), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(KEYINPUT69), .ZN(new_n368));
  INV_X1    g167(.A(G127gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(G134gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT69), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n367), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n365), .A2(new_n373), .A3(new_n310), .A4(new_n316), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n365), .A2(new_n373), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n325), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n374), .A2(new_n383), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n366), .A2(new_n363), .B1(new_n371), .B2(new_n370), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n368), .A2(new_n385), .B1(new_n361), .B2(new_n364), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n324), .A2(new_n386), .A3(KEYINPUT79), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n379), .B(new_n382), .C1(KEYINPUT4), .C2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT80), .B1(new_n324), .B2(new_n386), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n380), .A2(new_n391), .A3(new_n317), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n388), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n389), .B(KEYINPUT5), .C1(new_n393), .C2(new_n377), .ZN(new_n394));
  INV_X1    g193(.A(new_n382), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n374), .B2(KEYINPUT4), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n324), .A2(new_n386), .A3(KEYINPUT81), .A4(new_n375), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n387), .A3(KEYINPUT4), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n378), .A2(KEYINPUT5), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI211_X1 g202(.A(new_n354), .B(new_n356), .C1(new_n394), .C2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n394), .A2(new_n354), .A3(new_n403), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n356), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n354), .B1(new_n394), .B2(new_n403), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n404), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G226gat), .A2(G233gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n412), .B(KEYINPUT76), .Z(new_n413));
  NOR2_X1   g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT23), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT23), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(G169gat), .B2(G176gat), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n417), .B2(new_n414), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(G183gat), .A2(G190gat), .ZN(new_n421));
  MUX2_X1   g220(.A(KEYINPUT24), .B(new_n420), .S(new_n421), .Z(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(KEYINPUT25), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT64), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(KEYINPUT64), .B(new_n415), .C1(new_n417), .C2(new_n414), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n422), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT65), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT25), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n427), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n423), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT66), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(KEYINPUT66), .B(new_n423), .C1(new_n430), .C2(new_n431), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(new_n414), .ZN(new_n437));
  NOR3_X1   g236(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n421), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n439), .B(KEYINPUT68), .Z(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT27), .B(G183gat), .ZN(new_n441));
  INV_X1    g240(.A(G190gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  NOR2_X1   g244(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n434), .A2(new_n435), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n413), .B1(new_n448), .B2(new_n326), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n429), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT65), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n446), .B1(new_n453), .B2(new_n423), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(new_n412), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n296), .B1(new_n449), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT30), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n435), .A2(new_n447), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT66), .B1(new_n453), .B2(new_n423), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n413), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n412), .B1(new_n454), .B2(KEYINPUT29), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n320), .ZN(new_n462));
  XNOR2_X1  g261(.A(G8gat), .B(G36gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(G64gat), .B(G92gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n456), .A2(new_n457), .A3(new_n462), .A4(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n326), .B1(new_n458), .B2(new_n459), .ZN(new_n468));
  INV_X1    g267(.A(new_n413), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n455), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n462), .B(new_n466), .C1(new_n470), .C2(new_n320), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT30), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n466), .B1(new_n456), .B2(new_n462), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n350), .B1(new_n411), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n350), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT39), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n400), .A2(new_n397), .A3(new_n398), .ZN(new_n479));
  AOI211_X1 g278(.A(new_n478), .B(new_n377), .C1(new_n479), .C2(new_n382), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n384), .A2(new_n387), .A3(KEYINPUT4), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n397), .A2(new_n398), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n382), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT86), .B1(new_n483), .B2(new_n378), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n477), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n478), .B1(new_n401), .B2(new_n377), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(KEYINPUT86), .A3(new_n378), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n477), .B1(new_n393), .B2(new_n377), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n354), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT40), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n485), .A2(new_n489), .A3(KEYINPUT40), .A4(new_n354), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n492), .A2(new_n409), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n471), .A2(KEYINPUT30), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n471), .A2(KEYINPUT30), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n462), .B1(new_n470), .B2(new_n320), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n465), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n495), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n476), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(KEYINPUT37), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT87), .B(KEYINPUT38), .Z(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT37), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n504), .B(new_n462), .C1(new_n470), .C2(new_n320), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n501), .A2(new_n465), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n460), .A2(new_n461), .A3(new_n296), .ZN(new_n507));
  OAI211_X1 g306(.A(KEYINPUT37), .B(new_n507), .C1(new_n470), .C2(new_n296), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n505), .A2(new_n508), .A3(new_n465), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n506), .B1(new_n509), .B2(new_n503), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n410), .A2(new_n471), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n475), .B1(new_n500), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G227gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(new_n329), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n386), .B1(new_n458), .B2(new_n459), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n434), .A2(new_n380), .A3(new_n435), .A4(new_n447), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI211_X1 g320(.A(new_n515), .B(new_n519), .C1(new_n516), .C2(new_n517), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n516), .A2(new_n515), .A3(new_n517), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT32), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT33), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G43gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT71), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT72), .ZN(new_n530));
  XNOR2_X1  g329(.A(G71gat), .B(G99gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n525), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n532), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n524), .B(KEYINPUT32), .C1(new_n526), .C2(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n533), .A2(KEYINPUT73), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT73), .B1(new_n533), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n523), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n521), .A2(new_n522), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(new_n533), .A3(new_n535), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n540), .A2(KEYINPUT36), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT75), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT36), .ZN(new_n544));
  INV_X1    g343(.A(new_n540), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n539), .B1(new_n535), .B2(new_n533), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n542), .B1(new_n538), .B2(new_n541), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n513), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n498), .A2(KEYINPUT30), .A3(new_n471), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n410), .B1(new_n551), .B2(new_n467), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n540), .A2(new_n350), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n538), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT35), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n533), .A2(new_n535), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n523), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n540), .A3(new_n350), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT88), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT35), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n552), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n411), .A2(new_n474), .A3(new_n561), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT88), .B1(new_n563), .B2(new_n558), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n555), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n288), .B1(new_n550), .B2(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(G57gat), .A2(G64gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(G57gat), .A2(G64gat), .ZN(new_n568));
  INV_X1    g367(.A(G71gat), .ZN(new_n569));
  INV_X1    g368(.A(G78gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n567), .B(new_n568), .C1(new_n571), .C2(KEYINPUT9), .ZN(new_n572));
  XOR2_X1   g371(.A(G71gat), .B(G78gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G127gat), .B(G155gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT20), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n580), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n574), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n208), .B1(KEYINPUT21), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT99), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n583), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G183gat), .B(G211gat), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n587), .A2(new_n589), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G99gat), .B(G106gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT100), .ZN(new_n594));
  NAND2_X1  g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT7), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n594), .B(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n249), .A2(new_n602), .B1(KEYINPUT41), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n267), .A2(new_n255), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n604), .B1(new_n605), .B2(new_n602), .ZN(new_n606));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n607), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(KEYINPUT101), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n608), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n584), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n594), .A2(new_n601), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n594), .A2(new_n601), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(new_n574), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n584), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n618), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n623), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(new_n618), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n628), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n592), .A2(new_n616), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n566), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n410), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g439(.A(G8gat), .B1(new_n637), .B2(new_n474), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT42), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT16), .B(G8gat), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n637), .A2(new_n474), .A3(new_n643), .ZN(new_n644));
  MUX2_X1   g443(.A(new_n642), .B(KEYINPUT42), .S(new_n644), .Z(G1325gat));
  INV_X1    g444(.A(G15gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n545), .A2(new_n546), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n637), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(KEYINPUT102), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(KEYINPUT102), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n548), .A2(new_n549), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n638), .A2(G15gat), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT103), .ZN(G1326gat));
  NOR2_X1   g454(.A1(new_n637), .A2(new_n350), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT43), .B(G22gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1327gat));
  NOR2_X1   g457(.A1(new_n590), .A2(new_n591), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT105), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n660), .A2(new_n288), .A3(new_n635), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n550), .A2(new_n565), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n663), .A3(new_n616), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT106), .ZN(new_n665));
  INV_X1    g464(.A(new_n616), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n550), .B2(new_n565), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n668), .A3(new_n663), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT44), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n661), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n229), .B1(new_n674), .B2(new_n411), .ZN(new_n675));
  INV_X1    g474(.A(new_n635), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n592), .A2(new_n616), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT104), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n566), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(new_n411), .A3(new_n229), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT45), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n675), .A2(new_n681), .ZN(G1328gat));
  OAI21_X1  g481(.A(G36gat), .B1(new_n674), .B2(new_n474), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n679), .A2(G36gat), .A3(new_n474), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT46), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(G1329gat));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n212), .B1(new_n673), .B2(new_n652), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n678), .A2(new_n566), .A3(new_n212), .A4(new_n647), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT107), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n687), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n652), .ZN(new_n693));
  AOI211_X1 g492(.A(new_n693), .B(new_n661), .C1(new_n670), .C2(new_n672), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n690), .B(KEYINPUT47), .C1(new_n694), .C2(new_n212), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(G1330gat));
  NAND3_X1  g495(.A1(new_n673), .A2(G50gat), .A3(new_n476), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n210), .B1(new_n679), .B2(new_n350), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n697), .A2(KEYINPUT48), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT48), .B1(new_n697), .B2(new_n698), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(G1331gat));
  NOR4_X1   g500(.A1(new_n592), .A2(new_n287), .A3(new_n616), .A4(new_n676), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n662), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n662), .A2(KEYINPUT108), .A3(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n411), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT109), .B(G57gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1332gat));
  INV_X1    g509(.A(KEYINPUT49), .ZN(new_n711));
  INV_X1    g510(.A(G64gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n499), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n707), .A2(KEYINPUT110), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT110), .B1(new_n707), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(new_n712), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1333gat));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n707), .B2(new_n648), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n705), .A2(KEYINPUT111), .A3(new_n647), .A4(new_n706), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n569), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n705), .A2(G71gat), .A3(new_n652), .A4(new_n706), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT50), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n726), .A3(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1334gat));
  NOR2_X1   g527(.A1(new_n707), .A2(new_n350), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(new_n570), .ZN(G1335gat));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n667), .A2(new_n668), .A3(new_n663), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n668), .B1(new_n667), .B2(new_n663), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n672), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n287), .A2(new_n659), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n635), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n731), .B1(new_n738), .B2(new_n411), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n736), .B1(new_n670), .B2(new_n672), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(KEYINPUT112), .A3(new_n410), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n739), .A2(G85gat), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n662), .A2(new_n743), .A3(new_n616), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(new_n735), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n667), .A2(new_n743), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(KEYINPUT51), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n744), .A2(new_n735), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(new_n746), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n410), .A2(new_n598), .A3(new_n635), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n742), .B1(new_n752), .B2(new_n753), .ZN(G1336gat));
  AOI21_X1  g553(.A(new_n599), .B1(new_n740), .B2(new_n499), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n499), .A2(new_n599), .A3(new_n635), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n748), .B2(new_n751), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT52), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n734), .A2(new_n499), .A3(new_n737), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT114), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n734), .A2(new_n761), .A3(new_n499), .A4(new_n737), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n599), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n757), .A2(KEYINPUT52), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n758), .B1(new_n763), .B2(new_n764), .ZN(G1337gat));
  OAI21_X1  g564(.A(G99gat), .B1(new_n738), .B2(new_n693), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n648), .A2(G99gat), .A3(new_n676), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n752), .B2(new_n767), .ZN(G1338gat));
  NAND3_X1  g567(.A1(new_n734), .A2(new_n476), .A3(new_n737), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n676), .A2(new_n350), .A3(G106gat), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n752), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n748), .A2(new_n751), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n772), .B(KEYINPUT115), .Z(new_n776));
  AOI22_X1  g575(.A1(new_n775), .A2(new_n776), .B1(new_n769), .B2(G106gat), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n770), .A2(new_n774), .B1(new_n777), .B2(new_n771), .ZN(G1339gat));
  NOR2_X1   g577(.A1(new_n592), .A2(new_n616), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(new_n288), .A3(new_n676), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n624), .A2(new_n625), .A3(new_n618), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT116), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n624), .A2(new_n783), .A3(new_n625), .A4(new_n618), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n626), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n632), .B1(new_n626), .B2(new_n786), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT55), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n789), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(new_n634), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n792), .A2(KEYINPUT117), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(KEYINPUT117), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n253), .A2(new_n261), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n796), .A2(new_n254), .B1(new_n263), .B2(new_n264), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n277), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n795), .A2(new_n283), .A3(new_n616), .A4(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n287), .A2(new_n795), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n280), .A2(new_n281), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n280), .A2(new_n281), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n635), .B(new_n798), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT118), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n283), .A2(new_n806), .A3(new_n635), .A4(new_n798), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n801), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n800), .B1(new_n808), .B2(new_n666), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n780), .B1(new_n809), .B2(new_n660), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n499), .A2(new_n411), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n538), .A2(new_n553), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(G113gat), .B1(new_n814), .B2(new_n287), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n559), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n359), .A3(new_n288), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n815), .A2(new_n817), .ZN(G1340gat));
  NAND2_X1  g617(.A1(new_n635), .A2(new_n357), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT119), .Z(new_n820));
  NAND2_X1  g619(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G120gat), .B1(new_n816), .B2(new_n676), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1341gat));
  AOI21_X1  g622(.A(G127gat), .B1(new_n814), .B2(new_n659), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n660), .A2(G127gat), .ZN(new_n825));
  OR3_X1    g624(.A1(new_n816), .A2(KEYINPUT120), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT120), .B1(new_n816), .B2(new_n825), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(G1342gat));
  NOR2_X1   g627(.A1(new_n666), .A2(G134gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n813), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT56), .Z(new_n831));
  OAI21_X1  g630(.A(G134gat), .B1(new_n816), .B2(new_n666), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1343gat));
  NOR3_X1   g632(.A1(new_n652), .A2(new_n411), .A3(new_n499), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT57), .B1(new_n810), .B2(new_n476), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n476), .A2(KEYINPUT57), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n791), .A2(new_n634), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(new_n790), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n283), .B2(new_n286), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n804), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n283), .A2(KEYINPUT121), .A3(new_n635), .A4(new_n798), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n799), .B1(new_n843), .B2(new_n616), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n592), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n836), .B1(new_n845), .B2(new_n780), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n287), .B(new_n834), .C1(new_n835), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(G141gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n652), .A2(new_n350), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n812), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n288), .A2(G141gat), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT58), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n848), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1344gat));
  INV_X1    g656(.A(G148gat), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n850), .A2(new_n858), .A3(new_n635), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n350), .A2(KEYINPUT57), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n844), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT122), .B(new_n799), .C1(new_n843), .C2(new_n616), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n659), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n780), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n810), .A2(new_n476), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT57), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n867), .A2(new_n635), .A3(new_n834), .A4(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n860), .B1(new_n870), .B2(G148gat), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n635), .B(new_n834), .C1(new_n835), .C2(new_n846), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n872), .A2(new_n860), .A3(G148gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n859), .B1(new_n871), .B2(new_n873), .ZN(G1345gat));
  OAI211_X1 g673(.A(new_n660), .B(new_n834), .C1(new_n835), .C2(new_n846), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G155gat), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n812), .A2(new_n301), .A3(new_n659), .A4(new_n849), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT123), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1346gat));
  OAI211_X1 g681(.A(new_n616), .B(new_n834), .C1(new_n835), .C2(new_n846), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G162gat), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n812), .A2(new_n302), .A3(new_n616), .A4(new_n849), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT124), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1347gat));
  NAND2_X1  g689(.A1(new_n499), .A2(new_n411), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n810), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n813), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n275), .B1(new_n894), .B2(new_n288), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n893), .A2(G169gat), .A3(new_n287), .A4(new_n559), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT125), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n899), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1348gat));
  INV_X1    g700(.A(new_n894), .ZN(new_n902));
  AOI21_X1  g701(.A(G176gat), .B1(new_n902), .B2(new_n635), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n893), .A2(new_n559), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n635), .A2(G176gat), .ZN(new_n906));
  OR3_X1    g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n905), .B1(new_n904), .B2(new_n906), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(G1349gat));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT127), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n893), .A2(new_n441), .A3(new_n813), .A4(new_n659), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n910), .A2(KEYINPUT127), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n893), .A2(new_n559), .A3(new_n660), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G183gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n911), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AND4_X1   g717(.A1(new_n917), .A2(new_n912), .A3(new_n914), .A4(new_n911), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(G1350gat));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n442), .A3(new_n616), .ZN(new_n921));
  OAI21_X1  g720(.A(G190gat), .B1(new_n904), .B2(new_n666), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(KEYINPUT61), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(KEYINPUT61), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(G1351gat));
  AND2_X1   g724(.A1(new_n893), .A2(new_n849), .ZN(new_n926));
  AOI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n287), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n652), .A2(new_n891), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n867), .A2(new_n869), .A3(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n287), .A2(G197gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1352gat));
  NOR2_X1   g730(.A1(new_n676), .A2(G204gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n893), .A2(new_n849), .A3(new_n932), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT62), .Z(new_n934));
  NAND4_X1  g733(.A1(new_n867), .A2(new_n635), .A3(new_n869), .A4(new_n928), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G204gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1353gat));
  NAND3_X1  g736(.A1(new_n926), .A2(new_n291), .A3(new_n659), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n867), .A2(new_n659), .A3(new_n869), .A4(new_n928), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  NAND3_X1  g741(.A1(new_n867), .A2(new_n869), .A3(new_n928), .ZN(new_n943));
  OAI21_X1  g742(.A(G218gat), .B1(new_n943), .B2(new_n666), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n292), .A3(new_n616), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1355gat));
endmodule


