

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597;

  BUF_X1 U326 ( .A(n413), .Z(n536) );
  INV_X1 U327 ( .A(KEYINPUT67), .ZN(n315) );
  XNOR2_X1 U328 ( .A(n308), .B(n307), .ZN(n310) );
  XNOR2_X1 U329 ( .A(n306), .B(n305), .ZN(n307) );
  INV_X1 U330 ( .A(KEYINPUT37), .ZN(n487) );
  NAND2_X1 U331 ( .A1(n486), .A2(n591), .ZN(n488) );
  NOR2_X1 U332 ( .A1(n498), .A2(n594), .ZN(n486) );
  XOR2_X1 U333 ( .A(n441), .B(n440), .Z(n294) );
  XOR2_X1 U334 ( .A(n397), .B(n374), .Z(n295) );
  XNOR2_X1 U335 ( .A(G22GAT), .B(G155GAT), .ZN(n371) );
  XNOR2_X1 U336 ( .A(n388), .B(KEYINPUT47), .ZN(n394) );
  XNOR2_X1 U337 ( .A(n371), .B(G78GAT), .ZN(n448) );
  XNOR2_X1 U338 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n395) );
  NOR2_X1 U339 ( .A1(n394), .A2(n393), .ZN(n396) );
  XNOR2_X1 U340 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U341 ( .A(n396), .B(n395), .ZN(n546) );
  XNOR2_X1 U342 ( .A(n404), .B(n403), .ZN(n408) );
  INV_X1 U343 ( .A(n564), .ZN(n438) );
  XNOR2_X1 U344 ( .A(n348), .B(n347), .ZN(n349) );
  OR2_X1 U345 ( .A1(n500), .A2(n532), .ZN(n489) );
  AND2_X1 U346 ( .A1(n439), .A2(n438), .ZN(n583) );
  XNOR2_X1 U347 ( .A(n316), .B(n315), .ZN(n359) );
  XNOR2_X1 U348 ( .A(n350), .B(n349), .ZN(n390) );
  XNOR2_X1 U349 ( .A(n488), .B(n487), .ZN(n532) );
  XOR2_X1 U350 ( .A(KEYINPUT38), .B(n489), .Z(n490) );
  XOR2_X1 U351 ( .A(n385), .B(n384), .Z(n591) );
  XOR2_X1 U352 ( .A(n370), .B(n369), .Z(n574) );
  XNOR2_X1 U353 ( .A(n312), .B(n311), .ZN(n548) );
  XNOR2_X1 U354 ( .A(n490), .B(KEYINPUT102), .ZN(n517) );
  XNOR2_X1 U355 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U356 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U357 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  XNOR2_X1 U358 ( .A(n494), .B(n493), .ZN(G1330GAT) );
  XNOR2_X1 U359 ( .A(G176GAT), .B(KEYINPUT18), .ZN(n296) );
  XNOR2_X1 U360 ( .A(n296), .B(KEYINPUT17), .ZN(n297) );
  XOR2_X1 U361 ( .A(n297), .B(KEYINPUT19), .Z(n299) );
  XNOR2_X1 U362 ( .A(G169GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U363 ( .A(n299), .B(n298), .ZN(n410) );
  XOR2_X1 U364 ( .A(G71GAT), .B(KEYINPUT79), .Z(n301) );
  XNOR2_X1 U365 ( .A(G183GAT), .B(KEYINPUT80), .ZN(n300) );
  XNOR2_X1 U366 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U367 ( .A(n410), .B(n302), .Z(n312) );
  XOR2_X1 U368 ( .A(G120GAT), .B(KEYINPUT0), .Z(n304) );
  XNOR2_X1 U369 ( .A(G113GAT), .B(KEYINPUT78), .ZN(n303) );
  XNOR2_X1 U370 ( .A(n304), .B(n303), .ZN(n431) );
  XOR2_X1 U371 ( .A(G43GAT), .B(G134GAT), .Z(n358) );
  XNOR2_X1 U372 ( .A(n431), .B(n358), .ZN(n308) );
  AND2_X1 U373 ( .A1(G227GAT), .A2(G233GAT), .ZN(n306) );
  INV_X1 U374 ( .A(KEYINPUT20), .ZN(n305) );
  XOR2_X1 U375 ( .A(G15GAT), .B(G127GAT), .Z(n376) );
  XNOR2_X1 U376 ( .A(G99GAT), .B(n376), .ZN(n309) );
  XNOR2_X1 U377 ( .A(n310), .B(n309), .ZN(n311) );
  INV_X1 U378 ( .A(n548), .ZN(n456) );
  XOR2_X1 U379 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n314) );
  XNOR2_X1 U380 ( .A(G36GAT), .B(G29GAT), .ZN(n313) );
  XNOR2_X1 U381 ( .A(n314), .B(n313), .ZN(n316) );
  XOR2_X1 U382 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n318) );
  XNOR2_X1 U383 ( .A(G1GAT), .B(KEYINPUT29), .ZN(n317) );
  XNOR2_X1 U384 ( .A(n318), .B(n317), .ZN(n331) );
  XOR2_X1 U385 ( .A(G22GAT), .B(G197GAT), .Z(n320) );
  XNOR2_X1 U386 ( .A(G50GAT), .B(G43GAT), .ZN(n319) );
  XNOR2_X1 U387 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U388 ( .A(G113GAT), .B(G15GAT), .Z(n322) );
  XNOR2_X1 U389 ( .A(G169GAT), .B(G141GAT), .ZN(n321) );
  XNOR2_X1 U390 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U391 ( .A(n324), .B(n323), .Z(n329) );
  XOR2_X1 U392 ( .A(KEYINPUT66), .B(KEYINPUT68), .Z(n326) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U394 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U395 ( .A(G8GAT), .B(n327), .ZN(n328) );
  XNOR2_X1 U396 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U397 ( .A(n331), .B(n330), .Z(n332) );
  XOR2_X1 U398 ( .A(n359), .B(n332), .Z(n577) );
  INV_X1 U399 ( .A(n577), .ZN(n584) );
  XNOR2_X1 U400 ( .A(G71GAT), .B(G57GAT), .ZN(n333) );
  XNOR2_X1 U401 ( .A(n333), .B(KEYINPUT13), .ZN(n375) );
  XOR2_X1 U402 ( .A(G99GAT), .B(G85GAT), .Z(n356) );
  XNOR2_X1 U403 ( .A(n375), .B(n356), .ZN(n335) );
  AND2_X1 U404 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U405 ( .A(n335), .B(n334), .ZN(n338) );
  INV_X1 U406 ( .A(n338), .ZN(n337) );
  INV_X1 U407 ( .A(KEYINPUT69), .ZN(n336) );
  NAND2_X1 U408 ( .A1(n337), .A2(n336), .ZN(n340) );
  NAND2_X1 U409 ( .A1(n338), .A2(KEYINPUT69), .ZN(n339) );
  NAND2_X1 U410 ( .A1(n340), .A2(n339), .ZN(n343) );
  XNOR2_X1 U411 ( .A(G106GAT), .B(G204GAT), .ZN(n341) );
  XNOR2_X1 U412 ( .A(n341), .B(G148GAT), .ZN(n440) );
  XOR2_X1 U413 ( .A(n440), .B(KEYINPUT33), .Z(n342) );
  XNOR2_X1 U414 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U415 ( .A(G92GAT), .B(G64GAT), .Z(n409) );
  XOR2_X1 U416 ( .A(n344), .B(n409), .Z(n350) );
  XOR2_X1 U417 ( .A(KEYINPUT32), .B(KEYINPUT70), .Z(n346) );
  XNOR2_X1 U418 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n345) );
  XNOR2_X1 U419 ( .A(n346), .B(n345), .ZN(n348) );
  XNOR2_X1 U420 ( .A(G176GAT), .B(G78GAT), .ZN(n347) );
  INV_X1 U421 ( .A(KEYINPUT41), .ZN(n351) );
  XNOR2_X1 U422 ( .A(n390), .B(n351), .ZN(n566) );
  NOR2_X1 U423 ( .A1(n584), .A2(n566), .ZN(n353) );
  INV_X1 U424 ( .A(KEYINPUT46), .ZN(n352) );
  XNOR2_X1 U425 ( .A(n353), .B(n352), .ZN(n387) );
  XOR2_X1 U426 ( .A(KEYINPUT9), .B(KEYINPUT73), .Z(n355) );
  XNOR2_X1 U427 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n354) );
  XNOR2_X1 U428 ( .A(n355), .B(n354), .ZN(n357) );
  XOR2_X1 U429 ( .A(n357), .B(n356), .Z(n361) );
  XNOR2_X1 U430 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U431 ( .A(G92GAT), .B(G106GAT), .Z(n363) );
  NAND2_X1 U432 ( .A1(G232GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U433 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U434 ( .A(n365), .B(n364), .Z(n370) );
  XOR2_X1 U435 ( .A(G50GAT), .B(G162GAT), .Z(n441) );
  XOR2_X1 U436 ( .A(KEYINPUT10), .B(KEYINPUT72), .Z(n367) );
  XNOR2_X1 U437 ( .A(G190GAT), .B(KEYINPUT74), .ZN(n366) );
  XNOR2_X1 U438 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n441), .B(n368), .ZN(n369) );
  XOR2_X1 U440 ( .A(G8GAT), .B(G183GAT), .Z(n397) );
  XOR2_X1 U441 ( .A(n448), .B(KEYINPUT14), .Z(n373) );
  NAND2_X1 U442 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U443 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n295), .B(n377), .ZN(n385) );
  XOR2_X1 U446 ( .A(KEYINPUT75), .B(G64GAT), .Z(n379) );
  XNOR2_X1 U447 ( .A(G1GAT), .B(G211GAT), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U449 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n381) );
  XNOR2_X1 U450 ( .A(KEYINPUT15), .B(KEYINPUT12), .ZN(n380) );
  XNOR2_X1 U451 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U452 ( .A(n383), .B(n382), .Z(n384) );
  XOR2_X1 U453 ( .A(KEYINPUT113), .B(n591), .Z(n580) );
  AND2_X1 U454 ( .A1(n574), .A2(n580), .ZN(n386) );
  NAND2_X1 U455 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U456 ( .A(KEYINPUT36), .B(n574), .ZN(n594) );
  NOR2_X1 U457 ( .A1(n594), .A2(n591), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n389), .B(KEYINPUT45), .ZN(n391) );
  NAND2_X1 U459 ( .A1(n391), .A2(n390), .ZN(n392) );
  NOR2_X1 U460 ( .A1(n392), .A2(n577), .ZN(n393) );
  XOR2_X1 U461 ( .A(n397), .B(G204GAT), .Z(n404) );
  XOR2_X1 U462 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n399) );
  XNOR2_X1 U463 ( .A(G197GAT), .B(G211GAT), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U465 ( .A(G218GAT), .B(KEYINPUT21), .Z(n400) );
  XOR2_X1 U466 ( .A(n401), .B(n400), .Z(n452) );
  INV_X1 U467 ( .A(n452), .ZN(n402) );
  XOR2_X1 U468 ( .A(G36GAT), .B(n402), .Z(n403) );
  XOR2_X1 U469 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n406) );
  NAND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U472 ( .A(n408), .B(n407), .Z(n412) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U474 ( .A(n412), .B(n411), .Z(n413) );
  INV_X1 U475 ( .A(n536), .ZN(n414) );
  NOR2_X1 U476 ( .A1(n546), .A2(n414), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n415), .B(KEYINPUT54), .ZN(n439) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n421) );
  XOR2_X1 U479 ( .A(KEYINPUT74), .B(G85GAT), .Z(n417) );
  XNOR2_X1 U480 ( .A(G29GAT), .B(G155GAT), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U482 ( .A(G134GAT), .B(G162GAT), .Z(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n437) );
  XOR2_X1 U485 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n423) );
  XNOR2_X1 U486 ( .A(KEYINPUT4), .B(KEYINPUT88), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n435) );
  XOR2_X1 U488 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n425) );
  XNOR2_X1 U489 ( .A(G127GAT), .B(G148GAT), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U491 ( .A(G57GAT), .B(KEYINPUT5), .Z(n427) );
  XNOR2_X1 U492 ( .A(G1GAT), .B(KEYINPUT85), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U494 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U495 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n430) );
  XNOR2_X1 U496 ( .A(n430), .B(KEYINPUT2), .ZN(n447) );
  XNOR2_X1 U497 ( .A(n431), .B(n447), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U499 ( .A(n435), .B(n434), .Z(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n564) );
  NAND2_X1 U501 ( .A1(G228GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n294), .B(n442), .ZN(n446) );
  XOR2_X1 U503 ( .A(KEYINPUT82), .B(KEYINPUT24), .Z(n444) );
  XNOR2_X1 U504 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n443) );
  XNOR2_X1 U505 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U506 ( .A(n446), .B(n445), .Z(n450) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U509 ( .A(n452), .B(n451), .Z(n468) );
  NAND2_X1 U510 ( .A1(n583), .A2(n468), .ZN(n454) );
  XOR2_X1 U511 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n455) );
  NOR2_X1 U513 ( .A1(n456), .A2(n455), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n457), .B(KEYINPUT121), .ZN(n579) );
  INV_X1 U515 ( .A(n579), .ZN(n576) );
  INV_X1 U516 ( .A(n566), .ZN(n520) );
  NAND2_X1 U517 ( .A1(n576), .A2(n520), .ZN(n461) );
  XOR2_X1 U518 ( .A(G176GAT), .B(KEYINPUT122), .Z(n459) );
  XNOR2_X1 U519 ( .A(KEYINPUT57), .B(KEYINPUT56), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  INV_X1 U522 ( .A(n574), .ZN(n495) );
  NAND2_X1 U523 ( .A1(n576), .A2(n495), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n463) );
  XNOR2_X1 U525 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n462) );
  NAND2_X1 U526 ( .A1(n390), .A2(n577), .ZN(n466) );
  XOR2_X1 U527 ( .A(n466), .B(KEYINPUT71), .Z(n500) );
  INV_X1 U528 ( .A(KEYINPUT95), .ZN(n479) );
  INV_X1 U529 ( .A(KEYINPUT27), .ZN(n467) );
  XNOR2_X1 U530 ( .A(n536), .B(n467), .ZN(n481) );
  INV_X1 U531 ( .A(n481), .ZN(n472) );
  NOR2_X1 U532 ( .A1(n468), .A2(n548), .ZN(n470) );
  XNOR2_X1 U533 ( .A(KEYINPUT92), .B(KEYINPUT26), .ZN(n469) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U535 ( .A(KEYINPUT91), .B(n471), .Z(n582) );
  NAND2_X1 U536 ( .A1(n472), .A2(n582), .ZN(n562) );
  XNOR2_X1 U537 ( .A(n562), .B(KEYINPUT93), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n548), .A2(n536), .ZN(n473) );
  NAND2_X1 U539 ( .A1(n473), .A2(n468), .ZN(n474) );
  XNOR2_X1 U540 ( .A(n474), .B(KEYINPUT94), .ZN(n475) );
  XNOR2_X1 U541 ( .A(KEYINPUT25), .B(n475), .ZN(n476) );
  NOR2_X1 U542 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U543 ( .A(n479), .B(n478), .ZN(n480) );
  NOR2_X1 U544 ( .A1(n480), .A2(n564), .ZN(n485) );
  XOR2_X1 U545 ( .A(n468), .B(KEYINPUT28), .Z(n541) );
  NOR2_X1 U546 ( .A1(n541), .A2(n481), .ZN(n482) );
  NAND2_X1 U547 ( .A1(n564), .A2(n482), .ZN(n547) );
  XOR2_X1 U548 ( .A(KEYINPUT81), .B(n548), .Z(n483) );
  NOR2_X1 U549 ( .A1(n547), .A2(n483), .ZN(n484) );
  NOR2_X1 U550 ( .A1(n485), .A2(n484), .ZN(n498) );
  NAND2_X1 U551 ( .A1(n517), .A2(n548), .ZN(n494) );
  XOR2_X1 U552 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n492) );
  INV_X1 U553 ( .A(G43GAT), .ZN(n491) );
  XOR2_X1 U554 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n502) );
  NOR2_X1 U555 ( .A1(n495), .A2(n591), .ZN(n496) );
  XOR2_X1 U556 ( .A(KEYINPUT16), .B(n496), .Z(n497) );
  NOR2_X1 U557 ( .A1(n498), .A2(n497), .ZN(n499) );
  XOR2_X1 U558 ( .A(KEYINPUT96), .B(n499), .Z(n521) );
  NOR2_X1 U559 ( .A1(n521), .A2(n500), .ZN(n510) );
  NAND2_X1 U560 ( .A1(n510), .A2(n564), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U562 ( .A(G1GAT), .B(n503), .ZN(G1324GAT) );
  NAND2_X1 U563 ( .A1(n536), .A2(n510), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n504), .B(KEYINPUT98), .ZN(n505) );
  XNOR2_X1 U565 ( .A(G8GAT), .B(n505), .ZN(G1325GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n507) );
  NAND2_X1 U567 ( .A1(n510), .A2(n548), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(n509) );
  XOR2_X1 U569 ( .A(G15GAT), .B(KEYINPUT99), .Z(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(G1326GAT) );
  XOR2_X1 U571 ( .A(G22GAT), .B(KEYINPUT101), .Z(n512) );
  NAND2_X1 U572 ( .A1(n510), .A2(n541), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n512), .B(n511), .ZN(G1327GAT) );
  XOR2_X1 U574 ( .A(G29GAT), .B(KEYINPUT39), .Z(n514) );
  NAND2_X1 U575 ( .A1(n517), .A2(n564), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n514), .B(n513), .ZN(G1328GAT) );
  XOR2_X1 U577 ( .A(G36GAT), .B(KEYINPUT103), .Z(n516) );
  NAND2_X1 U578 ( .A1(n517), .A2(n536), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1329GAT) );
  XOR2_X1 U580 ( .A(G50GAT), .B(KEYINPUT105), .Z(n519) );
  NAND2_X1 U581 ( .A1(n517), .A2(n541), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(G1331GAT) );
  NAND2_X1 U583 ( .A1(n520), .A2(n584), .ZN(n531) );
  NOR2_X1 U584 ( .A1(n521), .A2(n531), .ZN(n522) );
  XNOR2_X1 U585 ( .A(KEYINPUT106), .B(n522), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n527), .A2(n564), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(KEYINPUT42), .ZN(n524) );
  XNOR2_X1 U588 ( .A(G57GAT), .B(n524), .ZN(G1332GAT) );
  NAND2_X1 U589 ( .A1(n527), .A2(n536), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U591 ( .A1(n527), .A2(n548), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n529) );
  NAND2_X1 U594 ( .A1(n541), .A2(n527), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U596 ( .A(G78GAT), .B(n530), .Z(G1335GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n534) );
  NOR2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n542), .A2(n564), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G85GAT), .B(n535), .ZN(G1336GAT) );
  NAND2_X1 U602 ( .A1(n536), .A2(n542), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n537), .B(KEYINPUT110), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G92GAT), .B(n538), .ZN(G1337GAT) );
  XOR2_X1 U605 ( .A(G99GAT), .B(KEYINPUT111), .Z(n540) );
  NAND2_X1 U606 ( .A1(n542), .A2(n548), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1338GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n544) );
  NAND2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(G106GAT), .B(n545), .Z(G1339GAT) );
  NOR2_X1 U612 ( .A1(n546), .A2(n547), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n558) );
  NOR2_X1 U614 ( .A1(n584), .A2(n558), .ZN(n550) );
  XOR2_X1 U615 ( .A(G113GAT), .B(n550), .Z(G1340GAT) );
  NOR2_X1 U616 ( .A1(n558), .A2(n566), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n552) );
  XNOR2_X1 U618 ( .A(G120GAT), .B(KEYINPUT115), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1341GAT) );
  NOR2_X1 U621 ( .A1(n580), .A2(n558), .ZN(n556) );
  XNOR2_X1 U622 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(G127GAT), .B(n557), .Z(G1342GAT) );
  NOR2_X1 U625 ( .A1(n574), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(G134GAT), .B(n561), .Z(G1343GAT) );
  NOR2_X1 U629 ( .A1(n546), .A2(n562), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n573) );
  NOR2_X1 U631 ( .A1(n584), .A2(n573), .ZN(n565) );
  XOR2_X1 U632 ( .A(G141GAT), .B(n565), .Z(G1344GAT) );
  NOR2_X1 U633 ( .A1(n566), .A2(n573), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G148GAT), .B(n569), .ZN(G1345GAT) );
  NOR2_X1 U637 ( .A1(n591), .A2(n573), .ZN(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U640 ( .A(G155GAT), .B(n572), .ZN(G1346GAT) );
  NOR2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U642 ( .A(G162GAT), .B(n575), .Z(G1347GAT) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(G169GAT), .B(n578), .ZN(G1348GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G183GAT), .B(n581), .Z(G1350GAT) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n593) );
  NOR2_X1 U648 ( .A1(n584), .A2(n593), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G197GAT), .B(n587), .ZN(G1352GAT) );
  NOR2_X1 U652 ( .A1(n390), .A2(n593), .ZN(n589) );
  XNOR2_X1 U653 ( .A(KEYINPUT61), .B(KEYINPUT125), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U655 ( .A(G204GAT), .B(n590), .Z(G1353GAT) );
  NOR2_X1 U656 ( .A1(n591), .A2(n593), .ZN(n592) );
  XOR2_X1 U657 ( .A(G211GAT), .B(n592), .Z(G1354GAT) );
  NOR2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n596) );
  XNOR2_X1 U659 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n595) );
  XNOR2_X1 U660 ( .A(n596), .B(n595), .ZN(n597) );
  XOR2_X1 U661 ( .A(G218GAT), .B(n597), .Z(G1355GAT) );
endmodule

