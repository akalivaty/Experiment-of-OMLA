//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT67), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n467), .A2(new_n464), .A3(G101), .A4(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n463), .A2(G137), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  OR2_X1    g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n472), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n469), .B1(new_n464), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n462), .A2(new_n464), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n464), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OR3_X1    g055(.A1(new_n462), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT68), .B1(new_n462), .B2(G2105), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n480), .B1(new_n483), .B2(G136), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT69), .ZN(G162));
  NAND2_X1  g060(.A1(new_n464), .A2(G138), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n470), .B2(new_n471), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT70), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n460), .B2(new_n461), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n488), .A2(KEYINPUT71), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n472), .A2(new_n499), .A3(KEYINPUT72), .A4(new_n492), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n493), .A2(new_n501), .A3(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n489), .A2(new_n495), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(G2105), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n506), .B1(new_n476), .B2(G126), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT73), .B1(new_n514), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(G543), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n519), .A2(G88), .A3(new_n520), .A4(new_n510), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n513), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n516), .B1(KEYINPUT5), .B2(new_n517), .ZN(new_n526));
  NOR3_X1   g101(.A1(new_n514), .A2(KEYINPUT73), .A3(G543), .ZN(new_n527));
  OAI211_X1 g102(.A(G62), .B(new_n520), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n519), .A2(KEYINPUT74), .A3(G62), .A4(new_n520), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n523), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n522), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI211_X1 g109(.A(KEYINPUT75), .B(new_n523), .C1(new_n530), .C2(new_n531), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(G166));
  AND2_X1   g111(.A1(new_n519), .A2(new_n520), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n537), .A2(G89), .A3(new_n510), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(G63), .A3(G651), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT76), .B(KEYINPUT7), .Z(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n512), .A2(G51), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n538), .A2(new_n539), .A3(new_n542), .A4(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  AOI22_X1  g120(.A1(new_n537), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n523), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n512), .A2(G52), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n537), .A2(new_n510), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n547), .A2(new_n551), .ZN(G171));
  AOI22_X1  g127(.A1(new_n537), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n523), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n512), .A2(G43), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n549), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n519), .A2(new_n520), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OR3_X1    g144(.A1(new_n511), .A2(KEYINPUT9), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n511), .B2(new_n569), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n549), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n537), .A2(KEYINPUT77), .A3(new_n510), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G91), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n568), .B(new_n572), .C1(new_n576), .C2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  NAND2_X1  g154(.A1(new_n528), .A2(new_n529), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n580), .A2(new_n531), .A3(new_n524), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT75), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n532), .A2(new_n533), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n583), .A2(new_n584), .A3(new_n522), .ZN(G303));
  NAND3_X1  g160(.A1(new_n574), .A2(G87), .A3(new_n575), .ZN(new_n586));
  INV_X1    g161(.A(G74), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n523), .B1(new_n565), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(G49), .B2(new_n512), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G288));
  NAND3_X1  g166(.A1(new_n574), .A2(G86), .A3(new_n575), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n519), .A2(G61), .A3(new_n520), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n523), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n595), .A2(new_n596), .B1(new_n512), .B2(G48), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n592), .A2(new_n597), .A3(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n537), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n523), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n512), .A2(G47), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n549), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n601), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n576), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n574), .A2(KEYINPUT10), .A3(G92), .A4(new_n575), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n565), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(new_n512), .B2(G54), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G321));
  XNOR2_X1  g193(.A(G321), .B(KEYINPUT79), .ZN(G284));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT80), .ZN(G148));
  NAND3_X1  g201(.A1(new_n611), .A2(new_n624), .A3(new_n615), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n476), .A2(G123), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT81), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n483), .A2(G135), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n637), .A2(new_n638), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT82), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT83), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n654), .A2(new_n660), .A3(new_n656), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n659), .B2(new_n661), .ZN(G401));
  XNOR2_X1  g237(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT84), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n663), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  INV_X1    g247(.A(new_n668), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n671), .B(new_n672), .C1(new_n663), .C2(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n671), .B2(new_n672), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT86), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n680), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n680), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n689), .B(new_n690), .Z(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G33), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n481), .A2(G139), .A3(new_n482), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT25), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(KEYINPUT92), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT92), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n699), .A2(new_n704), .A3(new_n701), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(new_n464), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n698), .B1(new_n709), .B2(new_n697), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n710), .A2(KEYINPUT93), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(KEYINPUT93), .ZN(new_n712));
  AOI21_X1  g287(.A(G2072), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n483), .A2(G141), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT26), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n715), .B(new_n717), .C1(G129), .C2(new_n476), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(new_n697), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n697), .B2(G32), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT27), .B(G1996), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT24), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n697), .B1(new_n724), .B2(G34), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n724), .B2(G34), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G160), .B2(G29), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n727), .A2(G2084), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n713), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n711), .A2(G2072), .A3(new_n712), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(KEYINPUT94), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(KEYINPUT94), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT95), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n729), .B(KEYINPUT95), .C1(new_n731), .C2(new_n732), .ZN(new_n736));
  INV_X1    g311(.A(G16), .ZN(new_n737));
  NOR2_X1   g312(.A1(G168), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n737), .B2(G21), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT96), .B(G1966), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT97), .Z(new_n742));
  OAI22_X1  g317(.A1(new_n721), .A2(new_n722), .B1(new_n739), .B2(new_n740), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT30), .B(G28), .ZN(new_n744));
  OR2_X1    g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  NAND2_X1  g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n744), .A2(new_n697), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n747), .B1(new_n727), .B2(G2084), .C1(new_n636), .C2(new_n697), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n697), .A2(G35), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n697), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n752));
  INV_X1    g327(.A(G2090), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n751), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n742), .A2(new_n749), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G4), .A2(G16), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT91), .Z(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n617), .B2(G16), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1348), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n697), .A2(G26), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT28), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n483), .A2(G140), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n764));
  INV_X1    g339(.A(G116), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G2105), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n476), .B2(G128), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(G29), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G1341), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT89), .B(G16), .Z(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n558), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G19), .B2(new_n774), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n771), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT23), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n621), .B2(new_n737), .ZN(new_n780));
  INV_X1    g355(.A(G1956), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n737), .A2(G5), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G171), .B2(new_n737), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1961), .ZN(new_n785));
  INV_X1    g360(.A(G2078), .ZN(new_n786));
  NAND2_X1  g361(.A1(G164), .A2(G29), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G27), .B2(G29), .ZN(new_n788));
  OAI22_X1  g363(.A1(new_n776), .A2(new_n772), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n786), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n777), .A2(new_n782), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n756), .A2(new_n760), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n735), .A2(new_n736), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G25), .A2(G29), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n476), .A2(G119), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n464), .A2(G107), .ZN(new_n797));
  OAI21_X1  g372(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n481), .A2(new_n482), .ZN(new_n799));
  INV_X1    g374(.A(G131), .ZN(new_n800));
  OAI221_X1 g375(.A(new_n796), .B1(new_n797), .B2(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT87), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n795), .B1(new_n804), .B2(G29), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT35), .B(G1991), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT88), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n805), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n774), .A2(G24), .ZN(new_n810));
  INV_X1    g385(.A(G290), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n774), .ZN(new_n812));
  INV_X1    g387(.A(G1986), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n737), .A2(G23), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n590), .B2(new_n737), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n818));
  INV_X1    g393(.A(G1976), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT33), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(new_n816), .C1(new_n590), .C2(new_n737), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n819), .B1(new_n818), .B2(new_n821), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n774), .A2(G22), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G166), .B2(new_n774), .ZN(new_n826));
  INV_X1    g401(.A(G1971), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  MUX2_X1   g403(.A(G6), .B(G305), .S(G16), .Z(new_n829));
  XOR2_X1   g404(.A(KEYINPUT32), .B(G1981), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n824), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT34), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n815), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n824), .A2(new_n828), .A3(new_n831), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT90), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT34), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n836), .B1(new_n835), .B2(KEYINPUT34), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n834), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT36), .ZN(new_n841));
  OAI21_X1  g416(.A(KEYINPUT90), .B1(new_n832), .B2(new_n833), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n837), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n843), .A2(new_n844), .A3(new_n834), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n794), .B1(new_n841), .B2(new_n845), .ZN(G311));
  INV_X1    g421(.A(new_n794), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n840), .A2(KEYINPUT36), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n844), .B1(new_n843), .B2(new_n834), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(G150));
  NAND2_X1  g425(.A1(new_n617), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n537), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(new_n523), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n512), .A2(G55), .ZN(new_n855));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n549), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(KEYINPUT99), .B2(new_n558), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n558), .A2(KEYINPUT99), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n861), .B1(new_n558), .B2(KEYINPUT99), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n554), .A2(new_n557), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n858), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n869), .A3(new_n862), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n852), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n852), .A2(new_n871), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n875));
  XOR2_X1   g450(.A(KEYINPUT101), .B(G860), .Z(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n874), .B2(KEYINPUT39), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n874), .A2(new_n878), .A3(KEYINPUT39), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n859), .A2(new_n876), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT37), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(G145));
  XNOR2_X1  g459(.A(G162), .B(G160), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n636), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n768), .A2(new_n508), .ZN(new_n887));
  NAND3_X1  g462(.A1(G164), .A2(new_n763), .A3(new_n767), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n709), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n706), .A2(new_n708), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n887), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n719), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n476), .A2(G130), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n464), .A2(G118), .ZN(new_n897));
  OAI21_X1  g472(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n898));
  INV_X1    g473(.A(G142), .ZN(new_n899));
  OAI221_X1 g474(.A(new_n896), .B1(new_n897), .B2(new_n898), .C1(new_n799), .C2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n640), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n803), .B(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n890), .A2(new_n719), .A3(new_n892), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n895), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n886), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n895), .A2(new_n903), .ZN(new_n907));
  INV_X1    g482(.A(new_n902), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(G37), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n904), .A2(KEYINPUT103), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n895), .A2(new_n902), .A3(new_n912), .A4(new_n903), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n913), .A3(new_n909), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n914), .A2(KEYINPUT104), .A3(new_n886), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT104), .B1(new_n914), .B2(new_n886), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g493(.A1(new_n616), .A2(G299), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n621), .B1(new_n611), .B2(new_n615), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n919), .B2(new_n920), .ZN(new_n924));
  INV_X1    g499(.A(new_n627), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n871), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n627), .B1(new_n865), .B2(new_n870), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n923), .B(new_n924), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n919), .ZN(new_n929));
  INV_X1    g504(.A(new_n920), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(KEYINPUT41), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n919), .B2(new_n920), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n871), .B(new_n925), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n928), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n811), .B(new_n590), .ZN(new_n938));
  XNOR2_X1  g513(.A(G303), .B(G305), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(KEYINPUT106), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n928), .B(new_n942), .C1(new_n934), .C2(new_n935), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n937), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n937), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g520(.A(G868), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n858), .A2(G868), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(G295));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n947), .ZN(G331));
  XNOR2_X1  g524(.A(G171), .B(G168), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n865), .A2(new_n870), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n950), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n871), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n924), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n951), .B(new_n953), .C1(new_n954), .C2(new_n922), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n865), .A2(new_n870), .A3(new_n950), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n950), .B1(new_n865), .B2(new_n870), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n931), .B(new_n933), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n940), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(G37), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n953), .A2(new_n930), .A3(new_n929), .A4(new_n951), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n958), .A2(new_n963), .A3(new_n940), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n961), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n962), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n940), .B1(new_n958), .B2(new_n963), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OR3_X1    g546(.A1(new_n966), .A2(KEYINPUT43), .A3(new_n967), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT43), .B1(new_n966), .B2(new_n959), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(KEYINPUT44), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(G397));
  XNOR2_X1  g550(.A(new_n719), .B(G1996), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n768), .B(new_n770), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n804), .A2(new_n808), .ZN(new_n979));
  OAI22_X1  g554(.A1(new_n978), .A2(new_n979), .B1(G2067), .B2(new_n768), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n508), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n469), .B(G40), .C1(new_n464), .C2(new_n473), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n977), .A2(new_n719), .ZN(new_n989));
  OR3_X1    g564(.A1(new_n984), .A2(G1996), .A3(new_n985), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n989), .A2(new_n986), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n991), .B2(new_n990), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n978), .B1(new_n807), .B2(new_n803), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n979), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n986), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n986), .A2(new_n813), .A3(new_n811), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(KEYINPUT48), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT48), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  OAI221_X1 g576(.A(new_n987), .B1(new_n988), .B2(new_n993), .C1(new_n999), .C2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n988), .B2(new_n993), .ZN(new_n1003));
  INV_X1    g578(.A(G8), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n503), .B2(new_n507), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n985), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n982), .B2(new_n983), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1005), .A2(KEYINPUT109), .A3(KEYINPUT45), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n827), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n1012));
  INV_X1    g587(.A(new_n985), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1005), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1012), .A2(new_n753), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1004), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(G8), .B1(new_n534), .B2(new_n535), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT110), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n1021));
  NAND4_X1  g596(.A1(G303), .A2(new_n1021), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1022));
  OAI211_X1 g597(.A(KEYINPUT55), .B(G8), .C1(new_n534), .C2(new_n535), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT111), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1020), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1024), .A2(new_n1022), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1017), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n592), .A2(new_n1030), .A3(new_n598), .A4(new_n597), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n512), .A2(G48), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT113), .B(G86), .Z(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n549), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(G1981), .B1(new_n1034), .B2(new_n595), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1004), .B1(new_n1013), .B2(new_n1005), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(new_n1037), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n586), .A2(G1976), .A3(new_n589), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1045), .A2(KEYINPUT112), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1976), .B1(new_n586), .B2(new_n589), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1046), .B(new_n1041), .C1(KEYINPUT52), .C2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT52), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1041), .A2(KEYINPUT112), .A3(new_n1045), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1040), .A2(new_n1044), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n982), .A2(new_n1007), .A3(new_n983), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT109), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1971), .B1(new_n1055), .B2(new_n1006), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1016), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1024), .A2(new_n1022), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1020), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1058), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1029), .A2(new_n1052), .A3(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n786), .B(new_n1006), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1013), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1068));
  AOI211_X1 g643(.A(KEYINPUT50), .B(G1384), .C1(new_n503), .C2(new_n507), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT118), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1012), .A2(new_n1071), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1072));
  INV_X1    g647(.A(G1961), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n984), .A2(new_n1006), .A3(KEYINPUT53), .A4(new_n786), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1067), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G171), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1068), .A2(G2084), .A3(new_n1069), .ZN(new_n1078));
  INV_X1    g653(.A(new_n740), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n984), .B2(new_n1006), .ZN(new_n1080));
  OAI21_X1  g655(.A(G168), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1013), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1005), .A2(KEYINPUT45), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n740), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G2084), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1012), .A2(new_n1086), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(G286), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1081), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(new_n1004), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1085), .A2(G168), .A3(new_n1087), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G8), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1089), .A2(new_n1091), .B1(new_n1093), .B2(new_n1090), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1077), .B1(new_n1094), .B2(KEYINPUT62), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT51), .B1(new_n1092), .B2(G8), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1064), .A2(new_n1095), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1041), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G288), .A2(G1976), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1031), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1101), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT115), .B(new_n1031), .C1(new_n1102), .C2(new_n1104), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1029), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1107), .A2(new_n1108), .B1(new_n1109), .B2(new_n1052), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1081), .A2(new_n1004), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1029), .A2(new_n1063), .A3(new_n1052), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT63), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1100), .B(new_n1110), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  AND4_X1   g691(.A1(new_n1029), .A2(new_n1094), .A3(new_n1052), .A4(new_n1063), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n786), .A2(KEYINPUT123), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n786), .A2(KEYINPUT123), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1066), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n984), .A2(new_n1006), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n984), .A2(new_n1006), .A3(KEYINPUT124), .A4(new_n1121), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(new_n1067), .A3(new_n1074), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1118), .B1(new_n1127), .B2(G171), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1067), .A2(new_n1074), .A3(new_n1075), .A4(G301), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1128), .A2(KEYINPUT126), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1117), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1126), .A2(new_n1067), .A3(G301), .A4(new_n1074), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1077), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT125), .B1(new_n1134), .B2(new_n1118), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1136), .B(KEYINPUT54), .C1(new_n1077), .C2(new_n1133), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n1140));
  INV_X1    g715(.A(G1348), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1070), .A2(new_n1072), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1013), .A2(new_n1005), .A3(new_n770), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n616), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT56), .B(G2072), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1006), .B(new_n1145), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1055), .A2(KEYINPUT117), .A3(new_n1006), .A4(new_n1145), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n781), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1148), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(G299), .A2(KEYINPUT116), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT57), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1144), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1146), .A2(new_n1147), .B1(new_n781), .B2(new_n1150), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(new_n1154), .A3(new_n1149), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1140), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1154), .B1(new_n1157), .B2(new_n1149), .ZN(new_n1161));
  OAI211_X1 g736(.A(KEYINPUT119), .B(new_n1158), .C1(new_n1161), .C2(new_n1144), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT122), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT61), .B1(new_n1168), .B2(new_n1158), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT60), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1170), .A2(new_n617), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1013), .A2(new_n1005), .ZN(new_n1173));
  XOR2_X1   g748(.A(KEYINPUT58), .B(G1341), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(KEYINPUT120), .B(G1996), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1175), .B1(new_n1010), .B2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n558), .A2(KEYINPUT121), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1177), .A2(KEYINPUT59), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT59), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1172), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1164), .A2(KEYINPUT61), .A3(new_n1158), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n616), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1183), .B1(new_n1171), .B2(new_n1170), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1163), .B1(new_n1169), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1116), .B1(new_n1139), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n986), .A2(G1986), .A3(G290), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n997), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT108), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n996), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1003), .B1(new_n1187), .B2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g767(.A(G319), .ZN(new_n1194));
  OR2_X1    g768(.A1(G227), .A2(new_n1194), .ZN(new_n1195));
  OR3_X1    g769(.A1(G401), .A2(new_n1195), .A3(KEYINPUT127), .ZN(new_n1196));
  OAI21_X1  g770(.A(KEYINPUT127), .B1(G401), .B2(new_n1195), .ZN(new_n1197));
  AND3_X1   g771(.A1(new_n1196), .A2(new_n695), .A3(new_n1197), .ZN(new_n1198));
  NAND3_X1  g772(.A1(new_n969), .A2(new_n917), .A3(new_n1198), .ZN(G225));
  INV_X1    g773(.A(G225), .ZN(G308));
endmodule


