//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(KEYINPUT69), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n465), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT70), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT71), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  AOI211_X1 g051(.A(new_n475), .B(new_n476), .C1(new_n470), .C2(new_n472), .ZN(new_n477));
  OR2_X1    g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n463), .A2(new_n464), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(G137), .A3(new_n476), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n481));
  INV_X1    g056(.A(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G101), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n481), .B1(new_n480), .B2(new_n484), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  NOR2_X1   g064(.A1(new_n467), .A2(new_n468), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(new_n476), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT74), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n490), .B2(new_n476), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G124), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT73), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n490), .B2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n479), .A2(KEYINPUT73), .A3(new_n476), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G136), .ZN(new_n502));
  OR2_X1    g077(.A1(G100), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n496), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G162));
  NAND2_X1  g081(.A1(new_n476), .A2(G138), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n507), .B1(new_n463), .B2(new_n464), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT75), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT75), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n511), .B(KEYINPUT4), .C1(new_n490), .C2(new_n507), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n465), .A2(new_n469), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n516));
  INV_X1    g091(.A(G114), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(G2105), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(new_n491), .B2(G126), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT76), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT76), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n515), .A2(new_n522), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(G164));
  OR2_X1    g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n528), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT6), .B(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G88), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G50), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n531), .A2(new_n537), .ZN(G166));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  INV_X1    g115(.A(G51), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n526), .A2(new_n527), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n532), .A2(G89), .ZN(new_n544));
  NAND2_X1  g119(.A1(G63), .A2(G651), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(G168));
  AOI22_X1  g122(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n530), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n533), .A2(new_n550), .B1(new_n535), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(G171));
  AOI22_X1  g128(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n530), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  INV_X1    g131(.A(G43), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n533), .A2(new_n556), .B1(new_n535), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n543), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n533), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n567), .A2(G651), .B1(new_n568), .B2(G91), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n532), .A2(KEYINPUT77), .A3(G53), .A4(G543), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  NAND3_X1  g151(.A1(new_n532), .A2(G49), .A3(G543), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT78), .Z(new_n578));
  OR2_X1    g153(.A1(new_n528), .A2(G74), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n568), .A2(G87), .B1(new_n579), .B2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n526), .B2(new_n527), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n528), .A2(new_n532), .A3(G86), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n532), .A2(G48), .A3(G543), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n530), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT80), .B(G47), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n533), .A2(new_n593), .B1(new_n535), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n568), .A2(G92), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT10), .Z(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n543), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n535), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n603), .A2(G651), .B1(new_n604), .B2(G54), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NOR2_X1   g190(.A1(new_n606), .A2(G559), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  OR3_X1    g192(.A1(new_n616), .A2(KEYINPUT81), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT81), .B1(new_n616), .B2(new_n617), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n618), .B(new_n619), .C1(G868), .C2(new_n559), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n495), .A2(G123), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n501), .A2(G135), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(G111), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n624), .A2(KEYINPUT82), .B1(new_n625), .B2(G2105), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(KEYINPUT82), .B2(new_n624), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n622), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT83), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n465), .A2(new_n469), .A3(new_n483), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT13), .B(G2100), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n630), .A2(new_n634), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT85), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n646), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  INV_X1    g235(.A(new_n653), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n660), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(KEYINPUT87), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT19), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(KEYINPUT87), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  INV_X1    g249(.A(new_n671), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n666), .A2(new_n667), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n668), .A3(new_n677), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n674), .B(new_n678), .C1(new_n675), .C2(new_n677), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G33), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n501), .A2(G139), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT94), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT25), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n469), .A3(G127), .ZN(new_n692));
  INV_X1    g267(.A(G115), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n482), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n691), .B1(new_n694), .B2(G2105), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n687), .B1(new_n697), .B2(new_n686), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(G2072), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n495), .A2(G129), .ZN(new_n700));
  NAND3_X1  g275(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT95), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT26), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n483), .A2(G105), .ZN(new_n705));
  INV_X1    g280(.A(G141), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n500), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(new_n686), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n686), .B2(G32), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT27), .B(G1996), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G2084), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n686), .B1(KEYINPUT24), .B2(G34), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(KEYINPUT24), .B2(G34), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n488), .B2(G29), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n699), .B(new_n712), .C1(new_n713), .C2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT96), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G23), .ZN(new_n720));
  INV_X1    g295(.A(G288), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT33), .B(G1976), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n719), .A2(G22), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G166), .B2(new_n719), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(G1971), .Z(new_n727));
  MUX2_X1   g302(.A(G6), .B(G305), .S(G16), .Z(new_n728));
  XOR2_X1   g303(.A(KEYINPUT32), .B(G1981), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n724), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT89), .B(KEYINPUT34), .Z(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n686), .A2(G25), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n495), .A2(G119), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n501), .A2(G131), .ZN(new_n737));
  OR2_X1    g312(.A1(G95), .A2(G2105), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n738), .B(G2104), .C1(G107), .C2(new_n476), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n686), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT35), .B(G1991), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n719), .A2(G24), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n596), .B2(new_n719), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT88), .B(G1986), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n734), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n731), .A2(new_n733), .ZN(new_n750));
  OAI22_X1  g325(.A1(new_n749), .A2(new_n750), .B1(KEYINPUT90), .B2(KEYINPUT36), .ZN(new_n751));
  NAND2_X1  g326(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT91), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n751), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n686), .A2(G26), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n495), .A2(G128), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n501), .A2(G140), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n760));
  AND3_X1   g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n756), .B1(new_n761), .B2(new_n686), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT92), .Z(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G2067), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G2067), .ZN(new_n765));
  NOR2_X1   g340(.A1(G4), .A2(G16), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n607), .B2(G16), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G1348), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n719), .A2(G19), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n559), .B2(new_n719), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1341), .ZN(new_n771));
  INV_X1    g346(.A(new_n767), .ZN(new_n772));
  INV_X1    g347(.A(G1348), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n764), .A2(new_n765), .A3(new_n768), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT93), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n686), .A2(G35), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G162), .B2(new_n686), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT29), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2090), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n686), .A2(G27), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n686), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n782), .A2(G2078), .B1(new_n716), .B2(new_n713), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G2078), .B2(new_n782), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT31), .B(G11), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT98), .ZN(new_n786));
  INV_X1    g361(.A(G28), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n787), .B2(KEYINPUT30), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(KEYINPUT30), .B2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G171), .A2(new_n719), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G5), .B2(new_n719), .ZN(new_n792));
  INV_X1    g367(.A(G1961), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n719), .A2(G21), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G168), .B2(new_n719), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT97), .B(G1966), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n794), .B(new_n798), .C1(new_n793), .C2(new_n792), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n719), .A2(G20), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT23), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n611), .B2(new_n719), .ZN(new_n802));
  INV_X1    g377(.A(G1956), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  OAI221_X1 g379(.A(new_n804), .B1(new_n686), .B2(new_n629), .C1(new_n710), .C2(new_n711), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n780), .A2(new_n784), .A3(new_n799), .A4(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n718), .A2(new_n754), .A3(new_n776), .A4(new_n806), .ZN(G150));
  INV_X1    g382(.A(G150), .ZN(G311));
  AOI22_X1  g383(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(new_n530), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT100), .B(G93), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT99), .B(G55), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n604), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(KEYINPUT101), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n812), .B2(new_n814), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n810), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G860), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT37), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n607), .A2(G559), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT38), .ZN(new_n823));
  INV_X1    g398(.A(new_n559), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n559), .B(new_n810), .C1(new_n816), .C2(new_n818), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n823), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT102), .ZN(new_n831));
  INV_X1    g406(.A(G860), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n829), .B2(KEYINPUT39), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n821), .B1(new_n831), .B2(new_n833), .ZN(G145));
  XNOR2_X1  g409(.A(new_n629), .B(new_n505), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n488), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n708), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n839));
  INV_X1    g414(.A(new_n520), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n838), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n761), .A2(new_n520), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n845), .A2(new_n708), .A3(new_n841), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n696), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT104), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n845), .A2(new_n708), .A3(new_n841), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n708), .B1(new_n845), .B2(new_n841), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT103), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT103), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n844), .A2(new_n852), .A3(new_n846), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n848), .B1(new_n854), .B2(new_n697), .ZN(new_n855));
  AOI211_X1 g430(.A(KEYINPUT104), .B(new_n696), .C1(new_n851), .C2(new_n853), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n741), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n858), .A3(new_n697), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n696), .B1(new_n851), .B2(new_n853), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n859), .B(new_n740), .C1(new_n860), .C2(new_n848), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n495), .A2(G130), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n501), .A2(G142), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n476), .A2(G118), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n862), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n632), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n857), .A2(new_n861), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n867), .B1(new_n857), .B2(new_n861), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n837), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n857), .A2(new_n861), .ZN(new_n872));
  INV_X1    g447(.A(new_n867), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n874), .A2(new_n836), .A3(new_n868), .ZN(new_n875));
  INV_X1    g450(.A(G37), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g453(.A(new_n827), .B(KEYINPUT105), .ZN(new_n879));
  INV_X1    g454(.A(new_n616), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n606), .A2(G299), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n600), .A2(new_n611), .A3(new_n605), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(KEYINPUT106), .A3(new_n883), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n881), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n884), .B(KEYINPUT41), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(new_n881), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT42), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n596), .B(KEYINPUT107), .Z(new_n892));
  AND2_X1   g467(.A1(new_n892), .A2(G288), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(G288), .ZN(new_n894));
  XNOR2_X1  g469(.A(G166), .B(G305), .ZN(new_n895));
  OR3_X1    g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n893), .B2(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n888), .B(new_n900), .C1(new_n889), .C2(new_n881), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n891), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n899), .B1(new_n891), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(G868), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n819), .A2(new_n617), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(G295));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n905), .ZN(G331));
  INV_X1    g482(.A(new_n882), .ZN(new_n908));
  INV_X1    g483(.A(new_n883), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(G286), .B(G171), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n827), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n825), .A2(new_n911), .A3(new_n826), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(KEYINPUT109), .A3(new_n914), .ZN(new_n915));
  OR3_X1    g490(.A1(new_n827), .A2(KEYINPUT109), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n918), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n913), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n910), .A2(new_n917), .B1(new_n921), .B2(new_n889), .ZN(new_n922));
  AOI21_X1  g497(.A(G37), .B1(new_n922), .B2(new_n898), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n898), .B2(new_n922), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n925));
  INV_X1    g500(.A(new_n889), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n886), .A2(new_n887), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  OAI22_X1  g503(.A1(new_n926), .A2(new_n917), .B1(new_n921), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n899), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n917), .A2(new_n910), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n921), .A2(new_n889), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n898), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n876), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n925), .B1(KEYINPUT43), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n935), .A2(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(KEYINPUT110), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n923), .A2(new_n938), .A3(new_n930), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n939), .A3(KEYINPUT43), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT111), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n937), .A2(new_n939), .A3(new_n942), .A4(KEYINPUT43), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n936), .B1(new_n945), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT45), .B1(new_n520), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  OAI211_X1 g524(.A(G40), .B(new_n487), .C1(new_n474), .C2(new_n477), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n740), .B(new_n743), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT112), .ZN(new_n953));
  INV_X1    g528(.A(G2067), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n761), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n839), .A2(G2067), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n708), .B(G1996), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G1986), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n596), .B(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n951), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT123), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n524), .B2(new_n947), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n520), .A2(new_n964), .A3(new_n947), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n478), .A2(new_n966), .A3(G40), .A4(new_n487), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n965), .A2(new_n967), .A3(G2084), .ZN(new_n968));
  INV_X1    g543(.A(new_n797), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n950), .A2(new_n948), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n515), .A2(new_n522), .A3(new_n519), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n522), .B1(new_n515), .B2(new_n519), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT45), .B(new_n947), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n969), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n963), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n950), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n976), .A3(new_n949), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n797), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n947), .B1(new_n971), .B2(new_n972), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n980));
  AOI211_X1 g555(.A(KEYINPUT50), .B(G1384), .C1(new_n515), .C2(new_n519), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n950), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n713), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n978), .A2(KEYINPUT123), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G8), .ZN(new_n985));
  NOR2_X1   g560(.A1(G168), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n975), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT124), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT124), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n975), .A2(new_n984), .A3(new_n989), .A4(new_n986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n978), .A2(KEYINPUT123), .A3(new_n983), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT123), .B1(new_n978), .B2(new_n983), .ZN(new_n993));
  OAI21_X1  g568(.A(G168), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT125), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n995), .B2(KEYINPUT51), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n995), .B2(KEYINPUT51), .ZN(new_n997));
  OAI21_X1  g572(.A(G8), .B1(new_n968), .B2(new_n974), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n986), .A2(KEYINPUT51), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n994), .A2(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n991), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT62), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n979), .A2(new_n1004), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n1004), .B(G1384), .C1(new_n515), .C2(new_n519), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n950), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1971), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G2090), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n964), .B(new_n947), .C1(new_n971), .C2(new_n972), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n520), .A2(new_n947), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1012));
  AND4_X1   g587(.A1(new_n1009), .A2(new_n1010), .A3(new_n976), .A4(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(G8), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G166), .A2(new_n985), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(G166), .B2(new_n985), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1014), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n980), .A2(new_n982), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(G2090), .ZN(new_n1024));
  OAI211_X1 g599(.A(G8), .B(new_n1020), .C1(new_n1024), .C2(new_n1008), .ZN(new_n1025));
  OAI21_X1  g600(.A(G8), .B1(new_n950), .B2(new_n1011), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G305), .A2(G1981), .ZN(new_n1027));
  INV_X1    g602(.A(G1981), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n587), .A2(new_n588), .A3(new_n1028), .A4(new_n589), .ZN(new_n1029));
  OR2_X1    g604(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1027), .A2(KEYINPUT115), .A3(new_n1029), .A4(KEYINPUT49), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n578), .A2(G1976), .A3(new_n580), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1036), .B(G8), .C1(new_n950), .C2(new_n1011), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n721), .B2(G1976), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n1026), .A2(new_n1035), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1037), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(new_n1038), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1040), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1022), .A2(new_n1025), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G2078), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1005), .A2(new_n1047), .A3(new_n1007), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1048), .A2(new_n1049), .B1(new_n1023), .B2(new_n793), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n970), .A2(KEYINPUT53), .A3(new_n973), .A4(new_n1047), .ZN(new_n1051));
  AOI21_X1  g626(.A(G301), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT62), .B1(new_n991), .B2(new_n1000), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1003), .A2(new_n1046), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n985), .B(G286), .C1(new_n978), .C2(new_n983), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1022), .A2(new_n1025), .A3(new_n1055), .A4(new_n1045), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT116), .B(KEYINPUT63), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT63), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n998), .A2(new_n1059), .A3(G286), .ZN(new_n1060));
  OAI21_X1  g635(.A(G8), .B1(new_n1024), .B2(new_n1008), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1021), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1060), .A2(new_n1025), .A3(new_n1045), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1025), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1026), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1035), .A2(new_n1026), .ZN(new_n1067));
  OR2_X1    g642(.A1(G288), .A2(G1976), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1029), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1065), .A2(new_n1045), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1064), .A2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT126), .B(KEYINPUT54), .Z(new_n1072));
  NAND4_X1  g647(.A1(new_n487), .A2(KEYINPUT53), .A3(G40), .A4(new_n1047), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(G2105), .B2(new_n473), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1006), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n949), .A3(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1050), .A2(G301), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1072), .B1(new_n1077), .B2(new_n1052), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1050), .A2(new_n1076), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G171), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1050), .A2(new_n1051), .A3(G301), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(KEYINPUT54), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1078), .A2(new_n1082), .A3(new_n1046), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1001), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1348), .B1(new_n980), .B2(new_n982), .ZN(new_n1086));
  OR3_X1    g661(.A1(new_n950), .A2(G2067), .A3(new_n1011), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n773), .B1(new_n965), .B2(new_n967), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(KEYINPUT118), .A3(new_n1087), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n1091), .A3(new_n607), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT119), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1089), .A2(new_n1091), .A3(new_n1094), .A4(new_n607), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n1096));
  AND3_X1   g671(.A1(G299), .A2(new_n1096), .A3(KEYINPUT57), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT57), .B1(G299), .B2(new_n1096), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT56), .B(G2072), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1005), .A2(new_n1007), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n950), .B1(KEYINPUT50), .B2(new_n1011), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1956), .B1(new_n1103), .B2(new_n1010), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1100), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1093), .A2(new_n1095), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1010), .A2(new_n976), .A3(new_n1012), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n803), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1005), .A2(new_n1007), .A3(new_n1101), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1099), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1086), .A2(new_n1088), .A3(new_n1085), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT118), .B1(new_n1090), .B2(new_n1087), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1089), .A2(new_n1091), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n607), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1110), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1099), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT61), .B1(new_n1119), .B2(KEYINPUT122), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1105), .B(new_n1110), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1117), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT120), .B(G1996), .Z(new_n1129));
  NAND3_X1  g704(.A1(new_n1005), .A2(new_n1007), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n950), .A2(new_n1011), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  AOI22_X1  g708(.A1(new_n1130), .A2(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1005), .A2(KEYINPUT121), .A3(new_n1007), .A4(new_n1129), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1128), .B1(new_n1136), .B2(new_n559), .ZN(new_n1137));
  AOI211_X1 g712(.A(KEYINPUT59), .B(new_n824), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1138));
  OAI22_X1  g713(.A1(new_n1137), .A2(new_n1138), .B1(new_n1114), .B2(new_n607), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1111), .B1(new_n1127), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1071), .B1(new_n1084), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1054), .B1(new_n1141), .B2(KEYINPUT127), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1143), .B(new_n1071), .C1(new_n1084), .C2(new_n1140), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n962), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n951), .A2(new_n960), .A3(new_n596), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT48), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1149));
  AOI211_X1 g724(.A(new_n1148), .B(new_n1149), .C1(new_n959), .C2(new_n951), .ZN(new_n1150));
  INV_X1    g725(.A(new_n957), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n951), .B1(new_n1151), .B2(new_n838), .ZN(new_n1152));
  INV_X1    g727(.A(G1996), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n951), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(KEYINPUT46), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1154), .A2(KEYINPUT46), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1152), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n1157), .B(KEYINPUT47), .Z(new_n1158));
  NAND2_X1  g733(.A1(new_n958), .A2(new_n957), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n741), .A2(new_n743), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n955), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g736(.A(new_n1150), .B(new_n1158), .C1(new_n951), .C2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1145), .A2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g738(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1165));
  NAND3_X1  g739(.A1(new_n877), .A2(new_n935), .A3(new_n1165), .ZN(G225));
  INV_X1    g740(.A(G225), .ZN(G308));
endmodule


