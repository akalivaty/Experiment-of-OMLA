//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  NAND2_X1  g005(.A1(G229gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(G1gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT16), .ZN(new_n209));
  INV_X1    g008(.A(G15gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G22gat), .ZN(new_n211));
  INV_X1    g010(.A(G22gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G15gat), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(G1gat), .B1(new_n211), .B2(new_n213), .ZN(new_n215));
  OAI21_X1  g014(.A(G8gat), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n217));
  INV_X1    g016(.A(G8gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n217), .B(new_n218), .C1(G1gat), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT17), .ZN(new_n222));
  INV_X1    g021(.A(G50gat), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT15), .B1(new_n223), .B2(G43gat), .ZN(new_n224));
  INV_X1    g023(.A(G43gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(G50gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT91), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G29gat), .A2(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT90), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT90), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(G29gat), .A3(G36gat), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n223), .A2(G43gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n225), .A2(G50gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT91), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .A4(KEYINPUT15), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT14), .ZN(new_n237));
  INV_X1    g036(.A(G29gat), .ZN(new_n238));
  INV_X1    g037(.A(G36gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n227), .A2(new_n232), .A3(new_n236), .A4(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT92), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n225), .B2(G50gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n223), .A2(KEYINPUT92), .A3(G43gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n234), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT15), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n224), .A2(new_n226), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT89), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n240), .A2(new_n253), .ZN(new_n254));
  NOR3_X1   g053(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT89), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n256), .A3(new_n241), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n252), .B1(new_n257), .B2(new_n232), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n222), .B1(new_n250), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT93), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n221), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT17), .B1(new_n221), .B2(new_n260), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n242), .A2(new_n231), .A3(new_n229), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n236), .A4(new_n227), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n241), .B1(new_n255), .B2(KEYINPUT89), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n240), .A2(new_n253), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n232), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n251), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g070(.A(KEYINPUT18), .B(new_n207), .C1(new_n261), .C2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT94), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n221), .ZN(new_n274));
  INV_X1    g073(.A(new_n221), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(new_n269), .A3(new_n265), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n207), .B(KEYINPUT13), .Z(new_n278));
  AOI21_X1  g077(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n278), .ZN(new_n280));
  AOI211_X1 g079(.A(KEYINPUT94), .B(new_n280), .C1(new_n274), .C2(new_n276), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n272), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n207), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT17), .B1(new_n265), .B2(new_n269), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n275), .B1(new_n284), .B2(KEYINPUT93), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n262), .A2(new_n270), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n283), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(KEYINPUT18), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n206), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n207), .B1(new_n261), .B2(new_n271), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT18), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n250), .A2(new_n221), .A3(new_n258), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n265), .A2(new_n269), .B1(new_n216), .B2(new_n220), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n278), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT94), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n273), .A3(new_n278), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n206), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n292), .A2(new_n298), .A3(new_n299), .A4(new_n272), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n289), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n303));
  XOR2_X1   g102(.A(G211gat), .B(G218gat), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT22), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n306), .A2(new_n307), .B1(G211gat), .B2(G218gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n306), .B2(new_n307), .ZN(new_n309));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n305), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n303), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G155gat), .B(G162gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G141gat), .B(G148gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(KEYINPUT2), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  INV_X1    g120(.A(G162gat), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT2), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT77), .ZN(new_n324));
  XOR2_X1   g123(.A(G141gat), .B(G148gat), .Z(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n317), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n320), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT78), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT2), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n317), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n323), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n326), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n316), .A2(new_n328), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n313), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(KEYINPUT75), .A3(new_n311), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n315), .B(new_n320), .C1(new_n324), .C2(new_n326), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n303), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(new_n312), .B2(new_n313), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G228gat), .A2(G233gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n337), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n345), .B(KEYINPUT80), .Z(new_n349));
  AOI21_X1  g148(.A(new_n334), .B1(new_n314), .B2(new_n315), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n350), .A2(KEYINPUT81), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n344), .B1(new_n350), .B2(KEYINPUT81), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT82), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT82), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n355), .B(new_n349), .C1(new_n351), .C2(new_n352), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n348), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G78gat), .B(G106gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT31), .B(G50gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(new_n212), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n212), .A2(KEYINPUT83), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n363), .B2(new_n360), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n357), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n367));
  INV_X1    g166(.A(G226gat), .ZN(new_n368));
  INV_X1    g167(.A(G233gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT27), .B(G183gat), .ZN(new_n371));
  INV_X1    g170(.A(G190gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n373), .A2(KEYINPUT28), .ZN(new_n374));
  NAND2_X1  g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(new_n373), .B2(KEYINPUT28), .ZN(new_n377));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT66), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n380), .B1(KEYINPUT26), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n384), .B(KEYINPUT68), .Z(new_n385));
  OAI211_X1 g184(.A(new_n374), .B(new_n377), .C1(new_n383), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT23), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n381), .B(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n376), .B1(KEYINPUT67), .B2(KEYINPUT24), .ZN(new_n389));
  INV_X1    g188(.A(G183gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n372), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n376), .A2(KEYINPUT67), .A3(KEYINPUT24), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n380), .B(new_n388), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT25), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT25), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n388), .A2(new_n396), .A3(new_n380), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n376), .A2(KEYINPUT65), .A3(KEYINPUT24), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT65), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT24), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n375), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n400), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n398), .A2(new_n391), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n395), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n370), .B1(new_n405), .B2(new_n303), .ZN(new_n406));
  INV_X1    g205(.A(new_n370), .ZN(new_n407));
  AOI22_X1  g206(.A1(KEYINPUT25), .A2(new_n394), .B1(new_n397), .B2(new_n403), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(new_n386), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n367), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n339), .A2(new_n343), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT29), .B1(new_n408), .B2(new_n386), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT76), .B1(new_n412), .B2(new_n370), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n406), .A2(new_n409), .ZN(new_n415));
  INV_X1    g214(.A(new_n411), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G8gat), .B(G36gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n414), .A2(new_n417), .A3(new_n421), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(KEYINPUT30), .A3(new_n424), .ZN(new_n425));
  OR3_X1    g224(.A1(new_n418), .A2(KEYINPUT30), .A3(new_n422), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G1gat), .B(G29gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT0), .ZN(new_n429));
  XNOR2_X1  g228(.A(G57gat), .B(G85gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G225gat), .A2(G233gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT70), .B(G120gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(G113gat), .ZN(new_n435));
  INV_X1    g234(.A(G113gat), .ZN(new_n436));
  INV_X1    g235(.A(G120gat), .ZN(new_n437));
  INV_X1    g236(.A(G134gat), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n436), .A2(new_n437), .B1(new_n438), .B2(G127gat), .ZN(new_n439));
  OR2_X1    g238(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n440));
  INV_X1    g239(.A(G127gat), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n441), .A2(G134gat), .B1(KEYINPUT71), .B2(KEYINPUT1), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n435), .A2(new_n439), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT1), .B1(new_n436), .B2(new_n437), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(new_n436), .B2(new_n437), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT69), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n441), .B2(G134gat), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(G127gat), .B2(new_n438), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n446), .A2(new_n441), .A3(G134gat), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n327), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT4), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n336), .A2(new_n328), .A3(KEYINPUT3), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n451), .A3(new_n340), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n433), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT39), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n432), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n336), .A2(new_n328), .A3(new_n451), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n443), .A2(new_n450), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n334), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n433), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT39), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n459), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT40), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n454), .A2(new_n456), .A3(KEYINPUT5), .A4(new_n433), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n454), .A2(new_n456), .A3(new_n433), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n433), .B1(new_n460), .B2(new_n462), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT5), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n432), .B(new_n468), .C1(new_n469), .C2(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n459), .B(KEYINPUT40), .C1(new_n457), .C2(new_n464), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n467), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n366), .B1(new_n427), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT37), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n415), .B2(new_n411), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n410), .A2(new_n416), .A3(new_n413), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n414), .A2(new_n417), .A3(new_n477), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n422), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT85), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n482), .A2(new_n483), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n454), .A2(new_n456), .ZN(new_n490));
  INV_X1    g289(.A(new_n433), .ZN(new_n491));
  OAI22_X1  g290(.A1(new_n490), .A2(new_n491), .B1(new_n470), .B2(new_n471), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n492), .A2(KEYINPUT6), .A3(new_n432), .A4(new_n468), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n473), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n432), .B1(new_n492), .B2(new_n468), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n424), .B(new_n493), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n483), .A2(new_n485), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n499), .A2(KEYINPUT87), .A3(new_n482), .A4(new_n486), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n489), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n421), .B1(new_n418), .B2(KEYINPUT37), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n502), .A2(KEYINPUT88), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n418), .A2(KEYINPUT37), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n502), .B2(KEYINPUT88), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n484), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n476), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n354), .A2(new_n356), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n365), .B1(new_n508), .B2(new_n347), .ZN(new_n509));
  AOI211_X1 g308(.A(new_n364), .B(new_n348), .C1(new_n354), .C2(new_n356), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n468), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n431), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n513), .A2(KEYINPUT79), .A3(new_n494), .A4(new_n473), .ZN(new_n514));
  INV_X1    g313(.A(new_n473), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT79), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n425), .A2(new_n426), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n511), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n405), .A2(new_n461), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n408), .A2(new_n451), .A3(new_n386), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT73), .ZN(new_n524));
  NAND2_X1  g323(.A1(G227gat), .A2(G233gat), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n525), .B(KEYINPUT64), .Z(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(KEYINPUT34), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n523), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n524), .B1(new_n523), .B2(new_n527), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n523), .A2(new_n525), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT34), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G43gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT72), .ZN(new_n535));
  XOR2_X1   g334(.A(G71gat), .B(G99gat), .Z(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n526), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT33), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(KEYINPUT32), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n538), .B(KEYINPUT32), .C1(new_n539), .C2(new_n537), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n533), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n530), .A2(new_n532), .A3(new_n542), .A4(new_n543), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT36), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT36), .B1(new_n545), .B2(new_n546), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT84), .B1(new_n520), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n549), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n547), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT84), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n514), .A2(new_n517), .B1(new_n425), .B2(new_n426), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(new_n511), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n507), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n518), .A2(new_n519), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n533), .A2(new_n544), .ZN(new_n559));
  INV_X1    g358(.A(new_n546), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n511), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT35), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n513), .A2(new_n494), .A3(new_n473), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT35), .B1(new_n564), .B2(new_n493), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n565), .A2(new_n519), .A3(new_n561), .A4(new_n511), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n302), .B1(new_n557), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT99), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT99), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n574), .A3(new_n569), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G85gat), .ZN(new_n577));
  INV_X1    g376(.A(G92gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(KEYINPUT8), .A2(new_n569), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n577), .B2(new_n578), .ZN(new_n581));
  NAND4_X1  g380(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n582), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT98), .A2(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n587), .A2(new_n572), .A3(new_n575), .A4(new_n579), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n270), .A2(new_n589), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n270), .A2(new_n222), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n259), .A2(new_n588), .A3(new_n584), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G190gat), .B(G218gat), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n598), .A2(KEYINPUT101), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(KEYINPUT101), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G134gat), .B(G162gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n597), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n604), .B1(new_n597), .B2(new_n599), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n609));
  AND2_X1   g408(.A1(G57gat), .A2(G64gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(G57gat), .A2(G64gat), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G57gat), .ZN(new_n613));
  INV_X1    g412(.A(G64gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G57gat), .A2(G64gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(KEYINPUT95), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(G71gat), .ZN(new_n619));
  INV_X1    g418(.A(G78gat), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(KEYINPUT9), .ZN(new_n621));
  NAND2_X1  g420(.A1(G71gat), .A2(G78gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n610), .A2(new_n611), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT9), .ZN(new_n625));
  XNOR2_X1  g424(.A(G71gat), .B(G78gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n618), .A2(new_n623), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(KEYINPUT21), .ZN(new_n629));
  XNOR2_X1  g428(.A(G127gat), .B(G155gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n221), .B1(KEYINPUT21), .B2(new_n628), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT97), .ZN(new_n635));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT96), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n635), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G183gat), .B(G211gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n633), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n608), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n576), .A2(new_n583), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n587), .A2(new_n579), .B1(new_n572), .B2(new_n575), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n628), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n612), .A2(new_n617), .B1(new_n622), .B2(new_n621), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n626), .B1(new_n624), .B2(KEYINPUT9), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n584), .B(new_n588), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n589), .A2(KEYINPUT10), .A3(new_n628), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n644), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n647), .A2(new_n650), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n655), .B2(new_n644), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  OR2_X1    g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n642), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n568), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n518), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT102), .B(G1gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1324gat));
  NOR2_X1   g466(.A1(new_n664), .A2(new_n519), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n218), .B2(new_n668), .ZN(new_n671));
  MUX2_X1   g470(.A(new_n670), .B(new_n671), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n664), .B2(new_n553), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n561), .A2(new_n210), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n664), .B2(new_n674), .ZN(G1326gat));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n664), .B2(new_n511), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n568), .A2(KEYINPUT103), .A3(new_n366), .A4(new_n663), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(new_n641), .ZN(new_n682));
  INV_X1    g481(.A(new_n662), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n608), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n568), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n518), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n238), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT45), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n557), .A2(new_n567), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n608), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n520), .A2(new_n550), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n507), .A2(new_n694), .B1(new_n563), .B2(new_n566), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n691), .B1(new_n695), .B2(new_n608), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n289), .A2(KEYINPUT104), .A3(new_n300), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT104), .B1(new_n289), .B2(new_n300), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n684), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n697), .A2(new_n687), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n689), .B1(new_n238), .B2(new_n703), .ZN(G1328gat));
  NOR2_X1   g503(.A1(new_n519), .A2(G36gat), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n690), .A2(new_n301), .A3(new_n685), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT105), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT106), .B1(new_n707), .B2(KEYINPUT46), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n706), .A2(KEYINPUT105), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(KEYINPUT105), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n709), .A2(new_n710), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n697), .A2(new_n427), .A3(new_n702), .ZN(new_n715));
  AOI22_X1  g514(.A1(KEYINPUT46), .A2(new_n707), .B1(new_n715), .B2(G36gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1329gat));
  NAND4_X1  g516(.A1(new_n693), .A2(new_n696), .A3(new_n550), .A4(new_n702), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n225), .B1(new_n718), .B2(KEYINPUT108), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT108), .B2(new_n718), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n686), .A2(new_n225), .A3(new_n561), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(KEYINPUT47), .A3(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n723));
  INV_X1    g522(.A(new_n721), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n718), .A2(G43gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n726), .ZN(G1330gat));
  NOR2_X1   g526(.A1(KEYINPUT109), .A2(KEYINPUT48), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n511), .A2(G50gat), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n686), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n693), .A2(new_n696), .A3(new_n366), .A4(new_n702), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G50gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(KEYINPUT109), .A2(KEYINPUT48), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1331gat));
  NOR2_X1   g534(.A1(new_n642), .A2(new_n700), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n662), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n695), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n687), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n738), .B(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n519), .ZN(new_n743));
  NOR2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  AND2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n743), .B2(new_n744), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n742), .B2(new_n553), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n738), .A2(new_n619), .A3(new_n561), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(KEYINPUT50), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1334gat));
  NOR2_X1   g553(.A1(new_n742), .A2(new_n511), .ZN(new_n755));
  XNOR2_X1  g554(.A(KEYINPUT111), .B(G78gat), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n755), .B(new_n756), .Z(G1335gat));
  NOR2_X1   g556(.A1(new_n700), .A2(new_n641), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n683), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n697), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(new_n687), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n695), .A2(new_n763), .A3(new_n608), .A4(new_n759), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n507), .A2(new_n694), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n608), .B1(new_n767), .B2(new_n567), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT51), .B1(new_n768), .B2(new_n758), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n764), .B2(new_n765), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n687), .A2(new_n577), .A3(new_n662), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n762), .A2(new_n577), .B1(new_n773), .B2(new_n774), .ZN(G1336gat));
  NOR3_X1   g574(.A1(new_n519), .A2(G92gat), .A3(new_n683), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n771), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n693), .A2(new_n696), .A3(new_n427), .A4(new_n760), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n776), .B1(new_n769), .B2(new_n764), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n782), .B1(new_n784), .B2(KEYINPUT52), .ZN(new_n785));
  AOI211_X1 g584(.A(KEYINPUT113), .B(new_n778), .C1(new_n780), .C2(new_n783), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n781), .B1(new_n785), .B2(new_n786), .ZN(G1337gat));
  AND2_X1   g586(.A1(new_n761), .A2(new_n550), .ZN(new_n788));
  INV_X1    g587(.A(G99gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n561), .A2(new_n789), .A3(new_n662), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n788), .A2(new_n789), .B1(new_n773), .B2(new_n790), .ZN(G1338gat));
  NOR3_X1   g590(.A1(new_n511), .A2(G106gat), .A3(new_n683), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n771), .A2(new_n772), .A3(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n693), .A2(new_n696), .A3(new_n366), .A4(new_n760), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G106gat), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n769), .A2(new_n764), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n798), .A2(new_n792), .B1(G106gat), .B2(new_n794), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n793), .A2(new_n797), .B1(new_n799), .B2(new_n796), .ZN(G1339gat));
  INV_X1    g599(.A(KEYINPUT104), .ZN(new_n801));
  AOI22_X1  g600(.A1(KEYINPUT18), .A2(new_n287), .B1(new_n296), .B2(new_n297), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n299), .B1(new_n802), .B2(new_n292), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n282), .A2(new_n288), .A3(new_n206), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n652), .A2(new_n653), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n643), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n652), .A2(new_n653), .A3(new_n644), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(KEYINPUT54), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n659), .B1(new_n654), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n809), .A2(new_n811), .A3(KEYINPUT114), .A4(KEYINPUT55), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n814), .A2(new_n661), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n289), .A2(KEYINPUT104), .A3(new_n300), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n809), .A2(new_n811), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(KEYINPUT115), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n805), .A2(new_n816), .A3(new_n817), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n285), .A2(new_n286), .A3(new_n283), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n278), .B2(new_n277), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n826), .A2(new_n827), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n205), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(new_n300), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n662), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n607), .B1(new_n825), .B2(new_n833), .ZN(new_n834));
  AND4_X1   g633(.A1(new_n607), .A2(new_n832), .A3(new_n816), .A4(new_n824), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT117), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n814), .A2(new_n661), .A3(new_n815), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n822), .B2(new_n823), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n607), .A3(new_n832), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n662), .A2(new_n831), .A3(new_n300), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(new_n700), .B2(new_n839), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n837), .B(new_n840), .C1(new_n842), .C2(new_n607), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n836), .A2(new_n843), .A3(new_n682), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n736), .A2(new_n683), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n518), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n562), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n519), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n700), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n366), .B1(new_n844), .B2(new_n845), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n561), .B1(new_n851), .B2(KEYINPUT118), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n853), .B(new_n366), .C1(new_n844), .C2(new_n845), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n687), .A2(new_n519), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n302), .A2(new_n436), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n850), .B1(new_n857), .B2(new_n858), .ZN(G1340gat));
  OR3_X1    g658(.A1(new_n848), .A2(new_n434), .A3(new_n683), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n855), .A2(new_n683), .A3(new_n856), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n437), .ZN(G1341gat));
  NAND3_X1  g661(.A1(new_n849), .A2(new_n441), .A3(new_n641), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n855), .A2(new_n682), .A3(new_n856), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n441), .ZN(G1342gat));
  INV_X1    g664(.A(new_n846), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n847), .A2(new_n438), .A3(new_n519), .A4(new_n607), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT56), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n855), .A2(new_n608), .A3(new_n856), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n438), .ZN(G1343gat));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n550), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n816), .A2(new_n301), .A3(new_n820), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n607), .B1(new_n833), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n682), .B1(new_n874), .B2(new_n835), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n511), .B1(new_n875), .B2(new_n845), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n511), .B1(new_n844), .B2(new_n845), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n877), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G141gat), .B1(new_n881), .B2(new_n302), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n846), .A2(KEYINPUT119), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n553), .A2(new_n366), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n846), .B2(KEYINPUT119), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n302), .A2(G141gat), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT120), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n883), .A2(new_n885), .A3(new_n519), .A4(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n882), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G141gat), .B1(new_n881), .B2(new_n701), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(new_n888), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n892), .B2(new_n889), .ZN(G1344gat));
  NOR2_X1   g692(.A1(new_n683), .A2(G148gat), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n883), .A2(new_n885), .A3(new_n519), .A4(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  INV_X1    g695(.A(new_n875), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n642), .A2(new_n301), .A3(new_n662), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n877), .B(new_n366), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n856), .A2(new_n550), .A3(new_n683), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n899), .B(new_n900), .C1(new_n879), .C2(new_n877), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n896), .B1(new_n901), .B2(G148gat), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n896), .A2(G148gat), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n903), .B1(new_n880), .B2(new_n662), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n895), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT121), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n907), .B(new_n895), .C1(new_n902), .C2(new_n904), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1345gat));
  NAND2_X1  g708(.A1(new_n883), .A2(new_n885), .ZN(new_n910));
  NOR4_X1   g709(.A1(new_n910), .A2(G155gat), .A3(new_n427), .A4(new_n682), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n321), .B1(new_n880), .B2(new_n641), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n911), .A2(new_n912), .ZN(G1346gat));
  OAI21_X1  g712(.A(G162gat), .B1(new_n881), .B2(new_n608), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n519), .A2(new_n322), .A3(new_n607), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n910), .B2(new_n915), .ZN(G1347gat));
  NAND2_X1  g715(.A1(new_n427), .A2(new_n518), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n852), .A2(new_n854), .A3(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(G169gat), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n918), .A2(new_n919), .A3(new_n302), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n687), .B1(new_n844), .B2(new_n845), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(new_n427), .A3(new_n847), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n700), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n920), .A2(new_n923), .ZN(G1348gat));
  OAI21_X1  g723(.A(G176gat), .B1(new_n918), .B2(new_n683), .ZN(new_n925));
  INV_X1    g724(.A(G176gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n922), .A2(new_n926), .A3(new_n662), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1349gat));
  AND2_X1   g727(.A1(new_n641), .A2(new_n371), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT122), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  NOR4_X1   g729(.A1(new_n852), .A2(new_n854), .A3(new_n682), .A4(new_n917), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n390), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n934), .B(new_n930), .C1(new_n931), .C2(new_n390), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n922), .A2(new_n372), .A3(new_n607), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n937), .B(new_n938), .ZN(new_n939));
  OAI211_X1 g738(.A(KEYINPUT61), .B(G190gat), .C1(new_n918), .C2(new_n608), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n941));
  NOR4_X1   g740(.A1(new_n852), .A2(new_n854), .A3(new_n608), .A4(new_n917), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n372), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n939), .A2(new_n940), .A3(new_n943), .ZN(G1351gat));
  NAND4_X1  g743(.A1(new_n921), .A2(new_n427), .A3(new_n366), .A4(new_n553), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(new_n701), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n553), .A2(new_n518), .A3(new_n427), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT124), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n899), .B(new_n948), .C1(new_n879), .C2(new_n877), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n301), .A2(G197gat), .ZN(new_n950));
  OAI22_X1  g749(.A1(new_n946), .A2(G197gat), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(G1352gat));
  OR3_X1    g751(.A1(new_n945), .A2(G204gat), .A3(new_n683), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  OAI21_X1  g753(.A(G204gat), .B1(new_n949), .B2(new_n683), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(G1353gat));
  NOR2_X1   g756(.A1(new_n947), .A2(new_n682), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n899), .B(new_n958), .C1(new_n879), .C2(new_n877), .ZN(new_n959));
  OAI21_X1  g758(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n945), .A2(G211gat), .A3(new_n682), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n959), .B(new_n961), .C1(new_n963), .C2(new_n964), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n966), .A2(new_n967), .A3(KEYINPUT126), .A4(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1354gat));
  NOR2_X1   g772(.A1(new_n945), .A2(new_n608), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n607), .A2(G218gat), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT127), .ZN(new_n976));
  OAI22_X1  g775(.A1(new_n974), .A2(G218gat), .B1(new_n949), .B2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(G1355gat));
endmodule


