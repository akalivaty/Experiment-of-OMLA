//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164, new_n1165;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  AOI22_X1  g035(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT72), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT72), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  OR2_X1    g045(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(G137), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n464), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT73), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g051(.A(KEYINPUT73), .B(new_n464), .C1(new_n470), .C2(new_n473), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n472), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G125), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n467), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT71), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n467), .A2(G2104), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n469), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n483), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(G113), .A2(G2104), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n482), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n478), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G160));
  OAI21_X1  g070(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G112), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n482), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n499));
  INV_X1    g074(.A(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G136), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n503), .B(KEYINPUT74), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n482), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI211_X1 g081(.A(new_n498), .B(new_n504), .C1(G124), .C2(new_n506), .ZN(G162));
  OR2_X1    g082(.A1(new_n500), .A2(G114), .ZN(new_n508));
  OAI21_X1  g083(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(G126), .A2(G2105), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n470), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n471), .A2(new_n514), .A3(G138), .A4(new_n472), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n489), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n488), .B1(new_n469), .B2(new_n487), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n471), .A2(G138), .A3(new_n472), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT4), .B1(new_n470), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n513), .B1(new_n519), .B2(new_n521), .ZN(G164));
  XNOR2_X1  g097(.A(KEYINPUT5), .B(G543), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n523), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT6), .B(G651), .Z(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(G166));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT6), .B(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT75), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n532), .A2(G543), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT5), .B(G543), .Z(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n528), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n536), .A2(new_n543), .ZN(G168));
  NAND2_X1  g119(.A1(new_n535), .A2(G52), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n525), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n538), .A2(G90), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(new_n535), .A2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n537), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(G651), .B1(new_n538), .B2(G81), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n532), .A2(G543), .A3(new_n534), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n563), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n537), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(new_n538), .B2(G91), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n535), .A2(KEYINPUT76), .A3(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n573), .A2(KEYINPUT9), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n535), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT77), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n538), .A2(G87), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n580), .A2(KEYINPUT77), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n579), .A2(new_n581), .A3(new_n582), .A4(new_n583), .ZN(G288));
  AOI22_X1  g159(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n525), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n523), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n528), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n538), .A2(G85), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n591), .B1(new_n525), .B2(new_n592), .C1(new_n565), .C2(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NOR2_X1   g170(.A1(G301), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n538), .A2(G92), .ZN(new_n597));
  XOR2_X1   g172(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n598));
  XOR2_X1   g173(.A(new_n597), .B(new_n598), .Z(new_n599));
  INV_X1    g174(.A(G54), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n565), .A2(new_n600), .B1(new_n525), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(KEYINPUT80), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(KEYINPUT80), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n596), .B1(new_n611), .B2(new_n595), .ZN(G284));
  AOI21_X1  g187(.A(new_n596), .B1(new_n611), .B2(new_n595), .ZN(G321));
  NOR2_X1   g188(.A1(G286), .A2(new_n595), .ZN(new_n614));
  AND2_X1   g189(.A1(new_n572), .A2(new_n575), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT81), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n614), .B1(new_n616), .B2(new_n595), .ZN(G280));
  XNOR2_X1  g192(.A(G280), .B(KEYINPUT82), .ZN(G297));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n611), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n556), .A2(new_n595), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n610), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n595), .ZN(G323));
  XNOR2_X1  g198(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n624));
  XNOR2_X1  g199(.A(G323), .B(new_n624), .ZN(G282));
  NAND2_X1  g200(.A1(new_n486), .A2(new_n489), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n463), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n627), .B(new_n628), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  OAI221_X1 g208(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n481), .C2(G111), .ZN(new_n634));
  INV_X1    g209(.A(G135), .ZN(new_n635));
  INV_X1    g210(.A(G123), .ZN(new_n636));
  OAI221_X1 g211(.A(new_n634), .B1(new_n501), .B2(new_n635), .C1(new_n636), .C2(new_n505), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND3_X1  g213(.A1(new_n632), .A2(new_n633), .A3(new_n638), .ZN(G156));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT86), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n641), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT85), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2430), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n644), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  AND3_X1   g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(G401));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT87), .ZN(new_n658));
  NOR2_X1   g233(.A1(G2072), .A2(G2078), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n442), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n658), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n658), .A2(new_n660), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n660), .B(KEYINPUT17), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n662), .C1(new_n658), .C2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n658), .A3(new_n661), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n664), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n676), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT20), .Z(new_n680));
  AOI211_X1 g255(.A(new_n678), .B(new_n680), .C1(new_n673), .C2(new_n677), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G35), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G162), .B2(new_n688), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT29), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G2090), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G20), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT23), .Z(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G299), .B2(G16), .ZN(new_n696));
  INV_X1    g271(.A(G1956), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n693), .A2(G19), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n557), .B2(new_n693), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1341), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n688), .A2(G26), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  OAI221_X1 g278(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n481), .C2(G116), .ZN(new_n704));
  INV_X1    g279(.A(G128), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n505), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G140), .B2(new_n502), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n703), .B1(new_n707), .B2(new_n688), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G2067), .ZN(new_n709));
  NOR4_X1   g284(.A1(new_n692), .A2(new_n698), .A3(new_n701), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n688), .A2(G32), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n502), .A2(G141), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT26), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n715), .A2(new_n716), .B1(G105), .B2(new_n463), .ZN(new_n717));
  INV_X1    g292(.A(G129), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n505), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n711), .B1(new_n720), .B2(new_n688), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT27), .B(G1996), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n688), .A2(G27), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G164), .B2(new_n688), .ZN(new_n724));
  OAI22_X1  g299(.A1(new_n721), .A2(new_n722), .B1(G2078), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT31), .B(G11), .Z(new_n726));
  INV_X1    g301(.A(G28), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT96), .Z(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n727), .B2(KEYINPUT30), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n693), .A2(G21), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G286), .B2(G16), .ZN(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n731), .B1(new_n688), .B2(new_n637), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G2078), .B2(new_n724), .ZN(new_n736));
  NOR2_X1   g311(.A1(G171), .A2(new_n693), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G5), .B2(new_n693), .ZN(new_n738));
  INV_X1    g313(.A(G1961), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n738), .A2(new_n739), .B1(new_n734), .B2(new_n733), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n736), .B(new_n740), .C1(new_n739), .C2(new_n738), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n725), .B(new_n741), .C1(new_n721), .C2(new_n722), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n688), .A2(G33), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n626), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(new_n481), .ZN(new_n745));
  INV_X1    g320(.A(G139), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n501), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT25), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n745), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT94), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n743), .B1(new_n752), .B2(new_n688), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(G2072), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT24), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(G34), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(G34), .ZN(new_n757));
  AOI21_X1  g332(.A(G29), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n494), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT95), .B(G2084), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n753), .A2(G2072), .ZN(new_n762));
  AND3_X1   g337(.A1(new_n754), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n742), .A2(KEYINPUT97), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G4), .A2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT93), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n610), .B2(new_n693), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1348), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n710), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(KEYINPUT97), .B1(new_n742), .B2(new_n763), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n693), .A2(G22), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G166), .B2(new_n693), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1971), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT33), .B(G1976), .ZN(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G23), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT92), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G288), .B2(new_n693), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n774), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G6), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n589), .B2(G16), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(G1981), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n778), .A2(new_n775), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(G1981), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n779), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT91), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT34), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n502), .A2(G131), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n506), .A2(G119), .ZN(new_n792));
  NOR2_X1   g367(.A1(G95), .A2(G2105), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT88), .Z(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(G2104), .C1(G107), .C2(new_n481), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n791), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT89), .Z(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(new_n688), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G25), .B2(new_n688), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT35), .B(G1991), .Z(new_n800));
  AND2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n693), .A2(G24), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT90), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G290), .B2(G16), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(G1986), .Z(new_n806));
  NOR3_X1   g381(.A1(new_n801), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n789), .A2(new_n790), .A3(new_n807), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT36), .Z(new_n809));
  NOR2_X1   g384(.A1(new_n771), .A2(new_n809), .ZN(G311));
  OR2_X1    g385(.A1(new_n771), .A2(new_n809), .ZN(G150));
  NOR2_X1   g386(.A1(new_n610), .A2(new_n619), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n816), .A2(new_n817), .A3(new_n525), .ZN(new_n818));
  INV_X1    g393(.A(G55), .ZN(new_n819));
  INV_X1    g394(.A(new_n538), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT100), .B(G93), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n565), .A2(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n556), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n814), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n827));
  AOI21_X1  g402(.A(G860), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  INV_X1    g404(.A(new_n823), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G860), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT37), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n832), .ZN(G145));
  INV_X1    g408(.A(KEYINPUT105), .ZN(new_n834));
  INV_X1    g409(.A(new_n512), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n499), .A2(new_n835), .B1(new_n508), .B2(new_n510), .ZN(new_n836));
  INV_X1    g411(.A(new_n520), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n514), .B1(new_n499), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n515), .B1(new_n486), .B2(new_n489), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT101), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n836), .B(new_n842), .C1(new_n838), .C2(new_n839), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n720), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n752), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n707), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n752), .B(new_n720), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n849), .A2(new_n707), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n844), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  OAI221_X1 g426(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n481), .C2(G118), .ZN(new_n852));
  INV_X1    g427(.A(G130), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n505), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G142), .B2(new_n502), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n629), .B(new_n855), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n796), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n849), .A2(new_n707), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n846), .A2(new_n847), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n860), .A2(new_n861), .A3(new_n841), .A4(new_n843), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n851), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n494), .B(new_n637), .ZN(new_n864));
  XOR2_X1   g439(.A(G162), .B(new_n864), .Z(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n859), .B1(new_n851), .B2(new_n862), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n863), .B(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n834), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n851), .A2(new_n862), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT104), .B1(new_n872), .B2(new_n859), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n851), .A2(new_n859), .A3(new_n862), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n874), .A2(new_n865), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n867), .A2(new_n868), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n873), .A2(new_n875), .A3(KEYINPUT105), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n865), .B1(new_n874), .B2(new_n867), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT40), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n884));
  AOI211_X1 g459(.A(new_n884), .B(new_n881), .C1(new_n871), .C2(new_n877), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(new_n885), .ZN(G395));
  INV_X1    g461(.A(KEYINPUT106), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n606), .B1(new_n887), .B2(G299), .ZN(new_n888));
  NAND2_X1  g463(.A1(G299), .A2(new_n887), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n606), .A2(new_n615), .A3(KEYINPUT106), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT41), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n615), .A2(KEYINPUT106), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n606), .A3(new_n889), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(KEYINPUT108), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n900), .B(KEYINPUT41), .C1(new_n891), .C2(new_n892), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n622), .A2(new_n825), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n824), .B1(new_n610), .B2(G559), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT109), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n891), .B2(new_n892), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n894), .A2(new_n896), .A3(KEYINPUT107), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n902), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT42), .ZN(new_n916));
  XNOR2_X1  g491(.A(G166), .B(KEYINPUT110), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(G288), .ZN(new_n918));
  XNOR2_X1  g493(.A(G290), .B(G305), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n918), .B(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n907), .A2(new_n921), .A3(new_n912), .A4(new_n914), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n916), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n920), .B1(new_n916), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n830), .A2(new_n595), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(G295));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n926), .ZN(G331));
  NAND2_X1  g503(.A1(new_n824), .A2(G301), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n830), .A2(new_n556), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n823), .A2(new_n557), .ZN(new_n931));
  OAI21_X1  g506(.A(G171), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n929), .A2(new_n932), .A3(G168), .ZN(new_n933));
  AOI21_X1  g508(.A(G168), .B1(new_n929), .B2(new_n932), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n899), .A2(new_n935), .A3(new_n901), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n894), .B(new_n896), .C1(new_n933), .C2(new_n934), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n920), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n938), .A2(G37), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n920), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT43), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n935), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n920), .B1(new_n942), .B2(new_n911), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n935), .A2(new_n893), .A3(new_n898), .ZN(new_n944));
  AOI21_X1  g519(.A(G37), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n945), .A2(KEYINPUT43), .A3(new_n940), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT44), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(new_n939), .B2(new_n940), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n945), .A2(new_n949), .A3(new_n940), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n947), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n947), .B2(new_n952), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(G397));
  INV_X1    g531(.A(KEYINPUT117), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n478), .A2(G40), .A3(new_n493), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n478), .A2(KEYINPUT112), .A3(G40), .A4(new_n493), .ZN(new_n961));
  INV_X1    g536(.A(G1384), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n840), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1976), .ZN(new_n966));
  OR2_X1    g541(.A1(G288), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(G8), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT52), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT52), .B1(G288), .B2(new_n966), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n965), .A2(new_n967), .A3(G8), .A4(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1981), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n589), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(G1981), .B1(new_n586), .B2(new_n588), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n973), .A2(KEYINPUT49), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT49), .B1(new_n973), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n965), .A3(G8), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n969), .A2(new_n971), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n981));
  INV_X1    g556(.A(G8), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(G166), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n840), .A2(new_n986), .A3(new_n962), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n960), .A2(new_n961), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G2090), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n841), .A2(KEYINPUT45), .A3(new_n962), .A4(new_n843), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n963), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n990), .A2(new_n960), .A3(new_n961), .A4(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1971), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n988), .A2(new_n989), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n984), .B1(new_n995), .B2(new_n982), .ZN(new_n996));
  INV_X1    g571(.A(G2084), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n960), .A2(new_n997), .A3(new_n961), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n985), .A2(new_n987), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n963), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n840), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n960), .A2(new_n992), .A3(new_n961), .A4(new_n1003), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n998), .A2(new_n1002), .B1(new_n1004), .B2(new_n734), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1005), .A2(new_n982), .A3(G286), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n960), .A2(new_n961), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(new_n1002), .A3(new_n989), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n993), .A2(new_n994), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n980), .A2(new_n983), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT114), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(G8), .A3(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n979), .A2(new_n996), .A3(new_n1006), .A4(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT116), .B(KEYINPUT63), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n998), .A2(new_n1002), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1004), .A2(new_n734), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AND4_X1   g594(.A1(KEYINPUT63), .A2(new_n1019), .A3(G8), .A4(G168), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1010), .A2(G8), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n984), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1020), .A2(new_n1022), .A3(new_n1013), .A4(new_n979), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n969), .A2(new_n971), .A3(new_n978), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G288), .A2(G1976), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT115), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1027), .A2(new_n978), .B1(new_n972), .B2(new_n589), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n965), .A2(G8), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1013), .A2(new_n1025), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n957), .B1(new_n1024), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g607(.A(KEYINPUT117), .B(new_n1030), .C1(new_n1016), .C2(new_n1023), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1007), .A2(new_n1002), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n739), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n991), .B1(new_n844), .B2(G1384), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n958), .A2(new_n1038), .A3(G2078), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n990), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT123), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n993), .B2(G2078), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1037), .A2(new_n1039), .A3(KEYINPUT123), .A4(new_n990), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1036), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(G171), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OR3_X1    g622(.A1(new_n1004), .A2(new_n1038), .A3(G2078), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1036), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1043), .A2(G301), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT54), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT124), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1051), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1046), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1057), .B(G8), .C1(new_n1019), .C2(G286), .ZN(new_n1058));
  NOR2_X1   g633(.A1(G168), .A2(new_n982), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(KEYINPUT51), .B(new_n1060), .C1(new_n1005), .C2(new_n982), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n1019), .B2(new_n1059), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1005), .A2(KEYINPUT121), .A3(new_n1060), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1058), .B(new_n1061), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT122), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1019), .A2(new_n1062), .A3(new_n1059), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT121), .B1(new_n1005), .B2(new_n1060), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n1061), .A4(new_n1058), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n979), .A2(new_n996), .A3(new_n1013), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1043), .ZN(new_n1074));
  OAI21_X1  g649(.A(G171), .B1(new_n1049), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1036), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(new_n1050), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1073), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1056), .A2(new_n1072), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n572), .B2(new_n575), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n960), .A2(new_n961), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n985), .A2(new_n987), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n697), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT56), .B(G2072), .Z(new_n1089));
  OAI211_X1 g664(.A(new_n1085), .B(new_n1088), .C1(new_n993), .C2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n988), .A2(G1956), .B1(new_n993), .B2(new_n1089), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1090), .A2(new_n1093), .A3(KEYINPUT61), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT61), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1348), .ZN(new_n1097));
  INV_X1    g672(.A(G2067), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1098), .A2(new_n960), .A3(new_n961), .A4(new_n964), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1035), .A2(new_n1097), .B1(new_n1099), .B2(KEYINPUT118), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1099), .A2(KEYINPUT118), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n1101), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n606), .A3(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1100), .A2(new_n1101), .A3(KEYINPUT60), .A4(new_n607), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n993), .A2(G1996), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  AND2_X1   g684(.A1(new_n965), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n557), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT59), .B(new_n557), .C1(new_n1108), .C2(new_n1110), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1107), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1096), .A2(new_n1106), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n607), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1093), .B1(new_n1117), .B2(KEYINPUT119), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1102), .A2(KEYINPUT119), .A3(new_n606), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1090), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1081), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1080), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1116), .A2(new_n1081), .A3(new_n1120), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1034), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1066), .A2(new_n1125), .A3(new_n1071), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1072), .B2(KEYINPUT62), .ZN(new_n1130));
  AOI211_X1 g705(.A(KEYINPUT125), .B(new_n1125), .C1(new_n1066), .C2(new_n1071), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1128), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT126), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1128), .B(new_n1134), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1124), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1037), .A2(new_n1086), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n720), .B(G1996), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n707), .B(G2067), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n796), .B(new_n800), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(G290), .B(G1986), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1137), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1136), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1137), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1145), .A2(G1986), .A3(G290), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1149));
  AOI211_X1 g724(.A(new_n1148), .B(new_n1149), .C1(new_n1137), .C2(new_n1141), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1145), .A2(G1996), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT46), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1145), .B1(new_n720), .B2(new_n1139), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT47), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n797), .A2(new_n800), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1156), .A2(new_n1157), .B1(G2067), .B2(new_n847), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1150), .B(new_n1155), .C1(new_n1137), .C2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1144), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g735(.A1(new_n878), .A2(new_n882), .ZN(new_n1162));
  OR2_X1    g736(.A1(new_n950), .A2(new_n951), .ZN(new_n1163));
  INV_X1    g737(.A(G319), .ZN(new_n1164));
  NOR4_X1   g738(.A1(G229), .A2(new_n1164), .A3(G401), .A4(G227), .ZN(new_n1165));
  AND3_X1   g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1165), .ZN(G308));
  NAND3_X1  g740(.A1(new_n1162), .A2(new_n1163), .A3(new_n1165), .ZN(G225));
endmodule


