

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705;

  OR2_X1 U363 ( .A1(n669), .A2(G902), .ZN(n366) );
  NOR2_X1 U364 ( .A1(n701), .A2(n356), .ZN(n558) );
  XNOR2_X1 U365 ( .A(n457), .B(n458), .ZN(n586) );
  NOR2_X1 U366 ( .A1(n586), .A2(G902), .ZN(n352) );
  INV_X2 U367 ( .A(G953), .ZN(n692) );
  NOR2_X2 U368 ( .A1(n589), .A2(n674), .ZN(n591) );
  NOR2_X1 U369 ( .A1(n559), .A2(n629), .ZN(n556) );
  INV_X1 U370 ( .A(n567), .ZN(n638) );
  INV_X1 U371 ( .A(G146), .ZN(n392) );
  INV_X1 U372 ( .A(n456), .ZN(n457) );
  XNOR2_X1 U373 ( .A(n392), .B(G125), .ZN(n433) );
  INV_X1 U374 ( .A(G134), .ZN(n421) );
  NAND2_X1 U375 ( .A1(n381), .A2(n380), .ZN(n583) );
  NAND2_X1 U376 ( .A1(n556), .A2(n555), .ZN(n357) );
  XNOR2_X1 U377 ( .A(n521), .B(n505), .ZN(n544) );
  XNOR2_X1 U378 ( .A(n422), .B(n421), .ZN(n462) );
  XNOR2_X1 U379 ( .A(n408), .B(n407), .ZN(n453) );
  XNOR2_X1 U380 ( .A(n416), .B(G128), .ZN(n422) );
  XOR2_X1 U381 ( .A(KEYINPUT68), .B(G131), .Z(n484) );
  XNOR2_X2 U382 ( .A(n357), .B(KEYINPUT32), .ZN(n703) );
  XNOR2_X1 U383 ( .A(KEYINPUT4), .B(KEYINPUT67), .ZN(n689) );
  XNOR2_X1 U384 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n434) );
  XNOR2_X1 U385 ( .A(n462), .B(n423), .ZN(n687) );
  XNOR2_X1 U386 ( .A(n361), .B(n360), .ZN(n538) );
  INV_X1 U387 ( .A(KEYINPUT74), .ZN(n360) );
  OR2_X1 U388 ( .A1(n631), .A2(n632), .ZN(n361) );
  OR2_X1 U389 ( .A1(G902), .A2(G237), .ZN(n493) );
  XNOR2_X1 U390 ( .A(G902), .B(KEYINPUT15), .ZN(n576) );
  XNOR2_X1 U391 ( .A(n429), .B(n428), .ZN(n510) );
  XNOR2_X1 U392 ( .A(n433), .B(n391), .ZN(n688) );
  XNOR2_X1 U393 ( .A(G140), .B(KEYINPUT10), .ZN(n391) );
  NOR2_X2 U394 ( .A1(n544), .A2(n545), .ZN(n348) );
  INV_X1 U395 ( .A(G143), .ZN(n416) );
  XNOR2_X1 U396 ( .A(G116), .B(KEYINPUT3), .ZN(n407) );
  XOR2_X1 U397 ( .A(G113), .B(G119), .Z(n408) );
  XOR2_X1 U398 ( .A(KEYINPUT18), .B(KEYINPUT77), .Z(n414) );
  NAND2_X1 U399 ( .A1(n614), .A2(KEYINPUT80), .ZN(n398) );
  XNOR2_X1 U400 ( .A(n368), .B(n367), .ZN(n381) );
  INV_X1 U401 ( .A(n702), .ZN(n380) );
  INV_X1 U402 ( .A(KEYINPUT48), .ZN(n367) );
  XNOR2_X1 U403 ( .A(n378), .B(n377), .ZN(n432) );
  XNOR2_X1 U404 ( .A(G119), .B(KEYINPUT23), .ZN(n377) );
  XNOR2_X1 U405 ( .A(n379), .B(G137), .ZN(n378) );
  XNOR2_X1 U406 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n379) );
  XNOR2_X1 U407 ( .A(n473), .B(n472), .ZN(n668) );
  XNOR2_X1 U408 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U409 ( .A(n466), .B(n465), .ZN(n473) );
  XNOR2_X1 U410 ( .A(n489), .B(n490), .ZN(n666) );
  XNOR2_X1 U411 ( .A(G122), .B(G143), .ZN(n475) );
  XNOR2_X1 U412 ( .A(n363), .B(n687), .ZN(n456) );
  XNOR2_X1 U413 ( .A(n539), .B(KEYINPUT33), .ZN(n650) );
  NAND2_X1 U414 ( .A1(n538), .A2(n560), .ZN(n539) );
  XNOR2_X1 U415 ( .A(n395), .B(n534), .ZN(n627) );
  NAND2_X1 U416 ( .A1(n623), .A2(n621), .ZN(n395) );
  INV_X1 U417 ( .A(n538), .ZN(n564) );
  NAND2_X1 U418 ( .A1(n657), .A2(n576), .ZN(n419) );
  XNOR2_X1 U419 ( .A(n500), .B(KEYINPUT28), .ZN(n501) );
  XNOR2_X1 U420 ( .A(n552), .B(n551), .ZN(n559) );
  INV_X1 U421 ( .A(n668), .ZN(n385) );
  AND2_X2 U422 ( .A1(n663), .A2(n662), .ZN(n670) );
  INV_X1 U423 ( .A(KEYINPUT47), .ZN(n353) );
  NOR2_X1 U424 ( .A1(G953), .A2(G237), .ZN(n479) );
  XNOR2_X1 U425 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n450) );
  XOR2_X1 U426 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n451) );
  NAND2_X1 U427 ( .A1(n372), .A2(n369), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n369) );
  AND2_X1 U429 ( .A1(n373), .A2(n612), .ZN(n372) );
  INV_X1 U430 ( .A(KEYINPUT46), .ZN(n370) );
  XNOR2_X1 U431 ( .A(KEYINPUT105), .B(KEYINPUT104), .ZN(n461) );
  INV_X1 U432 ( .A(G122), .ZN(n463) );
  XNOR2_X1 U433 ( .A(G116), .B(G107), .ZN(n464) );
  XOR2_X1 U434 ( .A(G104), .B(G113), .Z(n476) );
  NOR2_X1 U435 ( .A1(n619), .A2(n617), .ZN(n623) );
  XNOR2_X1 U436 ( .A(n365), .B(n364), .ZN(n537) );
  INV_X1 U437 ( .A(KEYINPUT66), .ZN(n364) );
  AND2_X1 U438 ( .A1(n585), .A2(n615), .ZN(n663) );
  XNOR2_X1 U439 ( .A(n354), .B(n675), .ZN(n657) );
  XNOR2_X1 U440 ( .A(n418), .B(n349), .ZN(n354) );
  XNOR2_X1 U441 ( .A(n417), .B(n420), .ZN(n349) );
  NAND2_X1 U442 ( .A1(n396), .A2(n575), .ZN(n662) );
  NOR2_X1 U443 ( .A1(n583), .A2(n398), .ZN(n397) );
  NOR2_X1 U444 ( .A1(n569), .A2(n512), .ZN(n514) );
  XNOR2_X1 U445 ( .A(n504), .B(KEYINPUT76), .ZN(n505) );
  XNOR2_X1 U446 ( .A(n510), .B(n430), .ZN(n631) );
  XNOR2_X1 U447 ( .A(n406), .B(n405), .ZN(n531) );
  XNOR2_X1 U448 ( .A(n491), .B(G475), .ZN(n405) );
  OR2_X1 U449 ( .A1(n666), .A2(G902), .ZN(n406) );
  INV_X1 U450 ( .A(n583), .ZN(n577) );
  XNOR2_X1 U451 ( .A(n437), .B(n436), .ZN(n669) );
  XNOR2_X1 U452 ( .A(G128), .B(G110), .ZN(n431) );
  XNOR2_X1 U453 ( .A(n667), .B(n346), .ZN(n404) );
  XNOR2_X1 U454 ( .A(n456), .B(n362), .ZN(n661) );
  XNOR2_X1 U455 ( .A(n425), .B(n424), .ZN(n426) );
  INV_X1 U456 ( .A(G140), .ZN(n424) );
  INV_X1 U457 ( .A(KEYINPUT42), .ZN(n393) );
  NOR2_X1 U458 ( .A1(n627), .A2(n535), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n358), .B(KEYINPUT35), .ZN(n701) );
  XNOR2_X1 U460 ( .A(n546), .B(n345), .ZN(n359) );
  INV_X1 U461 ( .A(KEYINPUT120), .ZN(n382) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(G60) );
  INV_X1 U463 ( .A(KEYINPUT60), .ZN(n400) );
  NAND2_X1 U464 ( .A1(n403), .A2(n402), .ZN(n401) );
  XNOR2_X1 U465 ( .A(n665), .B(n404), .ZN(n403) );
  NOR2_X1 U466 ( .A1(n374), .A2(n674), .ZN(G54) );
  XNOR2_X1 U467 ( .A(n376), .B(n375), .ZN(n374) );
  XNOR2_X1 U468 ( .A(n661), .B(n660), .ZN(n375) );
  NAND2_X1 U469 ( .A1(n670), .A2(G469), .ZN(n376) );
  INV_X1 U470 ( .A(KEYINPUT56), .ZN(n387) );
  AND2_X1 U471 ( .A1(G221), .A2(n467), .ZN(n340) );
  XOR2_X1 U472 ( .A(n440), .B(KEYINPUT25), .Z(n341) );
  XOR2_X1 U473 ( .A(n547), .B(KEYINPUT78), .Z(n342) );
  AND2_X1 U474 ( .A1(G210), .A2(n493), .ZN(n343) );
  XOR2_X1 U475 ( .A(n659), .B(n658), .Z(n344) );
  XNOR2_X1 U476 ( .A(KEYINPUT34), .B(KEYINPUT79), .ZN(n345) );
  XNOR2_X1 U477 ( .A(KEYINPUT59), .B(KEYINPUT89), .ZN(n346) );
  NOR2_X1 U478 ( .A1(G952), .A2(n692), .ZN(n674) );
  INV_X1 U479 ( .A(n674), .ZN(n402) );
  NAND2_X1 U480 ( .A1(n347), .A2(n517), .ZN(n351) );
  XNOR2_X1 U481 ( .A(n602), .B(KEYINPUT84), .ZN(n347) );
  XNOR2_X1 U482 ( .A(n420), .B(G146), .ZN(n363) );
  XNOR2_X2 U483 ( .A(n348), .B(KEYINPUT0), .ZN(n566) );
  XNOR2_X1 U484 ( .A(n350), .B(KEYINPUT30), .ZN(n512) );
  NAND2_X1 U485 ( .A1(n638), .A2(n621), .ZN(n350) );
  XNOR2_X1 U486 ( .A(n351), .B(KEYINPUT81), .ZN(n518) );
  XNOR2_X2 U487 ( .A(n352), .B(n459), .ZN(n567) );
  XNOR2_X1 U488 ( .A(n603), .B(n353), .ZN(n508) );
  NOR2_X2 U489 ( .A1(n535), .A2(n544), .ZN(n603) );
  NAND2_X1 U490 ( .A1(n355), .A2(n397), .ZN(n396) );
  NAND2_X1 U491 ( .A1(n355), .A2(n584), .ZN(n615) );
  NAND2_X1 U492 ( .A1(n355), .A2(n692), .ZN(n680) );
  XNOR2_X2 U493 ( .A(n399), .B(KEYINPUT45), .ZN(n355) );
  NAND2_X1 U494 ( .A1(n703), .A2(n599), .ZN(n356) );
  NAND2_X1 U495 ( .A1(n359), .A2(n342), .ZN(n358) );
  XNOR2_X1 U496 ( .A(n426), .B(n427), .ZN(n362) );
  NAND2_X1 U497 ( .A1(n629), .A2(n628), .ZN(n365) );
  XNOR2_X2 U498 ( .A(n366), .B(n341), .ZN(n629) );
  NAND2_X1 U499 ( .A1(n699), .A2(n704), .ZN(n371) );
  XNOR2_X1 U500 ( .A(n520), .B(KEYINPUT73), .ZN(n373) );
  XNOR2_X1 U501 ( .A(n411), .B(n427), .ZN(n412) );
  XNOR2_X1 U502 ( .A(n383), .B(n382), .ZN(G63) );
  NAND2_X1 U503 ( .A1(n384), .A2(n402), .ZN(n383) );
  XNOR2_X1 U504 ( .A(n386), .B(n385), .ZN(n384) );
  NAND2_X1 U505 ( .A1(n670), .A2(G478), .ZN(n386) );
  XNOR2_X1 U506 ( .A(n388), .B(n387), .ZN(G51) );
  NAND2_X1 U507 ( .A1(n389), .A2(n402), .ZN(n388) );
  XNOR2_X1 U508 ( .A(n390), .B(n344), .ZN(n389) );
  NAND2_X1 U509 ( .A1(n670), .A2(G210), .ZN(n390) );
  XNOR2_X1 U510 ( .A(n394), .B(n393), .ZN(n704) );
  NAND2_X1 U511 ( .A1(n577), .A2(n614), .ZN(n691) );
  NAND2_X1 U512 ( .A1(n574), .A2(n573), .ZN(n399) );
  XNOR2_X1 U513 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U514 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U515 ( .A(n409), .B(G122), .ZN(n411) );
  XNOR2_X1 U516 ( .A(n484), .B(G137), .ZN(n423) );
  XNOR2_X1 U517 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U518 ( .A(n550), .B(KEYINPUT71), .ZN(n551) );
  XNOR2_X1 U519 ( .A(n688), .B(n340), .ZN(n436) );
  XNOR2_X1 U520 ( .A(n474), .B(G478), .ZN(n532) );
  XNOR2_X1 U521 ( .A(n586), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U522 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U523 ( .A(n530), .B(n529), .ZN(n699) );
  INV_X1 U524 ( .A(KEYINPUT80), .ZN(n578) );
  XNOR2_X1 U525 ( .A(G101), .B(n689), .ZN(n420) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(KEYINPUT72), .Z(n409) );
  XNOR2_X1 U527 ( .A(G107), .B(G110), .ZN(n410) );
  XNOR2_X1 U528 ( .A(n410), .B(G104), .ZN(n427) );
  XOR2_X2 U529 ( .A(n453), .B(n412), .Z(n675) );
  NAND2_X1 U530 ( .A1(G224), .A2(n692), .ZN(n413) );
  XNOR2_X1 U531 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U532 ( .A(n415), .B(KEYINPUT17), .Z(n418) );
  XNOR2_X1 U533 ( .A(n422), .B(n433), .ZN(n417) );
  XNOR2_X2 U534 ( .A(n419), .B(n343), .ZN(n503) );
  XOR2_X1 U535 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n496) );
  NAND2_X1 U536 ( .A1(G227), .A2(n692), .ZN(n425) );
  NOR2_X1 U537 ( .A1(G902), .A2(n661), .ZN(n429) );
  XNOR2_X1 U538 ( .A(KEYINPUT69), .B(G469), .ZN(n428) );
  INV_X1 U539 ( .A(KEYINPUT1), .ZN(n430) );
  INV_X1 U540 ( .A(n631), .ZN(n563) );
  XNOR2_X1 U541 ( .A(n432), .B(n431), .ZN(n437) );
  NAND2_X1 U542 ( .A1(n692), .A2(G234), .ZN(n435) );
  XNOR2_X1 U543 ( .A(n435), .B(n434), .ZN(n467) );
  XOR2_X1 U544 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n439) );
  NAND2_X1 U545 ( .A1(G234), .A2(n576), .ZN(n438) );
  XNOR2_X1 U546 ( .A(n439), .B(n438), .ZN(n447) );
  NAND2_X1 U547 ( .A1(n447), .A2(G217), .ZN(n440) );
  NAND2_X1 U548 ( .A1(G237), .A2(G234), .ZN(n441) );
  XNOR2_X1 U549 ( .A(n441), .B(KEYINPUT14), .ZN(n444) );
  NAND2_X1 U550 ( .A1(G952), .A2(n444), .ZN(n442) );
  XNOR2_X1 U551 ( .A(KEYINPUT90), .B(n442), .ZN(n648) );
  NOR2_X1 U552 ( .A1(n648), .A2(G953), .ZN(n443) );
  XNOR2_X1 U553 ( .A(n443), .B(KEYINPUT91), .ZN(n542) );
  NAND2_X1 U554 ( .A1(G902), .A2(n444), .ZN(n540) );
  NOR2_X1 U555 ( .A1(G900), .A2(n540), .ZN(n445) );
  NAND2_X1 U556 ( .A1(G953), .A2(n445), .ZN(n446) );
  NAND2_X1 U557 ( .A1(n542), .A2(n446), .ZN(n513) );
  NAND2_X1 U558 ( .A1(n447), .A2(G221), .ZN(n448) );
  XOR2_X1 U559 ( .A(KEYINPUT21), .B(n448), .Z(n628) );
  NAND2_X1 U560 ( .A1(n513), .A2(n628), .ZN(n449) );
  NOR2_X1 U561 ( .A1(n629), .A2(n449), .ZN(n499) );
  XNOR2_X1 U562 ( .A(KEYINPUT70), .B(G472), .ZN(n459) );
  XNOR2_X1 U563 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U564 ( .A(n453), .B(n452), .Z(n455) );
  NAND2_X1 U565 ( .A1(n479), .A2(G210), .ZN(n454) );
  XNOR2_X1 U566 ( .A(n455), .B(n454), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n567), .B(KEYINPUT107), .ZN(n460) );
  XNOR2_X1 U568 ( .A(n460), .B(KEYINPUT6), .ZN(n554) );
  INV_X1 U569 ( .A(n554), .ZN(n560) );
  XNOR2_X1 U570 ( .A(n462), .B(n461), .ZN(n466) );
  NAND2_X1 U571 ( .A1(G217), .A2(n467), .ZN(n471) );
  XOR2_X1 U572 ( .A(KEYINPUT9), .B(KEYINPUT106), .Z(n469) );
  XNOR2_X1 U573 ( .A(KEYINPUT7), .B(KEYINPUT103), .ZN(n468) );
  XNOR2_X1 U574 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U575 ( .A1(n668), .A2(G902), .ZN(n474) );
  INV_X1 U576 ( .A(n532), .ZN(n506) );
  XNOR2_X1 U577 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n491) );
  XNOR2_X1 U578 ( .A(n476), .B(n475), .ZN(n490) );
  INV_X1 U579 ( .A(n688), .ZN(n488) );
  XOR2_X1 U580 ( .A(KEYINPUT99), .B(KEYINPUT97), .Z(n478) );
  XNOR2_X1 U581 ( .A(KEYINPUT98), .B(KEYINPUT100), .ZN(n477) );
  XNOR2_X1 U582 ( .A(n478), .B(n477), .ZN(n483) );
  XOR2_X1 U583 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n481) );
  NAND2_X1 U584 ( .A1(n479), .A2(G214), .ZN(n480) );
  XNOR2_X1 U585 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U586 ( .A(n483), .B(n482), .ZN(n486) );
  XNOR2_X1 U587 ( .A(n484), .B(KEYINPUT12), .ZN(n485) );
  NOR2_X1 U588 ( .A1(n506), .A2(n531), .ZN(n605) );
  AND2_X1 U589 ( .A1(n560), .A2(n605), .ZN(n492) );
  NAND2_X1 U590 ( .A1(n499), .A2(n492), .ZN(n522) );
  NOR2_X1 U591 ( .A1(n563), .A2(n522), .ZN(n494) );
  NAND2_X1 U592 ( .A1(G214), .A2(n493), .ZN(n621) );
  NAND2_X1 U593 ( .A1(n494), .A2(n621), .ZN(n495) );
  XNOR2_X1 U594 ( .A(n496), .B(n495), .ZN(n497) );
  NOR2_X1 U595 ( .A1(n503), .A2(n497), .ZN(n498) );
  XOR2_X1 U596 ( .A(KEYINPUT111), .B(n498), .Z(n702) );
  AND2_X1 U597 ( .A1(n638), .A2(n499), .ZN(n500) );
  NAND2_X1 U598 ( .A1(n501), .A2(n510), .ZN(n502) );
  XNOR2_X1 U599 ( .A(n502), .B(KEYINPUT112), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n503), .A2(n621), .ZN(n521) );
  XNOR2_X1 U601 ( .A(KEYINPUT19), .B(KEYINPUT65), .ZN(n504) );
  AND2_X1 U602 ( .A1(n506), .A2(n531), .ZN(n607) );
  NOR2_X1 U603 ( .A1(n605), .A2(n607), .ZN(n618) );
  XOR2_X1 U604 ( .A(KEYINPUT83), .B(n618), .Z(n571) );
  NAND2_X1 U605 ( .A1(n603), .A2(n571), .ZN(n507) );
  NAND2_X1 U606 ( .A1(n508), .A2(n507), .ZN(n519) );
  NAND2_X1 U607 ( .A1(KEYINPUT47), .A2(n618), .ZN(n509) );
  XNOR2_X1 U608 ( .A(KEYINPUT82), .B(n509), .ZN(n517) );
  NAND2_X1 U609 ( .A1(n537), .A2(n510), .ZN(n511) );
  XNOR2_X1 U610 ( .A(n511), .B(KEYINPUT94), .ZN(n569) );
  NAND2_X1 U611 ( .A1(n514), .A2(n513), .ZN(n525) );
  NOR2_X1 U612 ( .A1(n532), .A2(n531), .ZN(n515) );
  XNOR2_X1 U613 ( .A(n515), .B(KEYINPUT109), .ZN(n547) );
  NOR2_X1 U614 ( .A1(n525), .A2(n547), .ZN(n516) );
  NAND2_X1 U615 ( .A1(n503), .A2(n516), .ZN(n602) );
  NAND2_X1 U616 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U617 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U618 ( .A(KEYINPUT36), .B(n523), .ZN(n524) );
  XNOR2_X1 U619 ( .A(KEYINPUT88), .B(n563), .ZN(n553) );
  NAND2_X1 U620 ( .A1(n524), .A2(n553), .ZN(n612) );
  INV_X1 U621 ( .A(n525), .ZN(n527) );
  XNOR2_X1 U622 ( .A(n503), .B(KEYINPUT38), .ZN(n617) );
  INV_X1 U623 ( .A(n617), .ZN(n526) );
  NAND2_X1 U624 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U625 ( .A(n528), .B(KEYINPUT39), .ZN(n536) );
  NAND2_X1 U626 ( .A1(n536), .A2(n605), .ZN(n530) );
  XOR2_X1 U627 ( .A(KEYINPUT113), .B(KEYINPUT40), .Z(n529) );
  NAND2_X1 U628 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U629 ( .A(n533), .B(KEYINPUT108), .ZN(n619) );
  INV_X1 U630 ( .A(KEYINPUT41), .ZN(n534) );
  NAND2_X1 U631 ( .A1(n536), .A2(n607), .ZN(n614) );
  INV_X1 U632 ( .A(n537), .ZN(n632) );
  INV_X1 U633 ( .A(n540), .ZN(n541) );
  NOR2_X1 U634 ( .A1(G898), .A2(n692), .ZN(n677) );
  NAND2_X1 U635 ( .A1(n541), .A2(n677), .ZN(n543) );
  AND2_X1 U636 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U637 ( .A1(n650), .A2(n566), .ZN(n546) );
  INV_X1 U638 ( .A(n628), .ZN(n548) );
  NOR2_X1 U639 ( .A1(n548), .A2(n619), .ZN(n549) );
  NAND2_X1 U640 ( .A1(n549), .A2(n566), .ZN(n552) );
  XOR2_X1 U641 ( .A(KEYINPUT64), .B(KEYINPUT22), .Z(n550) );
  AND2_X1 U642 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U643 ( .A1(n556), .A2(n631), .ZN(n557) );
  NAND2_X1 U644 ( .A1(n567), .A2(n557), .ZN(n599) );
  XNOR2_X1 U645 ( .A(n558), .B(KEYINPUT44), .ZN(n574) );
  NOR2_X1 U646 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U647 ( .A1(n561), .A2(n629), .ZN(n562) );
  NOR2_X1 U648 ( .A1(n563), .A2(n562), .ZN(n592) );
  NOR2_X1 U649 ( .A1(n567), .A2(n564), .ZN(n640) );
  NAND2_X1 U650 ( .A1(n566), .A2(n640), .ZN(n565) );
  XNOR2_X1 U651 ( .A(n565), .B(KEYINPUT31), .ZN(n608) );
  NAND2_X1 U652 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U653 ( .A1(n569), .A2(n568), .ZN(n595) );
  NOR2_X1 U654 ( .A1(n608), .A2(n595), .ZN(n570) );
  NOR2_X1 U655 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U656 ( .A1(n592), .A2(n572), .ZN(n573) );
  INV_X1 U657 ( .A(KEYINPUT2), .ZN(n575) );
  INV_X1 U658 ( .A(n576), .ZN(n585) );
  NAND2_X1 U659 ( .A1(n578), .A2(n614), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n614), .A2(KEYINPUT2), .ZN(n579) );
  NAND2_X1 U661 ( .A1(n579), .A2(KEYINPUT80), .ZN(n580) );
  NAND2_X1 U662 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U663 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U664 ( .A1(n670), .A2(G472), .ZN(n588) );
  XNOR2_X1 U665 ( .A(KEYINPUT63), .B(KEYINPUT87), .ZN(n590) );
  XNOR2_X1 U666 ( .A(n591), .B(n590), .ZN(G57) );
  XOR2_X1 U667 ( .A(G101), .B(n592), .Z(G3) );
  NAND2_X1 U668 ( .A1(n595), .A2(n605), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n593), .B(KEYINPUT114), .ZN(n594) );
  XNOR2_X1 U670 ( .A(G104), .B(n594), .ZN(G6) );
  XOR2_X1 U671 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n597) );
  NAND2_X1 U672 ( .A1(n595), .A2(n607), .ZN(n596) );
  XNOR2_X1 U673 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X1 U674 ( .A(G107), .B(n598), .ZN(G9) );
  XNOR2_X1 U675 ( .A(G110), .B(n599), .ZN(G12) );
  XOR2_X1 U676 ( .A(G128), .B(KEYINPUT29), .Z(n601) );
  NAND2_X1 U677 ( .A1(n607), .A2(n603), .ZN(n600) );
  XNOR2_X1 U678 ( .A(n601), .B(n600), .ZN(G30) );
  XNOR2_X1 U679 ( .A(G143), .B(n602), .ZN(G45) );
  NAND2_X1 U680 ( .A1(n603), .A2(n605), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n604), .B(G146), .ZN(G48) );
  NAND2_X1 U682 ( .A1(n608), .A2(n605), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n606), .B(G113), .ZN(G15) );
  NAND2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(G116), .ZN(G18) );
  XOR2_X1 U686 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n611) );
  XNOR2_X1 U687 ( .A(G125), .B(KEYINPUT37), .ZN(n610) );
  XNOR2_X1 U688 ( .A(n611), .B(n610), .ZN(n613) );
  XOR2_X1 U689 ( .A(n613), .B(n612), .Z(G27) );
  XNOR2_X1 U690 ( .A(G134), .B(n614), .ZN(G36) );
  NAND2_X1 U691 ( .A1(n662), .A2(n615), .ZN(n616) );
  XNOR2_X1 U692 ( .A(KEYINPUT86), .B(n616), .ZN(n654) );
  OR2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n625) );
  INV_X1 U696 ( .A(n623), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U698 ( .A1(n626), .A2(n650), .ZN(n645) );
  INV_X1 U699 ( .A(n627), .ZN(n649) );
  NOR2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U701 ( .A(KEYINPUT49), .B(n630), .ZN(n636) );
  XOR2_X1 U702 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n634) );
  NAND2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U706 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U707 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U708 ( .A(n641), .B(KEYINPUT118), .ZN(n642) );
  XNOR2_X1 U709 ( .A(n642), .B(KEYINPUT51), .ZN(n643) );
  NAND2_X1 U710 ( .A1(n649), .A2(n643), .ZN(n644) );
  NAND2_X1 U711 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U712 ( .A(KEYINPUT52), .B(n646), .Z(n647) );
  NOR2_X1 U713 ( .A1(n648), .A2(n647), .ZN(n652) );
  AND2_X1 U714 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U715 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U716 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U717 ( .A1(n655), .A2(G953), .ZN(n656) );
  XNOR2_X1 U718 ( .A(n656), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U719 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n659) );
  XNOR2_X1 U720 ( .A(n657), .B(KEYINPUT55), .ZN(n658) );
  XOR2_X1 U721 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n660) );
  AND2_X1 U722 ( .A1(n662), .A2(G475), .ZN(n664) );
  NAND2_X1 U723 ( .A1(n664), .A2(n663), .ZN(n665) );
  INV_X1 U724 ( .A(n666), .ZN(n667) );
  XOR2_X1 U725 ( .A(n669), .B(KEYINPUT121), .Z(n672) );
  NAND2_X1 U726 ( .A1(n670), .A2(G217), .ZN(n671) );
  XNOR2_X1 U727 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U728 ( .A1(n674), .A2(n673), .ZN(G66) );
  XOR2_X1 U729 ( .A(n675), .B(G101), .Z(n676) );
  NOR2_X1 U730 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U731 ( .A(KEYINPUT124), .B(n678), .Z(n679) );
  XNOR2_X1 U732 ( .A(KEYINPUT123), .B(n679), .ZN(n686) );
  XNOR2_X1 U733 ( .A(n680), .B(KEYINPUT122), .ZN(n684) );
  NAND2_X1 U734 ( .A1(G953), .A2(G224), .ZN(n681) );
  XNOR2_X1 U735 ( .A(KEYINPUT61), .B(n681), .ZN(n682) );
  NAND2_X1 U736 ( .A1(n682), .A2(G898), .ZN(n683) );
  NAND2_X1 U737 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U738 ( .A(n686), .B(n685), .ZN(G69) );
  XNOR2_X1 U739 ( .A(n688), .B(n687), .ZN(n690) );
  XNOR2_X1 U740 ( .A(n689), .B(n690), .ZN(n694) );
  XNOR2_X1 U741 ( .A(n694), .B(n691), .ZN(n693) );
  NAND2_X1 U742 ( .A1(n693), .A2(n692), .ZN(n698) );
  XNOR2_X1 U743 ( .A(G227), .B(n694), .ZN(n695) );
  NAND2_X1 U744 ( .A1(n695), .A2(G900), .ZN(n696) );
  NAND2_X1 U745 ( .A1(G953), .A2(n696), .ZN(n697) );
  NAND2_X1 U746 ( .A1(n698), .A2(n697), .ZN(G72) );
  XNOR2_X1 U747 ( .A(G131), .B(n699), .ZN(n700) );
  XNOR2_X1 U748 ( .A(n700), .B(KEYINPUT126), .ZN(G33) );
  XOR2_X1 U749 ( .A(n701), .B(G122), .Z(G24) );
  XOR2_X1 U750 ( .A(G140), .B(n702), .Z(G42) );
  XNOR2_X1 U751 ( .A(n703), .B(G119), .ZN(G21) );
  XOR2_X1 U752 ( .A(G137), .B(n704), .Z(n705) );
  XNOR2_X1 U753 ( .A(KEYINPUT125), .B(n705), .ZN(G39) );
endmodule

