

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n806), .A2(n753), .ZN(n519) );
  XOR2_X1 U553 ( .A(KEYINPUT105), .B(n739), .Z(n520) );
  INV_X1 U554 ( .A(KEYINPUT101), .ZN(n696) );
  XNOR2_X1 U555 ( .A(KEYINPUT31), .B(KEYINPUT103), .ZN(n728) );
  XNOR2_X1 U556 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U557 ( .A1(n731), .A2(n730), .ZN(n742) );
  NAND2_X1 U558 ( .A1(G160), .A2(G40), .ZN(n758) );
  AND2_X1 U559 ( .A1(n538), .A2(G2104), .ZN(n886) );
  NOR2_X1 U560 ( .A1(n642), .A2(G651), .ZN(n649) );
  XNOR2_X1 U561 ( .A(KEYINPUT65), .B(KEYINPUT23), .ZN(n536) );
  XNOR2_X1 U562 ( .A(n537), .B(n536), .ZN(n540) );
  NOR2_X1 U563 ( .A1(n548), .A2(n547), .ZN(G160) );
  INV_X1 U564 ( .A(G651), .ZN(n527) );
  XOR2_X1 U565 ( .A(KEYINPUT0), .B(G543), .Z(n642) );
  OR2_X1 U566 ( .A1(n527), .A2(n642), .ZN(n521) );
  XNOR2_X1 U567 ( .A(KEYINPUT69), .B(n521), .ZN(n652) );
  NAND2_X1 U568 ( .A1(n652), .A2(G76), .ZN(n522) );
  XNOR2_X1 U569 ( .A(KEYINPUT78), .B(n522), .ZN(n525) );
  NOR2_X1 U570 ( .A1(G543), .A2(G651), .ZN(n648) );
  NAND2_X1 U571 ( .A1(n648), .A2(G89), .ZN(n523) );
  XNOR2_X1 U572 ( .A(KEYINPUT4), .B(n523), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U574 ( .A(n526), .B(KEYINPUT5), .ZN(n533) );
  NOR2_X1 U575 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U576 ( .A(KEYINPUT1), .B(n528), .Z(n656) );
  NAND2_X1 U577 ( .A1(G63), .A2(n656), .ZN(n530) );
  NAND2_X1 U578 ( .A1(G51), .A2(n649), .ZN(n529) );
  NAND2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U580 ( .A(KEYINPUT6), .B(n531), .Z(n532) );
  NAND2_X1 U581 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U582 ( .A(n534), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U583 ( .A(G168), .B(KEYINPUT8), .ZN(n535) );
  XNOR2_X1 U584 ( .A(n535), .B(KEYINPUT79), .ZN(G286) );
  INV_X1 U585 ( .A(G2105), .ZN(n538) );
  NAND2_X1 U586 ( .A1(G101), .A2(n886), .ZN(n537) );
  NOR2_X1 U587 ( .A1(G2104), .A2(n538), .ZN(n881) );
  NAND2_X1 U588 ( .A1(G125), .A2(n881), .ZN(n539) );
  NAND2_X1 U589 ( .A1(n540), .A2(n539), .ZN(n548) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n880) );
  NAND2_X1 U591 ( .A1(n880), .A2(G113), .ZN(n541) );
  XNOR2_X1 U592 ( .A(n541), .B(KEYINPUT66), .ZN(n545) );
  XNOR2_X1 U593 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n543) );
  NOR2_X1 U594 ( .A1(G2105), .A2(G2104), .ZN(n542) );
  XNOR2_X2 U595 ( .A(n543), .B(n542), .ZN(n884) );
  NAND2_X1 U596 ( .A1(G137), .A2(n884), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U598 ( .A(KEYINPUT68), .B(n546), .ZN(n547) );
  NAND2_X1 U599 ( .A1(G138), .A2(n884), .ZN(n550) );
  NAND2_X1 U600 ( .A1(G102), .A2(n886), .ZN(n549) );
  NAND2_X1 U601 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U602 ( .A(n551), .B(KEYINPUT93), .ZN(n556) );
  NAND2_X1 U603 ( .A1(G126), .A2(n881), .ZN(n554) );
  NAND2_X1 U604 ( .A1(G114), .A2(n880), .ZN(n552) );
  XNOR2_X1 U605 ( .A(KEYINPUT92), .B(n552), .ZN(n553) );
  AND2_X1 U606 ( .A1(n554), .A2(n553), .ZN(n555) );
  AND2_X1 U607 ( .A1(n556), .A2(n555), .ZN(G164) );
  NAND2_X1 U608 ( .A1(G91), .A2(n648), .ZN(n558) );
  NAND2_X1 U609 ( .A1(G78), .A2(n652), .ZN(n557) );
  NAND2_X1 U610 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U611 ( .A1(G65), .A2(n656), .ZN(n560) );
  NAND2_X1 U612 ( .A1(G53), .A2(n649), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n560), .A2(n559), .ZN(n561) );
  OR2_X1 U614 ( .A1(n562), .A2(n561), .ZN(G299) );
  NAND2_X1 U615 ( .A1(G64), .A2(n656), .ZN(n564) );
  NAND2_X1 U616 ( .A1(G52), .A2(n649), .ZN(n563) );
  NAND2_X1 U617 ( .A1(n564), .A2(n563), .ZN(n570) );
  NAND2_X1 U618 ( .A1(n652), .A2(G77), .ZN(n565) );
  XOR2_X1 U619 ( .A(KEYINPUT71), .B(n565), .Z(n567) );
  NAND2_X1 U620 ( .A1(n648), .A2(G90), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U622 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U623 ( .A1(n570), .A2(n569), .ZN(G171) );
  INV_X1 U624 ( .A(G132), .ZN(G219) );
  INV_X1 U625 ( .A(G82), .ZN(G220) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G69), .ZN(G235) );
  INV_X1 U628 ( .A(G108), .ZN(G238) );
  INV_X1 U629 ( .A(G120), .ZN(G236) );
  NAND2_X1 U630 ( .A1(G94), .A2(G452), .ZN(n571) );
  XOR2_X1 U631 ( .A(KEYINPUT72), .B(n571), .Z(G173) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U633 ( .A(n572), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U634 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n574) );
  INV_X1 U635 ( .A(G223), .ZN(n830) );
  NAND2_X1 U636 ( .A1(G567), .A2(n830), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT73), .B(n575), .Z(G234) );
  NAND2_X1 U639 ( .A1(n648), .A2(G81), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G68), .A2(n652), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT13), .B(n579), .Z(n583) );
  NAND2_X1 U644 ( .A1(G56), .A2(n656), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT14), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT75), .ZN(n582) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n649), .A2(G43), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n978) );
  INV_X1 U650 ( .A(G860), .ZN(n623) );
  OR2_X1 U651 ( .A1(n978), .A2(n623), .ZN(G153) );
  INV_X1 U652 ( .A(G171), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G868), .A2(G301), .ZN(n596) );
  NAND2_X1 U654 ( .A1(G54), .A2(n649), .ZN(n592) );
  NAND2_X1 U655 ( .A1(G92), .A2(n648), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G79), .A2(n652), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n656), .A2(G66), .ZN(n588) );
  XOR2_X1 U659 ( .A(KEYINPUT76), .B(n588), .Z(n589) );
  NOR2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U662 ( .A(n593), .B(KEYINPUT15), .ZN(n594) );
  XNOR2_X1 U663 ( .A(KEYINPUT77), .B(n594), .ZN(n975) );
  INV_X1 U664 ( .A(G868), .ZN(n669) );
  NAND2_X1 U665 ( .A1(n975), .A2(n669), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n596), .A2(n595), .ZN(G284) );
  NOR2_X1 U667 ( .A1(G286), .A2(n669), .ZN(n598) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U669 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n623), .A2(G559), .ZN(n599) );
  INV_X1 U671 ( .A(n975), .ZN(n899) );
  NAND2_X1 U672 ( .A1(n599), .A2(n899), .ZN(n600) );
  XNOR2_X1 U673 ( .A(n600), .B(KEYINPUT80), .ZN(n601) );
  XNOR2_X1 U674 ( .A(KEYINPUT16), .B(n601), .ZN(G148) );
  NOR2_X1 U675 ( .A1(G559), .A2(n669), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n899), .A2(n602), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT81), .ZN(n605) );
  NOR2_X1 U678 ( .A1(n978), .A2(G868), .ZN(n604) );
  NOR2_X1 U679 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G99), .A2(n886), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G111), .A2(n880), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U683 ( .A(KEYINPUT82), .B(n608), .ZN(n613) );
  NAND2_X1 U684 ( .A1(G123), .A2(n881), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n884), .A2(G135), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n939) );
  XNOR2_X1 U689 ( .A(n939), .B(G2096), .ZN(n615) );
  INV_X1 U690 ( .A(G2100), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U692 ( .A1(G93), .A2(n648), .ZN(n617) );
  NAND2_X1 U693 ( .A1(G80), .A2(n652), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G67), .A2(n656), .ZN(n619) );
  NAND2_X1 U696 ( .A1(G55), .A2(n649), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n670) );
  NAND2_X1 U699 ( .A1(G559), .A2(n899), .ZN(n622) );
  XOR2_X1 U700 ( .A(n978), .B(n622), .Z(n666) );
  NAND2_X1 U701 ( .A1(n623), .A2(n666), .ZN(n624) );
  XNOR2_X1 U702 ( .A(n624), .B(KEYINPUT83), .ZN(n625) );
  XOR2_X1 U703 ( .A(n670), .B(n625), .Z(G145) );
  NAND2_X1 U704 ( .A1(n652), .A2(G72), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n648), .A2(G85), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G60), .A2(n656), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G47), .A2(n649), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U711 ( .A(KEYINPUT70), .B(n632), .Z(G290) );
  NAND2_X1 U712 ( .A1(G62), .A2(n656), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G50), .A2(n649), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U715 ( .A(KEYINPUT85), .B(n635), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G88), .A2(n648), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G75), .A2(n652), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U719 ( .A(KEYINPUT86), .B(n638), .Z(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(G303) );
  INV_X1 U721 ( .A(G303), .ZN(G166) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n641) );
  XNOR2_X1 U723 ( .A(n641), .B(KEYINPUT84), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G49), .A2(n649), .ZN(n644) );
  NAND2_X1 U725 ( .A1(G87), .A2(n642), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U727 ( .A1(n656), .A2(n645), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G86), .A2(n648), .ZN(n651) );
  NAND2_X1 U730 ( .A1(G48), .A2(n649), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n652), .A2(G73), .ZN(n653) );
  XOR2_X1 U733 ( .A(KEYINPUT2), .B(n653), .Z(n654) );
  NOR2_X1 U734 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U735 ( .A1(n656), .A2(G61), .ZN(n657) );
  NAND2_X1 U736 ( .A1(n658), .A2(n657), .ZN(G305) );
  XNOR2_X1 U737 ( .A(G290), .B(G166), .ZN(n665) );
  XNOR2_X1 U738 ( .A(KEYINPUT87), .B(KEYINPUT19), .ZN(n660) );
  XNOR2_X1 U739 ( .A(G288), .B(KEYINPUT88), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U741 ( .A(n661), .B(G305), .ZN(n663) );
  XNOR2_X1 U742 ( .A(n670), .B(G299), .ZN(n662) );
  XNOR2_X1 U743 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U744 ( .A(n665), .B(n664), .ZN(n898) );
  XNOR2_X1 U745 ( .A(n898), .B(n666), .ZN(n667) );
  NAND2_X1 U746 ( .A1(n667), .A2(G868), .ZN(n668) );
  XOR2_X1 U747 ( .A(KEYINPUT89), .B(n668), .Z(n672) );
  NAND2_X1 U748 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U749 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U756 ( .A1(G236), .A2(G238), .ZN(n678) );
  NOR2_X1 U757 ( .A1(G235), .A2(G237), .ZN(n677) );
  NAND2_X1 U758 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U759 ( .A(KEYINPUT90), .B(n679), .ZN(n835) );
  NAND2_X1 U760 ( .A1(G567), .A2(n835), .ZN(n684) );
  NOR2_X1 U761 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U763 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U764 ( .A1(G96), .A2(n682), .ZN(n834) );
  NAND2_X1 U765 ( .A1(G2106), .A2(n834), .ZN(n683) );
  NAND2_X1 U766 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U767 ( .A(KEYINPUT91), .B(n685), .ZN(G319) );
  INV_X1 U768 ( .A(G319), .ZN(n687) );
  NAND2_X1 U769 ( .A1(G661), .A2(G483), .ZN(n686) );
  NOR2_X1 U770 ( .A1(n687), .A2(n686), .ZN(n833) );
  NAND2_X1 U771 ( .A1(n833), .A2(G36), .ZN(G176) );
  XOR2_X1 U772 ( .A(KEYINPUT28), .B(KEYINPUT100), .Z(n694) );
  INV_X1 U773 ( .A(n758), .ZN(n688) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n759) );
  NAND2_X1 U775 ( .A1(n688), .A2(n759), .ZN(n689) );
  XNOR2_X1 U776 ( .A(n689), .B(KEYINPUT64), .ZN(n720) );
  INV_X1 U777 ( .A(n720), .ZN(n714) );
  NAND2_X1 U778 ( .A1(G2072), .A2(n714), .ZN(n690) );
  XOR2_X1 U779 ( .A(KEYINPUT27), .B(n690), .Z(n692) );
  INV_X1 U780 ( .A(n714), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(G1956), .ZN(n691) );
  NAND2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U783 ( .A1(n695), .A2(G299), .ZN(n693) );
  XNOR2_X1 U784 ( .A(n694), .B(n693), .ZN(n712) );
  NOR2_X1 U785 ( .A1(G299), .A2(n695), .ZN(n697) );
  XNOR2_X1 U786 ( .A(n697), .B(n696), .ZN(n710) );
  NAND2_X1 U787 ( .A1(n714), .A2(G1996), .ZN(n698) );
  XNOR2_X1 U788 ( .A(n698), .B(KEYINPUT26), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n733), .A2(G1341), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U791 ( .A1(n978), .A2(n701), .ZN(n705) );
  NAND2_X1 U792 ( .A1(G2067), .A2(n714), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n733), .A2(G1348), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n706) );
  NOR2_X1 U795 ( .A1(n975), .A2(n706), .ZN(n704) );
  NOR2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n708) );
  AND2_X1 U797 ( .A1(n975), .A2(n706), .ZN(n707) );
  NOR2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U801 ( .A(n713), .B(KEYINPUT29), .ZN(n719) );
  NOR2_X1 U802 ( .A1(G1961), .A2(n714), .ZN(n716) );
  XOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .Z(n955) );
  NOR2_X1 U804 ( .A1(n733), .A2(n955), .ZN(n715) );
  NOR2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U806 ( .A(n717), .B(KEYINPUT99), .ZN(n725) );
  NAND2_X1 U807 ( .A1(G171), .A2(n725), .ZN(n718) );
  NAND2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n731) );
  NAND2_X1 U809 ( .A1(n720), .A2(G8), .ZN(n806) );
  NOR2_X1 U810 ( .A1(G1966), .A2(n806), .ZN(n744) );
  NOR2_X1 U811 ( .A1(n733), .A2(G2084), .ZN(n741) );
  NOR2_X1 U812 ( .A1(n744), .A2(n741), .ZN(n721) );
  XNOR2_X1 U813 ( .A(KEYINPUT102), .B(n721), .ZN(n722) );
  NAND2_X1 U814 ( .A1(n722), .A2(G8), .ZN(n723) );
  XNOR2_X1 U815 ( .A(n723), .B(KEYINPUT30), .ZN(n724) );
  NOR2_X1 U816 ( .A1(G168), .A2(n724), .ZN(n727) );
  NOR2_X1 U817 ( .A1(G171), .A2(n725), .ZN(n726) );
  NOR2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U819 ( .A1(n742), .A2(G286), .ZN(n732) );
  XNOR2_X1 U820 ( .A(n732), .B(KEYINPUT104), .ZN(n738) );
  NOR2_X1 U821 ( .A1(n733), .A2(G2090), .ZN(n735) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n806), .ZN(n734) );
  NOR2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U824 ( .A1(n736), .A2(G303), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U826 ( .A1(G8), .A2(n520), .ZN(n740) );
  XNOR2_X1 U827 ( .A(n740), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U828 ( .A1(G8), .A2(n741), .ZN(n746) );
  INV_X1 U829 ( .A(n742), .ZN(n743) );
  NOR2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U831 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U832 ( .A1(n748), .A2(n747), .ZN(n804) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n754) );
  NOR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n754), .A2(n749), .ZN(n980) );
  XNOR2_X1 U836 ( .A(KEYINPUT106), .B(n980), .ZN(n751) );
  INV_X1 U837 ( .A(KEYINPUT33), .ZN(n750) );
  AND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n804), .A2(n752), .ZN(n794) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n983) );
  INV_X1 U841 ( .A(n983), .ZN(n753) );
  OR2_X1 U842 ( .A1(KEYINPUT33), .A2(n519), .ZN(n792) );
  NAND2_X1 U843 ( .A1(n754), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n755), .A2(n806), .ZN(n757) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n972) );
  INV_X1 U846 ( .A(n972), .ZN(n756) );
  NOR2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n790) );
  NOR2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n825) );
  XNOR2_X1 U849 ( .A(KEYINPUT37), .B(G2067), .ZN(n823) );
  NAND2_X1 U850 ( .A1(G104), .A2(n886), .ZN(n761) );
  NAND2_X1 U851 ( .A1(G140), .A2(n884), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U853 ( .A(KEYINPUT34), .B(n762), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n880), .A2(G116), .ZN(n763) );
  XNOR2_X1 U855 ( .A(n763), .B(KEYINPUT94), .ZN(n765) );
  NAND2_X1 U856 ( .A1(G128), .A2(n881), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U858 ( .A(KEYINPUT35), .B(n766), .Z(n767) );
  NOR2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U860 ( .A(KEYINPUT36), .B(n769), .ZN(n874) );
  NOR2_X1 U861 ( .A1(n823), .A2(n874), .ZN(n923) );
  NAND2_X1 U862 ( .A1(n825), .A2(n923), .ZN(n821) );
  NAND2_X1 U863 ( .A1(G95), .A2(n886), .ZN(n771) );
  NAND2_X1 U864 ( .A1(G131), .A2(n884), .ZN(n770) );
  NAND2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U866 ( .A(KEYINPUT96), .B(n772), .ZN(n777) );
  NAND2_X1 U867 ( .A1(G107), .A2(n880), .ZN(n774) );
  NAND2_X1 U868 ( .A1(G119), .A2(n881), .ZN(n773) );
  NAND2_X1 U869 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U870 ( .A(KEYINPUT95), .B(n775), .Z(n776) );
  NOR2_X1 U871 ( .A1(n777), .A2(n776), .ZN(n894) );
  INV_X1 U872 ( .A(G1991), .ZN(n951) );
  NOR2_X1 U873 ( .A1(n894), .A2(n951), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n884), .A2(G141), .ZN(n784) );
  NAND2_X1 U875 ( .A1(G117), .A2(n880), .ZN(n779) );
  NAND2_X1 U876 ( .A1(G129), .A2(n881), .ZN(n778) );
  NAND2_X1 U877 ( .A1(n779), .A2(n778), .ZN(n782) );
  NAND2_X1 U878 ( .A1(n886), .A2(G105), .ZN(n780) );
  XOR2_X1 U879 ( .A(KEYINPUT38), .B(n780), .Z(n781) );
  NOR2_X1 U880 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U881 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U882 ( .A(KEYINPUT97), .B(n785), .Z(n873) );
  AND2_X1 U883 ( .A1(n873), .A2(G1996), .ZN(n786) );
  NOR2_X1 U884 ( .A1(n787), .A2(n786), .ZN(n932) );
  INV_X1 U885 ( .A(n825), .ZN(n788) );
  NOR2_X1 U886 ( .A1(n932), .A2(n788), .ZN(n818) );
  INV_X1 U887 ( .A(n818), .ZN(n789) );
  AND2_X1 U888 ( .A1(n821), .A2(n789), .ZN(n805) );
  AND2_X1 U889 ( .A1(n790), .A2(n805), .ZN(n791) );
  AND2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U891 ( .A1(n794), .A2(n793), .ZN(n812) );
  NAND2_X1 U892 ( .A1(G8), .A2(G166), .ZN(n795) );
  NOR2_X1 U893 ( .A1(G2090), .A2(n795), .ZN(n796) );
  XNOR2_X1 U894 ( .A(n796), .B(KEYINPUT107), .ZN(n802) );
  NOR2_X1 U895 ( .A1(G1981), .A2(G305), .ZN(n797) );
  XOR2_X1 U896 ( .A(n797), .B(KEYINPUT24), .Z(n798) );
  NOR2_X1 U897 ( .A1(n806), .A2(n798), .ZN(n799) );
  XNOR2_X1 U898 ( .A(n799), .B(KEYINPUT98), .ZN(n800) );
  AND2_X1 U899 ( .A1(n805), .A2(n800), .ZN(n808) );
  INV_X1 U900 ( .A(n808), .ZN(n801) );
  AND2_X1 U901 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n810) );
  AND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n814) );
  XNOR2_X1 U907 ( .A(G1986), .B(G290), .ZN(n977) );
  NAND2_X1 U908 ( .A1(n977), .A2(n825), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n828) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n873), .ZN(n927) );
  AND2_X1 U911 ( .A1(n951), .A2(n894), .ZN(n940) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n815) );
  XNOR2_X1 U913 ( .A(KEYINPUT108), .B(n815), .ZN(n816) );
  NOR2_X1 U914 ( .A1(n940), .A2(n816), .ZN(n817) );
  NOR2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U916 ( .A1(n927), .A2(n819), .ZN(n820) );
  XNOR2_X1 U917 ( .A(n820), .B(KEYINPUT39), .ZN(n822) );
  NAND2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n823), .A2(n874), .ZN(n925) );
  NAND2_X1 U920 ( .A1(n824), .A2(n925), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U923 ( .A(KEYINPUT40), .B(n829), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U926 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  NOR2_X1 U931 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U933 ( .A(G1981), .B(KEYINPUT41), .ZN(n845) );
  XOR2_X1 U934 ( .A(G1956), .B(G1961), .Z(n837) );
  XNOR2_X1 U935 ( .A(G1986), .B(G1966), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U937 ( .A(G1971), .B(G1976), .Z(n839) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U940 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U941 ( .A(KEYINPUT114), .B(G2474), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(G229) );
  XOR2_X1 U944 ( .A(KEYINPUT43), .B(G2678), .Z(n847) );
  XNOR2_X1 U945 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT42), .B(G2090), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U951 ( .A(G2096), .B(G2100), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n855) );
  XOR2_X1 U953 ( .A(G2078), .B(G2084), .Z(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G227) );
  NAND2_X1 U955 ( .A1(G100), .A2(n886), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G112), .A2(n880), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n858), .B(KEYINPUT115), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G136), .A2(n884), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n863) );
  NAND2_X1 U961 ( .A1(n881), .A2(G124), .ZN(n861) );
  XOR2_X1 U962 ( .A(KEYINPUT44), .B(n861), .Z(n862) );
  NOR2_X1 U963 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U964 ( .A1(G103), .A2(n886), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G139), .A2(n884), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U967 ( .A1(G115), .A2(n880), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G127), .A2(n881), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n933) );
  XNOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n871), .B(KEYINPUT117), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n933), .B(n872), .ZN(n876) );
  XOR2_X1 U975 ( .A(n874), .B(n873), .Z(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U977 ( .A(n877), .B(G162), .Z(n879) );
  XNOR2_X1 U978 ( .A(G164), .B(n939), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n879), .B(n878), .ZN(n893) );
  NAND2_X1 U980 ( .A1(G118), .A2(n880), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G130), .A2(n881), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n891) );
  NAND2_X1 U983 ( .A1(n884), .A2(G142), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n885), .B(KEYINPUT116), .ZN(n888) );
  NAND2_X1 U985 ( .A1(G106), .A2(n886), .ZN(n887) );
  NAND2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U987 ( .A(n889), .B(KEYINPUT45), .Z(n890) );
  NOR2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U989 ( .A(n893), .B(n892), .Z(n896) );
  XOR2_X1 U990 ( .A(n894), .B(G160), .Z(n895) );
  XNOR2_X1 U991 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U992 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U993 ( .A(n898), .B(KEYINPUT118), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n978), .B(n899), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U996 ( .A(G286), .B(G171), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G37), .A2(n904), .ZN(G397) );
  XOR2_X1 U999 ( .A(G2438), .B(G2435), .Z(n906) );
  XNOR2_X1 U1000 ( .A(KEYINPUT110), .B(G2454), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1002 ( .A(n907), .B(G2430), .Z(n909) );
  XNOR2_X1 U1003 ( .A(G1341), .B(G1348), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n913) );
  XOR2_X1 U1005 ( .A(G2427), .B(KEYINPUT111), .Z(n911) );
  XNOR2_X1 U1006 ( .A(G2443), .B(G2446), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1008 ( .A(n913), .B(n912), .Z(n915) );
  XNOR2_X1 U1009 ( .A(KEYINPUT109), .B(G2451), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n916) );
  NAND2_X1 U1011 ( .A1(n916), .A2(G14), .ZN(n922) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n922), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(n922), .ZN(G401) );
  INV_X1 U1020 ( .A(n923), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n945) );
  XOR2_X1 U1022 ( .A(G160), .B(G2084), .Z(n930) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(KEYINPUT51), .B(n928), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n938) );
  XOR2_X1 U1028 ( .A(G2072), .B(n933), .Z(n935) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n936), .Z(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n943) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1034 ( .A(KEYINPUT119), .B(n941), .Z(n942) );
  NAND2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1037 ( .A(KEYINPUT52), .B(n946), .Z(n947) );
  NOR2_X1 U1038 ( .A1(KEYINPUT55), .A2(n947), .ZN(n948) );
  XOR2_X1 U1039 ( .A(KEYINPUT120), .B(n948), .Z(n949) );
  NAND2_X1 U1040 ( .A1(G29), .A2(n949), .ZN(n1027) );
  XNOR2_X1 U1041 ( .A(G2084), .B(G34), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(n950), .B(KEYINPUT54), .ZN(n967) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n964) );
  XNOR2_X1 U1044 ( .A(G25), .B(n951), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n952), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1046 ( .A(G1996), .B(G32), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G27), .B(n955), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(KEYINPUT53), .B(n962), .ZN(n963) );
  NOR2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(n965), .B(KEYINPUT121), .ZN(n966) );
  NOR2_X1 U1057 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1058 ( .A(KEYINPUT55), .B(n968), .Z(n969) );
  NOR2_X1 U1059 ( .A1(G29), .A2(n969), .ZN(n970) );
  XOR2_X1 U1060 ( .A(KEYINPUT122), .B(n970), .Z(n971) );
  NAND2_X1 U1061 ( .A1(G11), .A2(n971), .ZN(n1025) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT56), .ZN(n996) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G168), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(KEYINPUT57), .B(n974), .ZN(n994) );
  XNOR2_X1 U1066 ( .A(G1348), .B(n975), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n991) );
  XOR2_X1 U1068 ( .A(G1341), .B(n978), .Z(n979) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n989) );
  XNOR2_X1 U1070 ( .A(G171), .B(G1961), .ZN(n987) );
  XOR2_X1 U1071 ( .A(G1956), .B(KEYINPUT123), .Z(n981) );
  XNOR2_X1 U1072 ( .A(G299), .B(n981), .ZN(n985) );
  NAND2_X1 U1073 ( .A1(G1971), .A2(G303), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1079 ( .A(KEYINPUT124), .B(n992), .Z(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1081 ( .A1(n996), .A2(n995), .ZN(n1023) );
  INV_X1 U1082 ( .A(G16), .ZN(n1021) );
  XNOR2_X1 U1083 ( .A(KEYINPUT127), .B(G1966), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(n997), .B(G21), .ZN(n1011) );
  XNOR2_X1 U1085 ( .A(KEYINPUT125), .B(G1956), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(n998), .B(G20), .ZN(n1003) );
  XOR2_X1 U1087 ( .A(G1348), .B(KEYINPUT59), .Z(n999) );
  XNOR2_X1 U1088 ( .A(G4), .B(n999), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G6), .B(G1981), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G19), .B(G1341), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(KEYINPUT126), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(KEYINPUT60), .B(n1007), .Z(n1009) );
  XNOR2_X1 U1096 ( .A(G1961), .B(G5), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1018) );
  XNOR2_X1 U1099 ( .A(G1976), .B(G23), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(G1986), .B(G24), .Z(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(KEYINPUT58), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

