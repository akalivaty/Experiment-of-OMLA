//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1383,
    new_n1384;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n204), .A2(new_n205), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT65), .B(G238), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n219), .A2(G68), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G58), .A2(G232), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n211), .B(new_n218), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND2_X1  g0044(.A1(new_n203), .A2(G20), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n216), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n216), .A2(new_n248), .ZN(new_n249));
  OAI221_X1 g0049(.A(new_n245), .B1(new_n246), .B2(new_n247), .C1(new_n213), .C2(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n215), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT11), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n253), .A2(new_n254), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n251), .A2(new_n215), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G1), .B2(new_n216), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT12), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n260), .B1(new_n263), .B2(new_n203), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n262), .A2(KEYINPUT12), .A3(G68), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n259), .A2(new_n203), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n256), .A2(new_n257), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  OAI211_X1 g0071(.A(G1), .B(G13), .C1(new_n248), .C2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n272), .A2(new_n268), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n270), .B1(new_n273), .B2(G238), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n272), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G33), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n277), .A2(new_n279), .A3(G232), .A4(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT71), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n283), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G97), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT66), .B(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G226), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n276), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n275), .B1(new_n291), .B2(KEYINPUT72), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT13), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT66), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT66), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G1698), .ZN(new_n297));
  AND4_X1   g0097(.A1(new_n277), .A2(new_n279), .A3(new_n295), .A4(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n298), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n282), .A2(new_n284), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n272), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT72), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n292), .A2(new_n293), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n274), .B1(new_n301), .B2(new_n302), .ZN(new_n305));
  AOI211_X1 g0105(.A(KEYINPUT72), .B(new_n272), .C1(new_n299), .C2(new_n300), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT13), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n267), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n304), .B2(new_n307), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n293), .B1(new_n292), .B2(new_n303), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n305), .A2(KEYINPUT13), .A3(new_n306), .ZN(new_n315));
  OAI21_X1  g0115(.A(G169), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT14), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n308), .A2(new_n318), .A3(G169), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n304), .A2(new_n307), .A3(G179), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n267), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n313), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n283), .A2(G223), .A3(G1698), .ZN(new_n324));
  INV_X1    g0124(.A(G222), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n324), .B1(new_n247), .B2(new_n283), .C1(new_n288), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n276), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n270), .B1(new_n273), .B2(G226), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G169), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT8), .B(G58), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT67), .ZN(new_n333));
  INV_X1    g0133(.A(G150), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n333), .A2(new_n246), .B1(new_n334), .B2(new_n249), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n216), .B1(new_n212), .B2(new_n213), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n252), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n262), .A2(G50), .ZN(new_n338));
  INV_X1    g0138(.A(new_n259), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(G50), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  OR3_X1    g0141(.A1(new_n331), .A2(new_n341), .A3(KEYINPUT68), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT68), .B1(new_n331), .B2(new_n341), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n330), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n329), .A2(G200), .ZN(new_n348));
  XOR2_X1   g0148(.A(new_n348), .B(KEYINPUT70), .Z(new_n349));
  OR2_X1    g0149(.A1(new_n341), .A2(KEYINPUT9), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n341), .A2(KEYINPUT9), .B1(G190), .B2(new_n330), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT10), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT10), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n349), .A2(new_n350), .A3(new_n354), .A4(new_n351), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n347), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n270), .B1(new_n273), .B2(G232), .ZN(new_n357));
  INV_X1    g0157(.A(G87), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n248), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n295), .A2(new_n297), .A3(G223), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G226), .A2(G1698), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT73), .B1(new_n248), .B2(KEYINPUT3), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT73), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(new_n278), .A3(G33), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n363), .A2(new_n365), .A3(new_n277), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n359), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n357), .B(G179), .C1(new_n367), .C2(new_n272), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT75), .ZN(new_n369));
  INV_X1    g0169(.A(new_n270), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n272), .A2(new_n268), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n230), .ZN(new_n372));
  INV_X1    g0172(.A(new_n359), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n287), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n363), .A2(new_n365), .A3(new_n277), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n372), .B1(new_n376), .B2(new_n276), .ZN(new_n377));
  INV_X1    g0177(.A(G169), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n368), .B(new_n369), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n357), .B1(new_n367), .B2(new_n272), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G169), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n369), .B1(new_n382), .B2(new_n368), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n333), .A2(new_n259), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n263), .B2(new_n333), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n375), .A2(new_n216), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT7), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n375), .A2(new_n389), .A3(new_n216), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(G68), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n204), .A2(new_n205), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G20), .ZN(new_n394));
  INV_X1    g0194(.A(G159), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n249), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT74), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n396), .B1(new_n393), .B2(G20), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT74), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n391), .A2(KEYINPUT16), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n252), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n400), .B(KEYINPUT74), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT7), .B1(new_n283), .B2(G20), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n277), .A2(new_n279), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n389), .A3(new_n216), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n408), .A3(G68), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT16), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n386), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n384), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT18), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n384), .A2(new_n414), .A3(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n357), .B(new_n309), .C1(new_n367), .C2(new_n272), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n377), .B2(G200), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(new_n386), .C1(new_n404), .C2(new_n410), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n262), .A2(G77), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n259), .B2(new_n247), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G20), .A2(G77), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT15), .B(G87), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n427), .B1(new_n332), .B2(new_n249), .C1(new_n246), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n252), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n219), .A2(new_n283), .A3(G1698), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n407), .A2(G107), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(new_n288), .C2(new_n230), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n276), .ZN(new_n435));
  INV_X1    g0235(.A(G244), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n370), .B1(new_n371), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n431), .B1(new_n439), .B2(G200), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n309), .B2(new_n439), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n425), .B1(new_n252), .B2(new_n429), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n439), .B2(new_n378), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n437), .B1(new_n434), .B2(new_n276), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n444), .A2(KEYINPUT69), .A3(new_n344), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT69), .B1(new_n444), .B2(new_n344), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AND4_X1   g0249(.A1(new_n323), .A2(new_n356), .A3(new_n422), .A4(new_n449), .ZN(new_n450));
  AND2_X1   g0250(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n451));
  NOR2_X1   g0251(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n271), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT77), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(KEYINPUT77), .B(new_n271), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n261), .A2(G45), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n458), .B2(G41), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(G257), .A3(new_n272), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n455), .A2(new_n456), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT78), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n455), .A2(KEYINPUT78), .A3(new_n456), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(G274), .A3(new_n272), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT4), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n295), .A2(new_n297), .A3(G244), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n375), .B2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n277), .A2(new_n279), .A3(G250), .A4(G1698), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n283), .A2(new_n287), .A3(KEYINPUT4), .A4(G244), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n276), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n460), .A2(KEYINPUT79), .A3(G257), .A4(new_n272), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n463), .A2(new_n470), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT80), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n468), .B1(new_n464), .B2(new_n465), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(new_n467), .B1(new_n478), .B2(new_n276), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n485), .A2(KEYINPUT80), .A3(new_n480), .A4(new_n463), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n486), .A3(G190), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT6), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n488), .A2(new_n489), .A3(G107), .ZN(new_n490));
  XNOR2_X1  g0290(.A(G97), .B(G107), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n492), .A2(new_n216), .B1(new_n247), .B2(new_n249), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n406), .A2(new_n408), .A3(G107), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n252), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n263), .A2(new_n489), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n258), .B(new_n262), .C1(G1), .C2(new_n248), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G97), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n481), .B2(G200), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n487), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n363), .A2(new_n365), .A3(new_n216), .A4(new_n277), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT19), .ZN(new_n504));
  INV_X1    g0304(.A(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n358), .A2(new_n489), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n286), .A2(new_n216), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n246), .A2(KEYINPUT19), .A3(new_n489), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n203), .A2(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(new_n252), .B1(new_n263), .B2(new_n428), .ZN(new_n511));
  INV_X1    g0311(.A(new_n428), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n498), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n511), .A2(new_n516), .A3(new_n513), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n287), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n519));
  INV_X1    g0319(.A(G116), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT81), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT81), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G116), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n519), .A2(new_n375), .B1(new_n248), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n276), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n457), .A2(G250), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n276), .A2(new_n527), .B1(new_n269), .B2(new_n457), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(G169), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n525), .B2(new_n276), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n344), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n498), .A2(G87), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n511), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n311), .B1(new_n526), .B2(new_n529), .ZN(new_n535));
  AOI211_X1 g0335(.A(new_n309), .B(new_n528), .C1(new_n525), .C2(new_n276), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n518), .A2(new_n532), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(G169), .B1(new_n483), .B2(new_n486), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n500), .B1(new_n481), .B2(G179), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n502), .B(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n460), .A2(G270), .A3(new_n272), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n287), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n544));
  INV_X1    g0344(.A(G303), .ZN(new_n545));
  OAI22_X1  g0345(.A1(new_n544), .A2(new_n375), .B1(new_n545), .B2(new_n283), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n276), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n470), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n521), .A2(new_n523), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n497), .A2(new_n520), .B1(new_n262), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n524), .A2(G20), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n475), .B(new_n216), .C1(G33), .C2(new_n489), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n552), .A2(KEYINPUT20), .A3(new_n252), .A4(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n252), .B(new_n553), .C1(new_n549), .C2(new_n216), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT20), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n378), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n548), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n470), .A2(new_n547), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n551), .A2(new_n558), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n563), .A2(G179), .A3(new_n543), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n548), .A2(new_n559), .A3(KEYINPUT21), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n564), .B1(new_n548), .B2(G200), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n309), .B2(new_n548), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n505), .A2(G20), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT23), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n549), .A2(new_n216), .A3(G33), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n366), .A2(KEYINPUT22), .A3(new_n216), .A4(G87), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT22), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n216), .A2(G87), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n579), .B1(new_n407), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n574), .A3(new_n575), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n503), .A2(new_n579), .A3(new_n358), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT24), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n258), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT25), .B1(new_n263), .B2(new_n505), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n505), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n498), .A2(G107), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT83), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT83), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n582), .A2(new_n585), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n593), .B(new_n590), .C1(new_n594), .C2(new_n258), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n287), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n596));
  INV_X1    g0396(.A(G294), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n596), .A2(new_n375), .B1(new_n248), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n276), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n460), .A2(G264), .A3(new_n272), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n470), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(KEYINPUT84), .A3(G169), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n470), .A2(G179), .A3(new_n599), .A4(new_n600), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT84), .B1(new_n601), .B2(G169), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n592), .B(new_n595), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n470), .A2(new_n599), .A3(new_n600), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G190), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n586), .A2(new_n591), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n601), .A2(G200), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n571), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n450), .A2(new_n542), .A3(new_n613), .ZN(G372));
  NAND2_X1  g0414(.A1(new_n353), .A2(new_n355), .ZN(new_n615));
  INV_X1    g0415(.A(new_n312), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n616), .B(new_n267), .C1(new_n309), .C2(new_n308), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n431), .B1(new_n444), .B2(G169), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT69), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n439), .B2(G179), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n444), .A2(KEYINPUT69), .A3(new_n344), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n319), .A2(new_n320), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n378), .B1(new_n304), .B2(new_n307), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(new_n318), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n322), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n421), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n368), .B1(new_n377), .B2(new_n378), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n411), .A2(new_n414), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n414), .B1(new_n411), .B2(new_n629), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n615), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n346), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n518), .A2(new_n532), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n483), .A2(new_n486), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n378), .ZN(new_n639));
  INV_X1    g0439(.A(new_n540), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n538), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n540), .B1(new_n638), .B2(new_n378), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(KEYINPUT26), .A3(new_n538), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n637), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT84), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n607), .B2(new_n378), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n602), .A3(new_n603), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n568), .B1(new_n650), .B2(new_n609), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n639), .A2(new_n640), .B1(new_n487), .B2(new_n501), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(new_n538), .A4(new_n611), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n450), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n635), .A2(new_n655), .ZN(G369));
  AND2_X1   g0456(.A1(new_n595), .A2(new_n592), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n261), .A2(new_n216), .A3(G13), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(KEYINPUT85), .B(G343), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g0464(.A(new_n664), .B(KEYINPUT86), .Z(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n657), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n606), .A3(new_n611), .ZN(new_n668));
  INV_X1    g0468(.A(new_n606), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n666), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n665), .B1(new_n558), .B2(new_n551), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n567), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n571), .B2(new_n672), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n674), .A2(KEYINPUT87), .A3(G330), .ZN(new_n675));
  AOI21_X1  g0475(.A(KEYINPUT87), .B1(new_n674), .B2(G330), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n567), .A2(new_n665), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n612), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n609), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n649), .A2(new_n680), .A3(new_n665), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n677), .A2(new_n683), .ZN(G399));
  NOR2_X1   g0484(.A1(new_n506), .A2(G116), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n209), .A2(new_n271), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(G1), .ZN(new_n687));
  INV_X1    g0487(.A(new_n214), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n654), .A2(new_n665), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT29), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n644), .A2(KEYINPUT26), .A3(new_n538), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT26), .B1(new_n644), .B2(new_n538), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n636), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n567), .B1(new_n657), .B2(new_n649), .ZN(new_n697));
  INV_X1    g0497(.A(new_n611), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n541), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI211_X1 g0499(.A(KEYINPUT29), .B(new_n665), .C1(new_n696), .C2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n548), .A2(new_n344), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n531), .A2(new_n599), .A3(new_n600), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n483), .A2(new_n486), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n531), .A2(G179), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n707), .A2(new_n548), .A3(new_n601), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n705), .A2(new_n706), .B1(new_n708), .B2(new_n481), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n703), .A2(new_n548), .A3(new_n344), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(KEYINPUT30), .A3(new_n483), .A4(new_n486), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n665), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT31), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT88), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n613), .A2(new_n542), .A3(new_n665), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT88), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n712), .A2(new_n716), .A3(KEYINPUT31), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n705), .A2(new_n706), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n708), .A2(new_n481), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(new_n711), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n666), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n714), .A2(new_n715), .A3(new_n717), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n701), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n690), .B1(new_n727), .B2(G1), .ZN(G364));
  NOR2_X1   g0528(.A1(new_n675), .A2(new_n676), .ZN(new_n729));
  INV_X1    g0529(.A(new_n686), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n216), .A2(G13), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT89), .Z(new_n732));
  AOI21_X1  g0532(.A(new_n261), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n729), .B1(G330), .B2(new_n674), .C1(new_n730), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n730), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n283), .A2(new_n209), .ZN(new_n737));
  INV_X1    g0537(.A(G355), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n737), .A2(new_n738), .B1(G116), .B2(new_n209), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n375), .A2(new_n209), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n243), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(G45), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n214), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n739), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(G1), .B(G13), .C1(new_n216), .C2(G169), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n745), .A2(KEYINPUT90), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(KEYINPUT90), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n736), .B1(new_n744), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n216), .A2(G190), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT92), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT92), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n395), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT32), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n216), .B1(new_n756), .B2(G190), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT93), .Z(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G97), .ZN(new_n765));
  INV_X1    g0565(.A(new_n755), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n766), .A2(new_n344), .A3(G200), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n767), .A2(KEYINPUT91), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(KEYINPUT91), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G77), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n216), .A2(new_n309), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G179), .A3(new_n311), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n344), .A2(new_n311), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n774), .A2(new_n202), .B1(new_n776), .B2(new_n213), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n755), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n311), .A2(G179), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n755), .A2(new_n779), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n778), .A2(new_n203), .B1(new_n780), .B2(new_n505), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n773), .A2(new_n779), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n283), .B1(new_n782), .B2(new_n358), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n777), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n762), .A2(new_n765), .A3(new_n772), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT94), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  INV_X1    g0588(.A(G322), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n407), .B1(new_n774), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n778), .ZN(new_n791));
  INV_X1    g0591(.A(G317), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n791), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  INV_X1    g0596(.A(new_n767), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n795), .B1(new_n796), .B2(new_n780), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n763), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n790), .B(new_n799), .C1(G294), .C2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n776), .B(KEYINPUT95), .Z(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT96), .B(G326), .Z(new_n804));
  INV_X1    g0604(.A(new_n760), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(G329), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n782), .A2(KEYINPUT97), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n782), .A2(KEYINPUT97), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n801), .B(new_n806), .C1(new_n545), .C2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n787), .A2(new_n788), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n754), .B1(new_n811), .B2(new_n748), .ZN(new_n812));
  INV_X1    g0612(.A(new_n751), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n674), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n735), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  INV_X1    g0616(.A(KEYINPUT99), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n447), .B2(new_n665), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n622), .A2(KEYINPUT99), .A3(new_n666), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT100), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n441), .B(new_n447), .C1(new_n442), .C2(new_n665), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n821), .B1(new_n820), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n691), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n447), .A2(new_n817), .A3(new_n665), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT99), .B1(new_n622), .B2(new_n666), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(KEYINPUT100), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n567), .B1(new_n649), .B2(new_n680), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n541), .A2(new_n833), .A3(new_n698), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n832), .B(new_n665), .C1(new_n696), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n826), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n736), .B1(new_n836), .B2(new_n725), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n725), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n748), .A2(new_n749), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n736), .B1(new_n840), .B2(G77), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n780), .A2(new_n203), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n375), .B(new_n842), .C1(G58), .C2(new_n800), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n213), .B2(new_n809), .C1(new_n844), .C2(new_n760), .ZN(new_n845));
  INV_X1    g0645(.A(new_n774), .ZN(new_n846));
  INV_X1    g0646(.A(new_n776), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n846), .A2(G143), .B1(new_n847), .B2(G137), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n334), .B2(new_n778), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n771), .B2(G159), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n845), .B1(KEYINPUT34), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(KEYINPUT34), .B2(new_n850), .ZN(new_n852));
  XNOR2_X1  g0652(.A(KEYINPUT98), .B(G283), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n774), .A2(new_n597), .B1(new_n778), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n780), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(G87), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n407), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n854), .B(new_n857), .C1(G303), .C2(new_n847), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n809), .A2(new_n505), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n771), .B2(new_n549), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n805), .A2(G311), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n858), .A2(new_n860), .A3(new_n765), .A4(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n841), .B1(new_n864), .B2(new_n748), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n832), .B2(new_n750), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n838), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(G384));
  INV_X1    g0668(.A(new_n492), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n869), .A2(KEYINPUT35), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(KEYINPUT35), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(G116), .A3(new_n217), .A4(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(KEYINPUT101), .B(KEYINPUT36), .Z(new_n873));
  XNOR2_X1  g0673(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n214), .A2(G77), .A3(new_n392), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n213), .A2(G68), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n261), .B(G13), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT16), .B1(new_n405), .B2(new_n391), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n386), .B1(new_n404), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n661), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n384), .A2(new_n414), .A3(new_n411), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n414), .B1(new_n384), .B2(new_n411), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n419), .B(KEYINPUT17), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n881), .A2(new_n629), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n882), .A2(new_n888), .A3(new_n419), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n419), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n411), .B1(new_n384), .B2(new_n661), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n889), .A2(KEYINPUT37), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n879), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT102), .ZN(new_n896));
  INV_X1    g0696(.A(new_n882), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n416), .B2(new_n421), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n892), .A2(new_n893), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n895), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(KEYINPUT102), .B(new_n879), .C1(new_n887), .C2(new_n894), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT106), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n712), .B2(KEYINPUT31), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n721), .A2(KEYINPUT106), .A3(new_n722), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n715), .A2(new_n906), .A3(new_n907), .A4(new_n713), .ZN(new_n908));
  INV_X1    g0708(.A(new_n308), .ZN(new_n909));
  AOI22_X1  g0709(.A1(G179), .A2(new_n909), .B1(new_n625), .B2(new_n318), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n267), .B1(new_n910), .B2(new_n317), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n666), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n666), .A2(new_n322), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n627), .A2(new_n617), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n825), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n903), .A2(new_n904), .A3(new_n908), .A4(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n411), .A2(new_n629), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n411), .A2(new_n661), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(new_n921), .A3(new_n419), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n922), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT103), .B1(new_n922), .B2(KEYINPUT37), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n629), .A2(KEYINPUT75), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n379), .ZN(new_n926));
  INV_X1    g0726(.A(new_n661), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n399), .A2(new_n402), .A3(new_n409), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n252), .B(new_n403), .C1(new_n928), .C2(KEYINPUT16), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n926), .A2(new_n927), .B1(new_n929), .B2(new_n386), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(new_n891), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n923), .A2(new_n924), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n921), .B1(new_n632), .B2(new_n886), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n879), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n919), .B1(new_n934), .B2(new_n902), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n915), .A2(new_n908), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n918), .A2(new_n937), .A3(G330), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n450), .A2(new_n908), .A3(G330), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT107), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(KEYINPUT107), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n916), .A2(new_n917), .B1(new_n935), .B2(new_n936), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n450), .A3(new_n908), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n622), .A2(new_n665), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n835), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n912), .A2(new_n914), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n948), .A2(new_n904), .A3(new_n903), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n633), .A2(new_n927), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n911), .A2(new_n665), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT39), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT103), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n931), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n922), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n933), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n955), .B(new_n902), .C1(new_n960), .C2(KEYINPUT38), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(KEYINPUT104), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT104), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n934), .A2(new_n963), .A3(new_n955), .A4(new_n902), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n904), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n952), .B1(new_n954), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n693), .A2(new_n450), .A3(new_n700), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n968), .A2(new_n635), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n946), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n261), .B2(new_n732), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n946), .A2(new_n970), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n878), .B1(new_n972), .B2(new_n973), .ZN(G367));
  OAI21_X1  g0774(.A(new_n752), .B1(new_n209), .B2(new_n428), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n236), .A2(new_n740), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n736), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n807), .A2(KEYINPUT46), .A3(G116), .A4(new_n808), .ZN(new_n978));
  XOR2_X1   g0778(.A(KEYINPUT114), .B(G317), .Z(new_n979));
  OAI221_X1 g0779(.A(new_n978), .B1(new_n760), .B2(new_n979), .C1(new_n770), .C2(new_n853), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G294), .A2(new_n791), .B1(new_n855), .B2(G97), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n545), .B2(new_n774), .C1(new_n802), .C2(new_n798), .ZN(new_n982));
  INV_X1    g0782(.A(new_n782), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT46), .B1(new_n983), .B2(new_n549), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n375), .B1(new_n505), .B2(new_n763), .ZN(new_n985));
  NOR4_X1   g0785(.A1(new_n980), .A2(new_n982), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n855), .A2(G77), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n283), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT116), .Z(new_n989));
  OAI22_X1  g0789(.A1(new_n202), .A2(new_n782), .B1(new_n778), .B2(new_n395), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n803), .B2(G143), .ZN(new_n991));
  INV_X1    g0791(.A(G137), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n991), .B1(new_n213), .B2(new_n770), .C1(new_n992), .C2(new_n760), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT115), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n764), .A2(G68), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n334), .B2(new_n774), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n989), .B(new_n993), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n994), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n986), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT47), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n999), .A2(KEYINPUT47), .B1(new_n746), .B2(new_n747), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n977), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n665), .A2(new_n534), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n538), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT108), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(KEYINPUT108), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1003), .A2(new_n636), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(new_n813), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT113), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1008), .B(KEYINPUT43), .Z(new_n1012));
  INV_X1    g0812(.A(KEYINPUT42), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n666), .A2(new_n500), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n502), .B(new_n1014), .C1(new_n539), .C2(new_n540), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n644), .A2(new_n666), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT110), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1017), .A2(new_n679), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1018), .B1(new_n1017), .B2(new_n679), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1013), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1017), .A2(new_n679), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(KEYINPUT110), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1024), .A2(KEYINPUT42), .A3(new_n1019), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1015), .A2(KEYINPUT109), .A3(new_n1016), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(KEYINPUT109), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n669), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n644), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n666), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(KEYINPUT111), .B(new_n1012), .C1(new_n1026), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1029), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n606), .B1(new_n1034), .B2(new_n1027), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n665), .B1(new_n1035), .B2(new_n644), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1008), .A2(KEYINPUT43), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1036), .A2(new_n1025), .A3(new_n1022), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n1025), .A3(new_n1022), .ZN(new_n1040));
  AOI21_X1  g0840(.A(KEYINPUT111), .B1(new_n1040), .B2(new_n1012), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT112), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1012), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT111), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT112), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1045), .A2(new_n1046), .A3(new_n1033), .A4(new_n1038), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1034), .A2(new_n1027), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n677), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1051), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1042), .A2(new_n1053), .A3(new_n1047), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT44), .ZN(new_n1056));
  OR3_X1    g0856(.A1(new_n683), .A2(new_n1056), .A3(new_n1017), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1056), .B1(new_n683), .B2(new_n1017), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n683), .A2(new_n1017), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT45), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n683), .A2(KEYINPUT45), .A3(new_n1017), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n1059), .A2(new_n677), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n677), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n671), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n679), .B1(new_n1068), .B2(new_n678), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n729), .B(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n726), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n686), .B(KEYINPUT41), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n733), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1011), .B1(new_n1055), .B2(new_n1073), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n1042), .A2(new_n1053), .A3(new_n1047), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1053), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1073), .B(new_n1011), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1010), .B1(new_n1074), .B2(new_n1078), .ZN(G387));
  OAI22_X1  g0879(.A1(new_n737), .A2(new_n685), .B1(G107), .B2(new_n209), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n233), .A2(new_n742), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n685), .ZN(new_n1082));
  AOI211_X1 g0882(.A(G45), .B(new_n1082), .C1(G68), .C2(G77), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n332), .A2(G50), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT50), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n740), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1080), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n736), .B1(new_n1087), .B2(new_n753), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n797), .A2(new_n203), .B1(new_n780), .B2(new_n489), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n774), .A2(new_n213), .B1(new_n782), .B2(new_n247), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n1089), .A2(new_n375), .A3(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n776), .A2(new_n395), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT117), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n333), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n805), .A2(G150), .B1(new_n1094), .B2(new_n791), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n764), .A2(new_n512), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1091), .A2(new_n1093), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n803), .A2(G322), .B1(G311), .B2(new_n791), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT118), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n545), .B2(new_n770), .C1(new_n774), .C2(new_n979), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1101), .A2(KEYINPUT48), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n782), .A2(new_n597), .B1(new_n763), .B2(new_n853), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1101), .B2(KEYINPUT48), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(KEYINPUT49), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n375), .B1(new_n524), .B2(new_n780), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n805), .B2(new_n804), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT49), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1097), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1088), .B1(new_n1110), .B2(new_n748), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1068), .A2(new_n751), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1111), .A2(new_n1112), .B1(new_n1070), .B2(new_n734), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n727), .A2(new_n1070), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n730), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n727), .A2(new_n1070), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(G393));
  AND2_X1   g0917(.A1(new_n727), .A2(new_n1070), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n686), .B1(new_n1118), .B2(new_n1067), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1114), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1067), .A2(new_n734), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n752), .B1(new_n489), .B2(new_n209), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n240), .A2(new_n209), .A3(new_n375), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n736), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n797), .A2(new_n597), .B1(new_n782), .B2(new_n853), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(G303), .B2(new_n791), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n774), .A2(new_n798), .B1(new_n776), .B2(new_n792), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT52), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n805), .A2(G322), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n407), .B1(new_n780), .B2(new_n505), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n549), .B2(new_n800), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1127), .A2(new_n1129), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n774), .A2(new_n395), .B1(new_n776), .B2(new_n334), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT51), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n805), .A2(G143), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(new_n332), .C2(new_n770), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n856), .B1(new_n203), .B2(new_n782), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G50), .B2(new_n791), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n764), .A2(G77), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n366), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1133), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1125), .B1(new_n1142), .B2(new_n748), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n1049), .B2(new_n813), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1121), .A2(new_n1122), .A3(new_n1144), .ZN(G390));
  OAI211_X1 g0945(.A(new_n665), .B(new_n832), .C1(new_n696), .C2(new_n699), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n947), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n949), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n954), .B1(new_n934), .B2(new_n902), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n1149), .A3(KEYINPUT119), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT119), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n956), .A2(new_n957), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(new_n900), .A3(new_n959), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n933), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT38), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n902), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n953), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n323), .A2(new_n913), .B1(new_n911), .B2(new_n666), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n1146), .B2(new_n947), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1151), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1150), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n947), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n666), .B1(new_n646), .B2(new_n653), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n832), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n953), .B1(new_n1164), .B2(new_n1158), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1165), .A2(new_n962), .A3(new_n964), .A4(new_n965), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n832), .A2(G330), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n908), .A2(new_n949), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n724), .A2(new_n949), .A3(new_n1168), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1161), .A2(new_n1166), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n734), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT120), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT120), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1170), .A2(new_n1175), .A3(new_n734), .A4(new_n1172), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n968), .A2(new_n635), .A3(new_n939), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n949), .B1(new_n724), .B2(new_n1168), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n948), .B1(new_n1169), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1147), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n908), .A2(new_n1168), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1182), .B(new_n1171), .C1(new_n1183), .C2(new_n949), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1179), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1178), .A2(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1188), .A2(new_n1165), .B1(new_n1160), .B2(new_n1150), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1169), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1172), .B(new_n1185), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1187), .A2(new_n730), .A3(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n736), .B1(new_n840), .B2(new_n1094), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n771), .A2(G97), .B1(G294), .B2(new_n805), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n358), .B2(new_n809), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n842), .A2(new_n283), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n776), .A2(new_n796), .B1(new_n778), .B2(new_n505), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G116), .B2(new_n846), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1140), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n805), .A2(G125), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n774), .A2(new_n844), .B1(new_n780), .B2(new_n213), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G128), .B2(new_n847), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT54), .B(G143), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1200), .B(new_n1202), .C1(new_n770), .C2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n764), .A2(G159), .ZN(new_n1205));
  OR3_X1    g1005(.A1(new_n782), .A2(KEYINPUT53), .A3(new_n334), .ZN(new_n1206));
  OAI21_X1  g1006(.A(KEYINPUT53), .B1(new_n782), .B2(new_n334), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n407), .B1(new_n791), .B2(G137), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n1195), .A2(new_n1199), .B1(new_n1204), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1193), .B1(new_n1210), .B2(new_n748), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n966), .B2(new_n750), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1177), .A2(new_n1192), .A3(new_n1212), .ZN(G378));
  INV_X1    g1013(.A(new_n1179), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1191), .A2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n950), .B(new_n951), .C1(new_n1188), .C2(new_n953), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n615), .A2(new_n346), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n341), .A2(new_n927), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n615), .B(new_n346), .C1(new_n341), .C2(new_n927), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1219), .A2(new_n1220), .A3(new_n1222), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n944), .B2(G330), .ZN(new_n1227));
  AND4_X1   g1027(.A1(G330), .A2(new_n918), .A3(new_n937), .A4(new_n1226), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1216), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1226), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n938), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n944), .A2(G330), .A3(new_n1226), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n967), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1229), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1215), .A2(KEYINPUT57), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT122), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1215), .A2(new_n1234), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT57), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT122), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1215), .A2(new_n1234), .A3(new_n1240), .A4(KEYINPUT57), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1236), .A2(new_n1239), .A3(new_n730), .A4(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1234), .A2(new_n734), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n736), .B1(new_n840), .B2(G50), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n366), .A2(G41), .ZN(new_n1245));
  AOI211_X1 g1045(.A(G50), .B(new_n1245), .C1(new_n248), .C2(new_n271), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n797), .A2(new_n428), .B1(new_n520), .B2(new_n776), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n247), .A2(new_n782), .B1(new_n778), .B2(new_n489), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n774), .A2(new_n505), .B1(new_n780), .B2(new_n202), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n805), .A2(G283), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(new_n995), .A3(new_n1245), .A4(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT58), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1246), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1203), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G125), .A2(new_n847), .B1(new_n983), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(G128), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1256), .B1(new_n1257), .B2(new_n774), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G150), .B2(new_n764), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n767), .A2(G137), .B1(new_n791), .B2(G132), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT121), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT59), .ZN(new_n1263));
  AOI211_X1 g1063(.A(G33), .B(G41), .C1(new_n855), .C2(G159), .ZN(new_n1264));
  INV_X1    g1064(.A(G124), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1264), .B1(new_n1265), .B2(new_n760), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1254), .B1(new_n1253), .B2(new_n1252), .C1(new_n1263), .C2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1244), .B1(new_n1267), .B2(new_n748), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1226), .B2(new_n750), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1243), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1242), .A2(new_n1271), .ZN(G375));
  AND2_X1   g1072(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1158), .A2(new_n749), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n736), .B1(new_n840), .B2(G68), .ZN(new_n1276));
  OAI221_X1 g1076(.A(new_n366), .B1(new_n202), .B2(new_n780), .C1(new_n992), .C2(new_n774), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n797), .A2(new_n334), .B1(new_n844), .B2(new_n776), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1277), .B(new_n1278), .C1(new_n791), .C2(new_n1255), .ZN(new_n1279));
  OAI221_X1 g1079(.A(new_n1279), .B1(new_n1257), .B2(new_n760), .C1(new_n395), .C2(new_n809), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n764), .A2(G50), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n805), .A2(G303), .ZN(new_n1282));
  OAI221_X1 g1082(.A(new_n1282), .B1(new_n489), .B2(new_n809), .C1(new_n770), .C2(new_n505), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n847), .A2(G294), .B1(new_n791), .B2(new_n549), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n796), .B2(new_n774), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1286), .A2(new_n1096), .A3(new_n407), .A4(new_n987), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n1280), .A2(new_n1281), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT123), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n746), .B2(new_n747), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1276), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1274), .A2(new_n734), .B1(new_n1275), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1273), .A2(new_n1179), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1072), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(new_n1186), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(G381));
  AOI22_X1  g1098(.A1(new_n1191), .A2(new_n1214), .B1(new_n1229), .B2(new_n1233), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n730), .B1(new_n1299), .B2(KEYINPUT57), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1240), .B1(new_n1299), .B2(KEYINPUT57), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1270), .B1(new_n1302), .B2(new_n1241), .ZN(new_n1303));
  INV_X1    g1103(.A(G378), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OR4_X1    g1105(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1306));
  NOR4_X1   g1106(.A1(new_n1305), .A2(G387), .A3(G381), .A4(new_n1306), .ZN(new_n1307));
  XOR2_X1   g1107(.A(new_n1307), .B(KEYINPUT124), .Z(G407));
  OAI211_X1 g1108(.A(G407), .B(G213), .C1(new_n663), .C2(new_n1305), .ZN(G409));
  NAND2_X1  g1109(.A1(new_n662), .A2(G213), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1231), .A2(new_n1232), .A3(new_n967), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n967), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT125), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1229), .A2(new_n1314), .A3(new_n1233), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n734), .A3(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1215), .A2(new_n1296), .A3(new_n1234), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1269), .A3(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1310), .B1(new_n1318), .B2(G378), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT60), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1295), .B1(new_n1321), .B2(new_n1185), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1273), .A2(KEYINPUT60), .A3(new_n1179), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(new_n730), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1294), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n867), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1324), .A2(G384), .A3(new_n1294), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1320), .B(new_n1329), .C1(new_n1303), .C2(new_n1304), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(G393), .B(new_n815), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(KEYINPUT113), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1077), .ZN(new_n1337));
  AOI21_X1  g1137(.A(G390), .B1(new_n1337), .B2(new_n1010), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1010), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1121), .A2(new_n1122), .A3(new_n1144), .ZN(new_n1340));
  AOI211_X1 g1140(.A(new_n1339), .B(new_n1340), .C1(new_n1336), .C2(new_n1077), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1334), .B1(new_n1338), .B2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(G387), .A2(new_n1340), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1337), .A2(new_n1010), .A3(G390), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1333), .A3(new_n1344), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1310), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(G2897), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(new_n1328), .B(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1304), .B1(new_n1242), .B2(new_n1271), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1349), .B1(new_n1350), .B2(new_n1319), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT61), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1332), .A2(new_n1346), .A3(new_n1351), .A4(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(G375), .A2(G378), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1354), .A2(KEYINPUT63), .A3(new_n1320), .A4(new_n1329), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT126), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1319), .B1(G375), .B2(G378), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1358), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1329), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1357), .A2(new_n1359), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1353), .A2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT62), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1362), .B1(new_n1358), .B2(new_n1329), .ZN(new_n1363));
  NOR4_X1   g1163(.A1(new_n1350), .A2(new_n1319), .A3(KEYINPUT62), .A4(new_n1328), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1354), .A2(new_n1320), .ZN(new_n1366));
  AOI21_X1  g1166(.A(KEYINPUT61), .B1(new_n1366), .B2(new_n1349), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1346), .B1(new_n1365), .B2(new_n1367), .ZN(new_n1368));
  OAI21_X1  g1168(.A(KEYINPUT127), .B1(new_n1361), .B2(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1348), .ZN(new_n1370));
  XNOR2_X1  g1170(.A(new_n1328), .B(new_n1370), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1358), .A2(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1373));
  NOR3_X1   g1173(.A1(new_n1372), .A2(new_n1373), .A3(KEYINPUT61), .ZN(new_n1374));
  NAND4_X1  g1174(.A1(new_n1374), .A2(new_n1332), .A3(new_n1357), .A4(new_n1359), .ZN(new_n1375));
  INV_X1    g1175(.A(new_n1364), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1330), .A2(KEYINPUT62), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1367), .A2(new_n1376), .A3(new_n1377), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1378), .A2(new_n1373), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT127), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1375), .A2(new_n1379), .A3(new_n1380), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1369), .A2(new_n1381), .ZN(G405));
  NAND2_X1  g1182(.A1(new_n1305), .A2(new_n1354), .ZN(new_n1383));
  XNOR2_X1  g1183(.A(new_n1383), .B(new_n1329), .ZN(new_n1384));
  XNOR2_X1  g1184(.A(new_n1384), .B(new_n1346), .ZN(G402));
endmodule


