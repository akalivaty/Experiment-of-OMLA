

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592;

  NOR2_X2 U323 ( .A1(n484), .A2(n423), .ZN(n424) );
  XNOR2_X2 U324 ( .A(n342), .B(n341), .ZN(n343) );
  INV_X1 U325 ( .A(KEYINPUT105), .ZN(n457) );
  XNOR2_X1 U326 ( .A(n420), .B(n419), .ZN(n540) );
  XOR2_X1 U327 ( .A(n380), .B(n330), .Z(n291) );
  XOR2_X1 U328 ( .A(n332), .B(KEYINPUT9), .Z(n292) );
  XNOR2_X1 U329 ( .A(n390), .B(n293), .ZN(n295) );
  XNOR2_X1 U330 ( .A(n475), .B(n474), .ZN(n476) );
  INV_X1 U331 ( .A(KEYINPUT72), .ZN(n302) );
  XNOR2_X1 U332 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U333 ( .A(n305), .B(n304), .ZN(n307) );
  XNOR2_X1 U334 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n480) );
  XNOR2_X1 U335 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U336 ( .A(n457), .B(KEYINPUT37), .ZN(n458) );
  XNOR2_X1 U337 ( .A(n411), .B(n410), .ZN(n416) );
  OR2_X1 U338 ( .A1(n563), .A2(n492), .ZN(n493) );
  XNOR2_X1 U339 ( .A(n459), .B(n458), .ZN(n536) );
  XNOR2_X1 U340 ( .A(n495), .B(n494), .ZN(n496) );
  INV_X1 U341 ( .A(G36GAT), .ZN(n461) );
  XNOR2_X1 U342 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U343 ( .A(n461), .B(KEYINPUT106), .ZN(n462) );
  XNOR2_X1 U344 ( .A(n491), .B(n490), .ZN(G1349GAT) );
  XNOR2_X1 U345 ( .A(n463), .B(n462), .ZN(G1329GAT) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G71GAT), .Z(n390) );
  AND2_X1 U347 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(G148GAT), .B(G106GAT), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n294), .B(G78GAT), .ZN(n372) );
  XNOR2_X1 U350 ( .A(n295), .B(n372), .ZN(n298) );
  INV_X1 U351 ( .A(n298), .ZN(n297) );
  INV_X1 U352 ( .A(KEYINPUT33), .ZN(n296) );
  NAND2_X1 U353 ( .A1(n297), .A2(n296), .ZN(n300) );
  NAND2_X1 U354 ( .A1(n298), .A2(KEYINPUT33), .ZN(n299) );
  NAND2_X1 U355 ( .A1(n300), .A2(n299), .ZN(n305) );
  XNOR2_X1 U356 ( .A(G85GAT), .B(KEYINPUT70), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n301), .B(G99GAT), .ZN(n333) );
  XOR2_X1 U358 ( .A(n333), .B(KEYINPUT32), .Z(n303) );
  XOR2_X1 U359 ( .A(G57GAT), .B(KEYINPUT13), .Z(n349) );
  XNOR2_X1 U360 ( .A(n349), .B(KEYINPUT31), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U362 ( .A(G204GAT), .B(KEYINPUT71), .Z(n309) );
  XNOR2_X1 U363 ( .A(G92GAT), .B(G176GAT), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U365 ( .A(G64GAT), .B(n310), .ZN(n417) );
  XNOR2_X1 U366 ( .A(n311), .B(n417), .ZN(n583) );
  XOR2_X1 U367 ( .A(KEYINPUT67), .B(G197GAT), .Z(n313) );
  XNOR2_X1 U368 ( .A(G15GAT), .B(KEYINPUT68), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U370 ( .A(G141GAT), .B(G22GAT), .Z(n379) );
  XOR2_X1 U371 ( .A(n314), .B(n379), .Z(n318) );
  XOR2_X1 U372 ( .A(G43GAT), .B(KEYINPUT8), .Z(n316) );
  XNOR2_X1 U373 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n316), .B(n315), .ZN(n340) );
  XOR2_X1 U375 ( .A(G8GAT), .B(G169GAT), .Z(n409) );
  XNOR2_X1 U376 ( .A(n340), .B(n409), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U378 ( .A(n319), .B(G50GAT), .Z(n321) );
  XOR2_X1 U379 ( .A(G113GAT), .B(G1GAT), .Z(n436) );
  XNOR2_X1 U380 ( .A(n436), .B(G36GAT), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n321), .B(n320), .ZN(n326) );
  XOR2_X1 U382 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n323) );
  NAND2_X1 U383 ( .A1(G229GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U385 ( .A(KEYINPUT29), .B(n324), .Z(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n577) );
  NAND2_X1 U387 ( .A1(n583), .A2(n577), .ZN(n327) );
  XNOR2_X1 U388 ( .A(KEYINPUT73), .B(n327), .ZN(n503) );
  XOR2_X1 U389 ( .A(G162GAT), .B(G50GAT), .Z(n380) );
  XOR2_X1 U390 ( .A(KEYINPUT11), .B(G92GAT), .Z(n329) );
  XNOR2_X1 U391 ( .A(G218GAT), .B(KEYINPUT74), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n330) );
  NAND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n291), .B(n331), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(KEYINPUT10), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n292), .B(n334), .ZN(n338) );
  XOR2_X1 U397 ( .A(KEYINPUT65), .B(KEYINPUT75), .Z(n336) );
  XNOR2_X1 U398 ( .A(G134GAT), .B(G106GAT), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n338), .B(n337), .ZN(n342) );
  XNOR2_X1 U401 ( .A(G36GAT), .B(KEYINPUT76), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n339), .B(G190GAT), .ZN(n412) );
  XNOR2_X1 U403 ( .A(n412), .B(n340), .ZN(n341) );
  INV_X1 U404 ( .A(n343), .ZN(n499) );
  XOR2_X1 U405 ( .A(KEYINPUT36), .B(n499), .Z(n589) );
  XOR2_X1 U406 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n345) );
  XNOR2_X1 U407 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n353) );
  XOR2_X1 U409 ( .A(G183GAT), .B(G71GAT), .Z(n347) );
  XNOR2_X1 U410 ( .A(G78GAT), .B(G211GAT), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U412 ( .A(n348), .B(G22GAT), .Z(n351) );
  XNOR2_X1 U413 ( .A(G155GAT), .B(n349), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n366) );
  XOR2_X1 U416 ( .A(G8GAT), .B(KEYINPUT68), .Z(n355) );
  XNOR2_X1 U417 ( .A(G1GAT), .B(G64GAT), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U419 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n357) );
  XNOR2_X1 U420 ( .A(KEYINPUT15), .B(KEYINPUT77), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U422 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U423 ( .A(G127GAT), .B(G15GAT), .Z(n397) );
  XOR2_X1 U424 ( .A(KEYINPUT83), .B(KEYINPUT12), .Z(n361) );
  NAND2_X1 U425 ( .A1(G231GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n397), .B(n362), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n366), .B(n365), .ZN(n587) );
  XOR2_X1 U430 ( .A(KEYINPUT88), .B(KEYINPUT91), .Z(n368) );
  NAND2_X1 U431 ( .A1(G228GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U433 ( .A(n369), .B(KEYINPUT24), .Z(n374) );
  XOR2_X1 U434 ( .A(G155GAT), .B(KEYINPUT3), .Z(n371) );
  XNOR2_X1 U435 ( .A(KEYINPUT90), .B(KEYINPUT2), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n371), .B(n370), .ZN(n445) );
  XNOR2_X1 U437 ( .A(n445), .B(n372), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U439 ( .A(KEYINPUT22), .B(KEYINPUT92), .Z(n376) );
  XNOR2_X1 U440 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U442 ( .A(n378), .B(n377), .Z(n382) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n387) );
  XOR2_X1 U445 ( .A(KEYINPUT89), .B(G197GAT), .Z(n384) );
  XNOR2_X1 U446 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U448 ( .A(G211GAT), .B(n385), .Z(n411) );
  INV_X1 U449 ( .A(n411), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n387), .B(n386), .ZN(n484) );
  XOR2_X1 U451 ( .A(KEYINPUT20), .B(G99GAT), .Z(n389) );
  XNOR2_X1 U452 ( .A(G190GAT), .B(G43GAT), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n391) );
  XOR2_X1 U454 ( .A(n391), .B(n390), .Z(n396) );
  XOR2_X1 U455 ( .A(G134GAT), .B(KEYINPUT0), .Z(n437) );
  XOR2_X1 U456 ( .A(KEYINPUT18), .B(KEYINPUT85), .Z(n393) );
  XNOR2_X1 U457 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n392) );
  XNOR2_X1 U458 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U459 ( .A(G183GAT), .B(n394), .Z(n418) );
  XNOR2_X1 U460 ( .A(n437), .B(n418), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n396), .B(n395), .ZN(n401) );
  XOR2_X1 U462 ( .A(n397), .B(G169GAT), .Z(n399) );
  NAND2_X1 U463 ( .A1(G227GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U465 ( .A(n401), .B(n400), .Z(n406) );
  XOR2_X1 U466 ( .A(G176GAT), .B(KEYINPUT84), .Z(n403) );
  XNOR2_X1 U467 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U469 ( .A(G113GAT), .B(n404), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n451) );
  NAND2_X1 U471 ( .A1(n484), .A2(n451), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n407), .B(KEYINPUT26), .ZN(n563) );
  XOR2_X1 U473 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n408) );
  XOR2_X1 U474 ( .A(n412), .B(KEYINPUT97), .Z(n414) );
  NAND2_X1 U475 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U477 ( .A(n416), .B(n415), .Z(n420) );
  XOR2_X1 U478 ( .A(n418), .B(n417), .Z(n419) );
  XNOR2_X1 U479 ( .A(n540), .B(KEYINPUT27), .ZN(n452) );
  NOR2_X1 U480 ( .A1(n563), .A2(n452), .ZN(n421) );
  XOR2_X1 U481 ( .A(KEYINPUT100), .B(n421), .Z(n426) );
  NOR2_X1 U482 ( .A1(n451), .A2(n540), .ZN(n422) );
  XOR2_X1 U483 ( .A(KEYINPUT101), .B(n422), .Z(n423) );
  XNOR2_X1 U484 ( .A(KEYINPUT25), .B(n424), .ZN(n425) );
  NAND2_X1 U485 ( .A1(n426), .A2(n425), .ZN(n427) );
  XNOR2_X1 U486 ( .A(KEYINPUT102), .B(n427), .ZN(n450) );
  XOR2_X1 U487 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n429) );
  XNOR2_X1 U488 ( .A(G120GAT), .B(G57GAT), .ZN(n428) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U490 ( .A(G127GAT), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U491 ( .A(G162GAT), .B(G141GAT), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n449) );
  XOR2_X1 U494 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n435) );
  XNOR2_X1 U495 ( .A(KEYINPUT5), .B(KEYINPUT93), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n441) );
  XOR2_X1 U497 ( .A(G85GAT), .B(n436), .Z(n439) );
  XNOR2_X1 U498 ( .A(G29GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U500 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U501 ( .A1(G225GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U503 ( .A(n444), .B(KEYINPUT6), .Z(n447) );
  XNOR2_X1 U504 ( .A(n445), .B(KEYINPUT96), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n537) );
  NAND2_X1 U507 ( .A1(n450), .A2(n537), .ZN(n454) );
  OR2_X1 U508 ( .A1(n452), .A2(n537), .ZN(n565) );
  XNOR2_X1 U509 ( .A(n484), .B(KEYINPUT28), .ZN(n510) );
  NOR2_X1 U510 ( .A1(n565), .A2(n510), .ZN(n550) );
  NAND2_X1 U511 ( .A1(n451), .A2(n550), .ZN(n453) );
  NAND2_X1 U512 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n455), .B(KEYINPUT103), .ZN(n502) );
  NOR2_X1 U514 ( .A1(n587), .A2(n502), .ZN(n456) );
  NAND2_X1 U515 ( .A1(n589), .A2(n456), .ZN(n459) );
  NAND2_X1 U516 ( .A1(n503), .A2(n536), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n460), .B(KEYINPUT38), .ZN(n518) );
  NOR2_X1 U518 ( .A1(n518), .A2(n540), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n583), .B(KEYINPUT41), .ZN(n570) );
  XNOR2_X1 U520 ( .A(KEYINPUT110), .B(n570), .ZN(n553) );
  AND2_X1 U521 ( .A1(n577), .A2(n570), .ZN(n465) );
  INV_X1 U522 ( .A(KEYINPUT46), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n465), .B(n464), .ZN(n467) );
  NOR2_X1 U524 ( .A1(n587), .A2(n343), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n469) );
  XOR2_X1 U526 ( .A(KEYINPUT117), .B(KEYINPUT47), .Z(n468) );
  NAND2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n473) );
  INV_X1 U528 ( .A(n468), .ZN(n471) );
  INV_X1 U529 ( .A(n469), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n479) );
  NAND2_X1 U532 ( .A1(n589), .A2(n587), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n474) );
  NAND2_X1 U534 ( .A1(n583), .A2(n476), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n577), .A2(n477), .ZN(n478) );
  NOR2_X1 U536 ( .A1(n479), .A2(n478), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(n480), .ZN(n548) );
  NOR2_X1 U538 ( .A1(n548), .A2(n540), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n482), .B(KEYINPUT54), .ZN(n483) );
  NAND2_X1 U540 ( .A1(n483), .A2(n537), .ZN(n492) );
  NOR2_X1 U541 ( .A1(n492), .A2(n484), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(KEYINPUT55), .ZN(n486) );
  NOR2_X1 U543 ( .A1(n451), .A2(n486), .ZN(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT123), .B(n487), .Z(n580) );
  NAND2_X1 U545 ( .A1(n553), .A2(n580), .ZN(n491) );
  XOR2_X1 U546 ( .A(G176GAT), .B(KEYINPUT56), .Z(n489) );
  XNOR2_X1 U547 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT125), .B(n493), .ZN(n590) );
  NAND2_X1 U549 ( .A1(n590), .A2(n577), .ZN(n495) );
  XOR2_X1 U550 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n494) );
  XNOR2_X1 U551 ( .A(n496), .B(KEYINPUT59), .ZN(n498) );
  XOR2_X1 U552 ( .A(G197GAT), .B(KEYINPUT126), .Z(n497) );
  XNOR2_X1 U553 ( .A(n498), .B(n497), .ZN(G1352GAT) );
  NAND2_X1 U554 ( .A1(n499), .A2(n587), .ZN(n500) );
  XNOR2_X1 U555 ( .A(KEYINPUT16), .B(n500), .ZN(n501) );
  NOR2_X1 U556 ( .A1(n502), .A2(n501), .ZN(n522) );
  NAND2_X1 U557 ( .A1(n503), .A2(n522), .ZN(n511) );
  NOR2_X1 U558 ( .A1(n537), .A2(n511), .ZN(n505) );
  XNOR2_X1 U559 ( .A(KEYINPUT34), .B(KEYINPUT104), .ZN(n504) );
  XNOR2_X1 U560 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U561 ( .A(G1GAT), .B(n506), .Z(G1324GAT) );
  NOR2_X1 U562 ( .A1(n540), .A2(n511), .ZN(n507) );
  XOR2_X1 U563 ( .A(G8GAT), .B(n507), .Z(G1325GAT) );
  NOR2_X1 U564 ( .A1(n451), .A2(n511), .ZN(n509) );
  XNOR2_X1 U565 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n508) );
  XNOR2_X1 U566 ( .A(n509), .B(n508), .ZN(G1326GAT) );
  INV_X1 U567 ( .A(n510), .ZN(n544) );
  NOR2_X1 U568 ( .A1(n544), .A2(n511), .ZN(n512) );
  XOR2_X1 U569 ( .A(G22GAT), .B(n512), .Z(G1327GAT) );
  NOR2_X1 U570 ( .A1(n537), .A2(n518), .ZN(n513) );
  XNOR2_X1 U571 ( .A(G29GAT), .B(n513), .ZN(n514) );
  XNOR2_X1 U572 ( .A(n514), .B(KEYINPUT39), .ZN(G1328GAT) );
  XNOR2_X1 U573 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n516) );
  NOR2_X1 U574 ( .A1(n451), .A2(n518), .ZN(n515) );
  XNOR2_X1 U575 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U576 ( .A(G43GAT), .B(n517), .ZN(G1330GAT) );
  NOR2_X1 U577 ( .A1(n544), .A2(n518), .ZN(n519) );
  XOR2_X1 U578 ( .A(KEYINPUT108), .B(n519), .Z(n520) );
  XNOR2_X1 U579 ( .A(G50GAT), .B(n520), .ZN(G1331GAT) );
  INV_X1 U580 ( .A(n553), .ZN(n521) );
  NOR2_X1 U581 ( .A1(n577), .A2(n521), .ZN(n535) );
  NAND2_X1 U582 ( .A1(n535), .A2(n522), .ZN(n531) );
  NOR2_X1 U583 ( .A1(n531), .A2(n537), .ZN(n526) );
  XOR2_X1 U584 ( .A(KEYINPUT109), .B(KEYINPUT111), .Z(n524) );
  XNOR2_X1 U585 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n526), .B(n525), .ZN(G1332GAT) );
  NOR2_X1 U588 ( .A1(n540), .A2(n531), .ZN(n527) );
  XOR2_X1 U589 ( .A(KEYINPUT112), .B(n527), .Z(n528) );
  XNOR2_X1 U590 ( .A(G64GAT), .B(n528), .ZN(G1333GAT) );
  NOR2_X1 U591 ( .A1(n451), .A2(n531), .ZN(n530) );
  XNOR2_X1 U592 ( .A(G71GAT), .B(KEYINPUT113), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(G1334GAT) );
  NOR2_X1 U594 ( .A1(n544), .A2(n531), .ZN(n533) );
  XNOR2_X1 U595 ( .A(KEYINPUT43), .B(KEYINPUT114), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U597 ( .A(G78GAT), .B(n534), .ZN(G1335GAT) );
  NAND2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n543) );
  NOR2_X1 U599 ( .A1(n537), .A2(n543), .ZN(n539) );
  XNOR2_X1 U600 ( .A(G85GAT), .B(KEYINPUT115), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n539), .B(n538), .ZN(G1336GAT) );
  NOR2_X1 U602 ( .A1(n540), .A2(n543), .ZN(n541) );
  XOR2_X1 U603 ( .A(G92GAT), .B(n541), .Z(G1337GAT) );
  NOR2_X1 U604 ( .A1(n451), .A2(n543), .ZN(n542) );
  XOR2_X1 U605 ( .A(G99GAT), .B(n542), .Z(G1338GAT) );
  NOR2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U607 ( .A(KEYINPUT44), .B(KEYINPUT116), .ZN(n545) );
  XNOR2_X1 U608 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U609 ( .A(G106GAT), .B(n547), .Z(G1339GAT) );
  INV_X1 U610 ( .A(n451), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U612 ( .A1(n548), .A2(n551), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n559), .A2(n577), .ZN(n552) );
  XNOR2_X1 U614 ( .A(G113GAT), .B(n552), .ZN(G1340GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n555) );
  NAND2_X1 U616 ( .A1(n559), .A2(n553), .ZN(n554) );
  XNOR2_X1 U617 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U618 ( .A(G120GAT), .B(n556), .ZN(G1341GAT) );
  NAND2_X1 U619 ( .A1(n559), .A2(n587), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n557), .B(KEYINPUT50), .ZN(n558) );
  XNOR2_X1 U621 ( .A(G127GAT), .B(n558), .ZN(G1342GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n561) );
  NAND2_X1 U623 ( .A1(n559), .A2(n343), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U625 ( .A(G134GAT), .B(n562), .Z(G1343GAT) );
  OR2_X1 U626 ( .A1(n563), .A2(n548), .ZN(n564) );
  NOR2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n575) );
  NAND2_X1 U628 ( .A1(n577), .A2(n575), .ZN(n566) );
  XNOR2_X1 U629 ( .A(n566), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n568) );
  XNOR2_X1 U631 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT53), .B(n569), .Z(n572) );
  NAND2_X1 U634 ( .A1(n575), .A2(n570), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n572), .B(n571), .ZN(G1345GAT) );
  NAND2_X1 U636 ( .A1(n575), .A2(n587), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(KEYINPUT122), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G155GAT), .B(n574), .ZN(G1346GAT) );
  NAND2_X1 U639 ( .A1(n343), .A2(n575), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n580), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U643 ( .A1(n580), .A2(n587), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U645 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n343), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1351GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  INV_X1 U649 ( .A(n583), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n590), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n590), .A2(n587), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

