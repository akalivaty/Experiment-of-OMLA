//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1273, new_n1274;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G125), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT67), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n469), .B2(new_n461), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n463), .A2(G137), .A3(new_n465), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n463), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n465), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n467), .A2(new_n468), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(G136), .B2(new_n488), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT68), .Z(G162));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n465), .B2(G114), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n492), .A2(new_n494), .A3(new_n495), .A4(G2104), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n467), .B2(new_n468), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n500), .B(new_n503), .C1(new_n468), .C2(new_n467), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n498), .B1(new_n502), .B2(new_n504), .ZN(G164));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n512), .A2(new_n513), .B1(new_n506), .B2(new_n507), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n515), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n509), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n513), .A2(new_n512), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n508), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n527), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT70), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(new_n538), .A3(G651), .ZN(new_n539));
  INV_X1    g114(.A(new_n514), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n506), .A2(new_n507), .ZN(new_n541));
  INV_X1    g116(.A(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(G90), .A2(new_n540), .B1(new_n543), .B2(G52), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n537), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(G171));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n528), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT71), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(KEYINPUT71), .ZN(new_n552));
  AOI22_X1  g127(.A1(G81), .A2(new_n540), .B1(new_n543), .B2(G43), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g132(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n558));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n528), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n566), .B2(new_n514), .ZN(new_n567));
  OAI211_X1 g142(.A(G53), .B(G543), .C1(new_n506), .C2(new_n507), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n508), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT73), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n567), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G299));
  XNOR2_X1  g153(.A(new_n545), .B(KEYINPUT74), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n514), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n508), .A2(KEYINPUT75), .A3(G87), .A4(new_n518), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n583), .A2(new_n584), .B1(G49), .B2(new_n543), .ZN(new_n585));
  NOR3_X1   g160(.A1(new_n513), .A2(new_n512), .A3(G74), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT76), .B1(new_n586), .B2(new_n520), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n588), .B(G651), .C1(new_n518), .C2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n585), .A2(new_n590), .ZN(G288));
  OAI211_X1 g166(.A(G48), .B(G543), .C1(new_n506), .C2(new_n507), .ZN(new_n592));
  INV_X1    g167(.A(G86), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n514), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(G61), .B1(new_n513), .B2(new_n512), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n540), .A2(G85), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n543), .A2(G47), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n601), .B(new_n602), .C1(new_n520), .C2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT77), .Z(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n528), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n606), .B(KEYINPUT78), .C1(new_n607), .C2(new_n528), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n610), .A2(G651), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n540), .A2(KEYINPUT10), .A3(G92), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n514), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n613), .A2(new_n616), .B1(G54), .B2(new_n543), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G301), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G284));
  AOI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n577), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(new_n577), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(new_n618), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n554), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n618), .A2(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n629), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n463), .A2(new_n476), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT13), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n482), .A2(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n465), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT80), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n488), .A2(new_n643), .A3(G135), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(new_n488), .B2(G135), .ZN(new_n645));
  OAI221_X1 g220(.A(new_n640), .B1(new_n641), .B2(new_n642), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n638), .A2(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(G2096), .ZN(new_n649));
  NAND4_X1  g224(.A1(new_n639), .A2(new_n647), .A3(new_n648), .A4(new_n649), .ZN(G156));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n654), .B2(new_n653), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(G401));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT81), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n668), .B(KEYINPUT17), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n673), .B(new_n670), .C1(new_n667), .C2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n667), .A3(new_n669), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n681), .B2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  XNOR2_X1  g271(.A(KEYINPUT91), .B(KEYINPUT25), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(G115), .A2(G2104), .ZN(new_n700));
  INV_X1    g275(.A(G127), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n487), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G2105), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n488), .A2(G139), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n699), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(KEYINPUT92), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n699), .A2(new_n703), .A3(new_n707), .A4(new_n704), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G33), .B(new_n709), .S(G29), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(new_n443), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n476), .A2(G105), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT94), .ZN(new_n713));
  INV_X1    g288(.A(G141), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n463), .A2(new_n465), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT26), .Z(new_n718));
  INV_X1    g293(.A(G129), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n481), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n722), .B2(G32), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G2084), .ZN(new_n727));
  AND2_X1   g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  NOR2_X1   g303(.A1(KEYINPUT24), .A2(G34), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n722), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT93), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n479), .B2(new_n722), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n711), .B(new_n726), .C1(new_n727), .C2(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT95), .Z(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT82), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT82), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(G19), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n555), .B2(new_n738), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1341), .ZN(new_n741));
  NOR2_X1   g316(.A1(G5), .A2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT96), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n545), .B2(new_n735), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n722), .A2(G26), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT28), .Z(new_n748));
  INV_X1    g323(.A(G128), .ZN(new_n749));
  OAI21_X1  g324(.A(KEYINPUT89), .B1(new_n481), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT89), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n463), .A2(new_n751), .A3(G128), .A4(G2105), .ZN(new_n752));
  NOR2_X1   g327(.A1(G104), .A2(G2105), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT90), .Z(new_n754));
  INV_X1    g329(.A(G116), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n475), .B1(new_n755), .B2(G2105), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n750), .A2(new_n752), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n488), .A2(new_n758), .A3(G140), .ZN(new_n759));
  INV_X1    g334(.A(G140), .ZN(new_n760));
  OAI21_X1  g335(.A(KEYINPUT88), .B1(new_n715), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n748), .B1(new_n763), .B2(G29), .ZN(new_n764));
  INV_X1    g339(.A(G2067), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n741), .A2(new_n746), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n722), .A2(G35), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G162), .B2(new_n722), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT29), .B(G2090), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n626), .A2(new_n735), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G4), .B2(new_n735), .ZN(new_n773));
  INV_X1    g348(.A(G1348), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n732), .A2(new_n727), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n738), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G20), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT23), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n577), .B2(new_n735), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1956), .ZN(new_n783));
  NOR2_X1   g358(.A1(G168), .A2(new_n735), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n735), .B2(G21), .ZN(new_n785));
  INV_X1    g360(.A(G1966), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n724), .B2(new_n725), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT30), .B(G28), .ZN(new_n789));
  OR2_X1    g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  NAND2_X1  g365(.A1(KEYINPUT31), .A2(G11), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n789), .A2(new_n722), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n504), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n503), .B1(new_n463), .B2(new_n500), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n497), .B(new_n496), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G29), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n722), .A2(G27), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n792), .B1(new_n646), .B2(new_n722), .C1(new_n798), .C2(new_n444), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n444), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n785), .B2(new_n786), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n788), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n771), .A2(new_n778), .A3(new_n783), .A4(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n734), .A2(new_n767), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n738), .A2(G22), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G166), .B2(new_n738), .ZN(new_n806));
  INV_X1    g381(.A(G1971), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n735), .A2(G23), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G288), .B2(G16), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT33), .B(G1976), .Z(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n810), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n735), .A2(G6), .ZN(new_n815));
  INV_X1    g390(.A(G305), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n735), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT32), .B(G1981), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT84), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n808), .A2(new_n813), .A3(new_n814), .A4(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT85), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT34), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n779), .A2(G24), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT83), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G290), .B2(new_n738), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(G1986), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n722), .A2(G25), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n463), .A2(G131), .A3(new_n465), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n463), .A2(G119), .A3(G2105), .ZN(new_n830));
  OR2_X1    g405(.A1(G95), .A2(G2105), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n831), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n828), .B1(new_n834), .B2(new_n722), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT35), .B(G1991), .Z(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n835), .B(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n827), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n823), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT85), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n821), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT34), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT36), .B1(new_n840), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT86), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT86), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(KEYINPUT36), .C1(new_n840), .C2(new_n845), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n844), .A2(new_n823), .A3(new_n851), .A4(new_n839), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT87), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n804), .B1(new_n850), .B2(new_n854), .ZN(G311));
  NAND2_X1  g430(.A1(new_n850), .A2(new_n854), .ZN(new_n856));
  INV_X1    g431(.A(new_n804), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(G150));
  INV_X1    g433(.A(G55), .ZN(new_n859));
  INV_X1    g434(.A(G93), .ZN(new_n860));
  OAI22_X1  g435(.A1(new_n509), .A2(new_n859), .B1(new_n860), .B2(new_n514), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n520), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT97), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n555), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n554), .A2(new_n865), .A3(KEYINPUT97), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT38), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n626), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n876));
  XOR2_X1   g451(.A(KEYINPUT98), .B(G860), .Z(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n864), .A2(new_n877), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(G145));
  NOR2_X1   g456(.A1(new_n709), .A2(KEYINPUT100), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n706), .B2(new_n708), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n795), .A2(KEYINPUT99), .ZN(new_n886));
  INV_X1    g461(.A(new_n498), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n502), .A2(new_n504), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(new_n763), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n886), .A2(new_n890), .B1(new_n757), .B2(new_n762), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n892), .A2(new_n721), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n721), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n763), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n886), .A2(new_n762), .A3(new_n757), .A4(new_n890), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n885), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n721), .B1(new_n892), .B2(new_n893), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n895), .A3(new_n897), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n884), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n488), .A2(G142), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n463), .A2(G130), .A3(G2105), .ZN(new_n905));
  OR2_X1    g480(.A1(G106), .A2(G2105), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n906), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n834), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n908), .A2(new_n834), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT101), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n908), .A2(new_n834), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n914), .A3(new_n909), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n636), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n912), .A2(new_n915), .A3(new_n636), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n903), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT102), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n903), .A2(new_n924), .A3(new_n920), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI221_X4 g501(.A(KEYINPUT102), .B1(new_n919), .B2(new_n918), .C1(new_n899), .C2(new_n902), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n924), .B1(new_n903), .B2(new_n920), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT103), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n903), .A2(new_n920), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n926), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n646), .B(new_n479), .ZN(new_n933));
  XNOR2_X1  g508(.A(G162), .B(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n922), .A2(new_n925), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n935), .A2(new_n930), .ZN(new_n938));
  AOI21_X1  g513(.A(G37), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n936), .A2(KEYINPUT104), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT104), .B1(new_n936), .B2(new_n939), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT40), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n936), .A2(new_n939), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n936), .A2(KEYINPUT104), .A3(new_n939), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT40), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n943), .A2(new_n948), .ZN(G395));
  XNOR2_X1  g524(.A(G290), .B(KEYINPUT105), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(G288), .ZN(new_n951));
  XNOR2_X1  g526(.A(G303), .B(new_n816), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n954), .A2(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(KEYINPUT106), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n957));
  OR3_X1    g532(.A1(new_n953), .A2(new_n957), .A3(KEYINPUT42), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n953), .B2(KEYINPUT42), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n955), .A2(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n871), .B(new_n631), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n618), .B(new_n577), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n962), .A2(KEYINPUT41), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(KEYINPUT41), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n962), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n966), .B2(new_n961), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n960), .A2(KEYINPUT108), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n960), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(G868), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(G868), .B2(new_n864), .ZN(G295));
  OAI21_X1  g548(.A(new_n972), .B1(G868), .B2(new_n864), .ZN(G331));
  NOR2_X1   g549(.A1(G301), .A2(G286), .ZN(new_n975));
  NOR2_X1   g550(.A1(G171), .A2(G168), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n871), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n870), .B(new_n869), .C1(new_n975), .C2(new_n976), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n962), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n978), .A2(new_n964), .A3(new_n979), .A4(new_n963), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n953), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G37), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n953), .B1(new_n981), .B2(new_n982), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT43), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n983), .A2(new_n984), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n986), .A2(KEYINPUT109), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n990));
  AOI211_X1 g565(.A(new_n990), .B(new_n953), .C1(new_n981), .C2(new_n982), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(new_n992), .B2(KEYINPUT43), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n985), .B2(new_n986), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n992), .B2(new_n994), .ZN(new_n996));
  MUX2_X1   g571(.A(new_n993), .B(new_n996), .S(KEYINPUT44), .Z(G397));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n886), .A2(new_n998), .A3(new_n890), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n886), .A2(KEYINPUT110), .A3(new_n998), .A4(new_n890), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n474), .A2(G40), .A3(new_n477), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n469), .A2(new_n461), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n471), .B1(new_n1006), .B2(G2105), .ZN(new_n1007));
  AOI211_X1 g582(.A(KEYINPUT67), .B(new_n465), .C1(new_n469), .C2(new_n461), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(G1986), .A3(G290), .ZN(new_n1011));
  NOR2_X1   g586(.A1(G290), .A2(G1986), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT111), .Z(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n1015), .B(KEYINPUT112), .Z(new_n1016));
  XNOR2_X1  g591(.A(new_n1010), .B(KEYINPUT113), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n833), .A2(new_n837), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n834), .A2(new_n836), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1996), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1010), .A2(new_n1021), .A3(new_n721), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n763), .B(new_n765), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n1021), .B2(new_n721), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1020), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1016), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n474), .A2(G40), .A3(new_n477), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n466), .B2(new_n472), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n795), .A2(new_n1031), .A3(new_n998), .ZN(new_n1032));
  AND4_X1   g607(.A1(new_n727), .A2(new_n1028), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT45), .B1(new_n795), .B2(new_n998), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT117), .B1(new_n1034), .B2(new_n1009), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1384), .B1(new_n887), .B2(new_n888), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1030), .B(new_n1036), .C1(new_n1037), .C2(KEYINPUT45), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1002), .A2(G1384), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n795), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1033), .B1(new_n1041), .B2(new_n786), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G286), .A2(G8), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT51), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1043), .B(new_n1047), .C1(new_n1042), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1048), .B(new_n1047), .C1(new_n1042), .C2(G168), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1044), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n886), .A2(new_n890), .A3(new_n1039), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n795), .A2(new_n998), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1002), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1053), .A2(new_n1055), .A3(new_n444), .A4(new_n1030), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n745), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1057), .A2(G2078), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1035), .A2(new_n1061), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1058), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(KEYINPUT124), .A3(new_n620), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT124), .B1(new_n1063), .B2(new_n620), .ZN(new_n1066));
  NOR4_X1   g641(.A1(new_n1029), .A2(new_n470), .A3(new_n1057), .A4(G2078), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1053), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1004), .A2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1056), .A2(new_n1057), .B1(new_n745), .B2(new_n1059), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1069), .A2(new_n1070), .A3(G301), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1065), .A2(new_n1066), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1052), .B1(new_n1072), .B2(KEYINPUT54), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G303), .A2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G2090), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT116), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1031), .B1(new_n795), .B2(new_n998), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n1009), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1079), .B(new_n1032), .C1(new_n1080), .C2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1034), .A2(new_n1009), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1971), .B1(new_n1085), .B2(new_n1053), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1078), .B1(new_n1088), .B2(G8), .ZN(new_n1089));
  AND4_X1   g664(.A1(new_n1079), .A2(new_n1028), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1078), .B(G8), .C1(new_n1086), .C2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1048), .B1(new_n1030), .B2(new_n1037), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n585), .A2(KEYINPUT114), .A3(G1976), .A4(new_n590), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n583), .A2(new_n584), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n543), .A2(G49), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1094), .A2(new_n590), .A3(G1976), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1092), .A2(new_n1093), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1976), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT52), .B1(G288), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(G8), .B1(new_n1054), .B2(new_n1009), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n508), .A2(G86), .A3(new_n518), .ZN(new_n1103));
  INV_X1    g678(.A(G1981), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n599), .A2(new_n1103), .A3(new_n1104), .A4(new_n592), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n520), .B1(new_n596), .B2(new_n597), .ZN(new_n1106));
  OAI21_X1  g681(.A(G1981), .B1(new_n594), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT49), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1105), .A2(new_n1107), .A3(KEYINPUT49), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT115), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1105), .A2(new_n1107), .A3(new_n1112), .A4(KEYINPUT49), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1099), .A2(new_n1101), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1092), .A2(new_n1098), .A3(new_n1093), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT52), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1091), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT125), .B1(new_n1089), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1078), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1032), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1082), .B1(new_n1081), .B2(new_n1009), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1030), .B(KEYINPUT116), .C1(new_n1037), .C2(new_n1031), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1086), .B1(new_n1124), .B2(new_n1079), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1120), .B1(new_n1125), .B2(new_n1048), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1101), .A2(new_n1093), .A3(new_n1092), .A4(new_n1098), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1128), .A2(new_n1117), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1126), .A2(new_n1127), .A3(new_n1091), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1070), .A2(G301), .A3(new_n1062), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1133));
  OAI211_X1 g708(.A(KEYINPUT54), .B(new_n1132), .C1(new_n1133), .C2(new_n545), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1119), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT126), .B1(new_n1073), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1063), .A2(new_n620), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1069), .A2(new_n1070), .A3(G301), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(new_n1064), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1047), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1041), .A2(new_n786), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1033), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g721(.A(G8), .B(new_n1143), .C1(new_n1146), .C2(G286), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1049), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1141), .A2(new_n1142), .B1(new_n1148), .B2(new_n1044), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1119), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI22_X1  g727(.A1(G651), .A2(new_n564), .B1(new_n540), .B2(G91), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n575), .A2(KEYINPUT73), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT57), .B(new_n1153), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT120), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n577), .A2(new_n1158), .A3(KEYINPUT57), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n567), .B2(new_n570), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT56), .B(G2072), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1085), .A2(new_n1053), .A3(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1163), .B(new_n1165), .C1(G1956), .C2(new_n1124), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1124), .B2(G1956), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT61), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1059), .A2(new_n774), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1054), .A2(new_n1009), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n765), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(KEYINPUT60), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n618), .A2(KEYINPUT122), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1059), .A2(new_n774), .B1(new_n1172), .B2(new_n765), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n618), .A2(KEYINPUT122), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1178), .A2(new_n1179), .A3(KEYINPUT60), .A4(new_n1175), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1059), .A2(new_n774), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1173), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1177), .A2(new_n1180), .A3(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1085), .A2(new_n1021), .A3(new_n1053), .ZN(new_n1186));
  XOR2_X1   g761(.A(KEYINPUT58), .B(G1341), .Z(new_n1187));
  OAI21_X1  g762(.A(new_n1187), .B1(new_n1054), .B2(new_n1009), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n555), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1189), .A2(KEYINPUT59), .A3(new_n555), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1185), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1170), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT121), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1169), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1167), .A2(new_n1168), .A3(KEYINPUT121), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1197), .A2(KEYINPUT61), .A3(new_n1198), .A4(new_n1166), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n626), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1197), .A2(new_n1201), .A3(new_n1198), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(new_n1166), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1136), .A2(new_n1152), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1206), .A2(new_n1091), .ZN(new_n1207));
  NOR2_X1   g782(.A1(G288), .A2(G1976), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1128), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1102), .B1(new_n1209), .B2(new_n1105), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1089), .A2(new_n1118), .ZN(new_n1214));
  NOR3_X1   g789(.A1(new_n1042), .A2(new_n1048), .A3(G286), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1213), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1042), .A2(new_n1048), .ZN(new_n1217));
  NAND4_X1  g792(.A1(new_n1217), .A2(KEYINPUT63), .A3(G168), .A4(new_n1091), .ZN(new_n1218));
  OAI21_X1  g793(.A(G8), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1219));
  AND2_X1   g794(.A1(new_n1219), .A2(new_n1120), .ZN(new_n1220));
  OAI21_X1  g795(.A(KEYINPUT119), .B1(new_n1220), .B2(new_n1206), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1219), .A2(new_n1120), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT119), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1130), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1218), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1211), .B1(new_n1216), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT62), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1148), .A2(new_n1227), .A3(new_n1044), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1227), .B1(new_n1148), .B2(new_n1044), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1139), .A2(new_n1064), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1119), .A2(new_n1230), .A3(new_n1131), .ZN(new_n1231));
  NOR2_X1   g806(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1226), .B1(new_n1228), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1027), .B1(new_n1205), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1023), .A2(new_n721), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1017), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1010), .A2(new_n1021), .ZN(new_n1237));
  XNOR2_X1  g812(.A(new_n1237), .B(KEYINPUT46), .ZN(new_n1238));
  INV_X1    g813(.A(KEYINPUT47), .ZN(new_n1239));
  AND3_X1   g814(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g815(.A(new_n1239), .B1(new_n1238), .B2(new_n1236), .ZN(new_n1241));
  XNOR2_X1  g816(.A(new_n1014), .B(KEYINPUT48), .ZN(new_n1242));
  INV_X1    g817(.A(new_n1242), .ZN(new_n1243));
  OAI22_X1  g818(.A1(new_n1240), .A2(new_n1241), .B1(new_n1026), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g819(.A(new_n1017), .ZN(new_n1245));
  NAND3_X1  g820(.A1(new_n1025), .A2(new_n1022), .A3(new_n1018), .ZN(new_n1246));
  NAND3_X1  g821(.A1(new_n757), .A2(new_n765), .A3(new_n762), .ZN(new_n1247));
  AOI21_X1  g822(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g823(.A1(new_n1244), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g824(.A(new_n1249), .ZN(new_n1250));
  OAI21_X1  g825(.A(KEYINPUT127), .B1(new_n1234), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g826(.A(KEYINPUT127), .ZN(new_n1252));
  AND3_X1   g827(.A1(new_n1119), .A2(new_n1230), .A3(new_n1131), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1052), .A2(KEYINPUT62), .ZN(new_n1254));
  NAND3_X1  g829(.A1(new_n1253), .A2(new_n1254), .A3(new_n1228), .ZN(new_n1255));
  INV_X1    g830(.A(new_n1211), .ZN(new_n1256));
  INV_X1    g831(.A(new_n1218), .ZN(new_n1257));
  INV_X1    g832(.A(new_n1224), .ZN(new_n1258));
  AOI21_X1  g833(.A(new_n1223), .B1(new_n1130), .B2(new_n1222), .ZN(new_n1259));
  OAI21_X1  g834(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g835(.A1(new_n1126), .A2(new_n1091), .A3(new_n1130), .ZN(new_n1261));
  INV_X1    g836(.A(new_n1215), .ZN(new_n1262));
  OAI21_X1  g837(.A(new_n1212), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g838(.A(new_n1256), .B1(new_n1260), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g839(.A1(new_n1255), .A2(new_n1264), .ZN(new_n1265));
  AOI22_X1  g840(.A1(new_n1195), .A2(new_n1199), .B1(new_n1202), .B2(new_n1166), .ZN(new_n1266));
  NAND2_X1  g841(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1267));
  AOI21_X1  g842(.A(new_n1266), .B1(new_n1267), .B2(KEYINPUT126), .ZN(new_n1268));
  AOI21_X1  g843(.A(new_n1265), .B1(new_n1268), .B2(new_n1152), .ZN(new_n1269));
  OAI211_X1 g844(.A(new_n1252), .B(new_n1249), .C1(new_n1269), .C2(new_n1027), .ZN(new_n1270));
  NAND2_X1  g845(.A1(new_n1251), .A2(new_n1270), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g846(.A(G319), .ZN(new_n1273));
  NOR4_X1   g847(.A1(G229), .A2(new_n1273), .A3(G401), .A4(G227), .ZN(new_n1274));
  OAI211_X1 g848(.A(new_n993), .B(new_n1274), .C1(new_n940), .C2(new_n941), .ZN(G225));
  INV_X1    g849(.A(G225), .ZN(G308));
endmodule


