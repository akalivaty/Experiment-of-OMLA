

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592;

  NOR2_X2 U327 ( .A1(n575), .A2(n468), .ZN(n543) );
  XOR2_X1 U328 ( .A(KEYINPUT36), .B(n568), .Z(n589) );
  NOR2_X1 U329 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U330 ( .A(n389), .B(n388), .ZN(n568) );
  XOR2_X1 U331 ( .A(KEYINPUT38), .B(n488), .Z(n496) );
  XNOR2_X1 U332 ( .A(n332), .B(n331), .ZN(n542) );
  XOR2_X1 U333 ( .A(n299), .B(KEYINPUT22), .Z(n295) );
  XOR2_X1 U334 ( .A(n326), .B(n371), .Z(n296) );
  XNOR2_X1 U335 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n297) );
  NOR2_X1 U336 ( .A1(n589), .A2(n484), .ZN(n485) );
  XNOR2_X1 U337 ( .A(n420), .B(n382), .ZN(n383) );
  NOR2_X1 U338 ( .A1(n542), .A2(n466), .ZN(n472) );
  XNOR2_X1 U339 ( .A(n384), .B(n383), .ZN(n386) );
  INV_X1 U340 ( .A(G183GAT), .ZN(n454) );
  XOR2_X1 U341 ( .A(n452), .B(KEYINPUT120), .Z(n567) );
  XNOR2_X1 U342 ( .A(n454), .B(KEYINPUT122), .ZN(n455) );
  XNOR2_X1 U343 ( .A(n456), .B(n455), .ZN(G1350GAT) );
  XNOR2_X1 U344 ( .A(n297), .B(KEYINPUT2), .ZN(n326) );
  XOR2_X1 U345 ( .A(G50GAT), .B(G162GAT), .Z(n371) );
  NAND2_X1 U346 ( .A1(G228GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n296), .B(n298), .ZN(n299) );
  XOR2_X1 U348 ( .A(G22GAT), .B(G155GAT), .Z(n395) );
  XNOR2_X1 U349 ( .A(n395), .B(KEYINPUT24), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n295), .B(n300), .ZN(n304) );
  XOR2_X1 U351 ( .A(G211GAT), .B(KEYINPUT84), .Z(n302) );
  XNOR2_X1 U352 ( .A(KEYINPUT23), .B(G204GAT), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U354 ( .A(n304), .B(n303), .Z(n310) );
  XOR2_X1 U355 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n306) );
  XNOR2_X1 U356 ( .A(G197GAT), .B(G218GAT), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n306), .B(n305), .ZN(n426) );
  XOR2_X1 U358 ( .A(G78GAT), .B(G148GAT), .Z(n308) );
  XNOR2_X1 U359 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n340) );
  XNOR2_X1 U361 ( .A(n426), .B(n340), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n467) );
  XOR2_X1 U363 ( .A(KEYINPUT78), .B(G127GAT), .Z(n312) );
  XNOR2_X1 U364 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U366 ( .A(G113GAT), .B(n313), .ZN(n449) );
  INV_X1 U367 ( .A(n449), .ZN(n332) );
  XOR2_X1 U368 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n315) );
  XNOR2_X1 U369 ( .A(KEYINPUT88), .B(KEYINPUT1), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U371 ( .A(KEYINPUT5), .B(G57GAT), .Z(n317) );
  XNOR2_X1 U372 ( .A(G1GAT), .B(G148GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n330) );
  XOR2_X1 U375 ( .A(G134GAT), .B(KEYINPUT73), .Z(n374) );
  XOR2_X1 U376 ( .A(G85GAT), .B(G162GAT), .Z(n321) );
  XNOR2_X1 U377 ( .A(G29GAT), .B(G155GAT), .ZN(n320) );
  XNOR2_X1 U378 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U379 ( .A(n374), .B(n322), .Z(n324) );
  NAND2_X1 U380 ( .A1(G225GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U382 ( .A(n325), .B(KEYINPUT86), .Z(n328) );
  XNOR2_X1 U383 ( .A(n326), .B(KEYINPUT87), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n331) );
  INV_X1 U386 ( .A(n542), .ZN(n574) );
  AND2_X1 U387 ( .A1(n467), .A2(n574), .ZN(n431) );
  XOR2_X1 U388 ( .A(KEYINPUT71), .B(KEYINPUT31), .Z(n334) );
  XNOR2_X1 U389 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n333) );
  XNOR2_X1 U390 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U391 ( .A(G99GAT), .B(G85GAT), .Z(n373) );
  XNOR2_X1 U392 ( .A(n335), .B(n373), .ZN(n337) );
  AND2_X1 U393 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n339) );
  INV_X1 U395 ( .A(KEYINPUT32), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n340), .B(KEYINPUT70), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n348) );
  XOR2_X1 U399 ( .A(KEYINPUT13), .B(KEYINPUT69), .Z(n344) );
  XNOR2_X1 U400 ( .A(G71GAT), .B(G57GAT), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n344), .B(n343), .ZN(n393) );
  XOR2_X1 U402 ( .A(G64GAT), .B(G92GAT), .Z(n346) );
  XNOR2_X1 U403 ( .A(G176GAT), .B(G204GAT), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n425) );
  XOR2_X1 U405 ( .A(n393), .B(n425), .Z(n347) );
  XOR2_X1 U406 ( .A(n348), .B(n347), .Z(n582) );
  XOR2_X1 U407 ( .A(KEYINPUT41), .B(n582), .Z(n550) );
  XOR2_X1 U408 ( .A(G8GAT), .B(G113GAT), .Z(n350) );
  XNOR2_X1 U409 ( .A(G169GAT), .B(G141GAT), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U411 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n352) );
  XNOR2_X1 U412 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n366) );
  XNOR2_X1 U415 ( .A(G22GAT), .B(G50GAT), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n355), .B(G36GAT), .ZN(n357) );
  XNOR2_X1 U417 ( .A(G15GAT), .B(G1GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n356), .B(KEYINPUT67), .ZN(n391) );
  XOR2_X1 U419 ( .A(n357), .B(n391), .Z(n364) );
  XOR2_X1 U420 ( .A(G29GAT), .B(G43GAT), .Z(n359) );
  XNOR2_X1 U421 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n387) );
  XOR2_X1 U423 ( .A(n387), .B(KEYINPUT66), .Z(n361) );
  NAND2_X1 U424 ( .A1(G229GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n362), .B(G197GAT), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n560) );
  INV_X1 U429 ( .A(n560), .ZN(n578) );
  NOR2_X1 U430 ( .A1(n550), .A2(n578), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n367), .B(KEYINPUT46), .ZN(n390) );
  XOR2_X1 U432 ( .A(KEYINPUT74), .B(KEYINPUT10), .Z(n369) );
  XNOR2_X1 U433 ( .A(G92GAT), .B(KEYINPUT64), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U435 ( .A(n371), .B(n370), .Z(n381) );
  INV_X1 U436 ( .A(n374), .ZN(n372) );
  NAND2_X1 U437 ( .A1(n373), .A2(n372), .ZN(n377) );
  INV_X1 U438 ( .A(n373), .ZN(n375) );
  NAND2_X1 U439 ( .A1(n375), .A2(n374), .ZN(n376) );
  NAND2_X1 U440 ( .A1(n377), .A2(n376), .ZN(n379) );
  NAND2_X1 U441 ( .A1(G232GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n384) );
  XOR2_X1 U444 ( .A(G36GAT), .B(G190GAT), .Z(n420) );
  XNOR2_X1 U445 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n382) );
  INV_X1 U446 ( .A(KEYINPUT9), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n385), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n387), .B(G106GAT), .ZN(n388) );
  NOR2_X1 U449 ( .A1(n390), .A2(n568), .ZN(n409) );
  INV_X1 U450 ( .A(n391), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n408) );
  XNOR2_X1 U452 ( .A(G8GAT), .B(G183GAT), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n394), .B(G211GAT), .ZN(n423) );
  XOR2_X1 U454 ( .A(n423), .B(n395), .Z(n397) );
  XNOR2_X1 U455 ( .A(G127GAT), .B(G78GAT), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U457 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n399) );
  NAND2_X1 U458 ( .A1(G231GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U460 ( .A(n401), .B(n400), .Z(n406) );
  XOR2_X1 U461 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n403) );
  XNOR2_X1 U462 ( .A(G64GAT), .B(KEYINPUT75), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n404), .B(KEYINPUT15), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U466 ( .A(n408), .B(n407), .Z(n585) );
  XOR2_X1 U467 ( .A(KEYINPUT107), .B(n585), .Z(n534) );
  NAND2_X1 U468 ( .A1(n409), .A2(n534), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n410), .B(KEYINPUT47), .ZN(n415) );
  NOR2_X1 U470 ( .A1(n589), .A2(n585), .ZN(n411) );
  XNOR2_X1 U471 ( .A(KEYINPUT45), .B(n411), .ZN(n413) );
  AND2_X1 U472 ( .A1(n582), .A2(n578), .ZN(n412) );
  AND2_X1 U473 ( .A1(n413), .A2(n412), .ZN(n414) );
  XNOR2_X1 U474 ( .A(KEYINPUT48), .B(n416), .ZN(n545) );
  XOR2_X1 U475 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n418) );
  XNOR2_X1 U476 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U478 ( .A(G169GAT), .B(n419), .Z(n446) );
  XOR2_X1 U479 ( .A(KEYINPUT89), .B(n420), .Z(n422) );
  NAND2_X1 U480 ( .A1(G226GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n424) );
  XOR2_X1 U482 ( .A(n424), .B(n423), .Z(n428) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n446), .B(n429), .ZN(n461) );
  NOR2_X1 U486 ( .A1(n545), .A2(n461), .ZN(n430) );
  XNOR2_X1 U487 ( .A(KEYINPUT54), .B(n430), .ZN(n573) );
  NAND2_X1 U488 ( .A1(n431), .A2(n573), .ZN(n433) );
  XOR2_X1 U489 ( .A(KEYINPUT119), .B(KEYINPUT55), .Z(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n451) );
  XOR2_X1 U491 ( .A(G176GAT), .B(KEYINPUT80), .Z(n435) );
  XNOR2_X1 U492 ( .A(KEYINPUT81), .B(KEYINPUT79), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U494 ( .A(G71GAT), .B(KEYINPUT20), .Z(n437) );
  XNOR2_X1 U495 ( .A(G183GAT), .B(KEYINPUT83), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U497 ( .A(n439), .B(n438), .Z(n448) );
  XOR2_X1 U498 ( .A(G190GAT), .B(G99GAT), .Z(n441) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(G134GAT), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U501 ( .A(G15GAT), .B(n442), .Z(n444) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n524) );
  NAND2_X1 U507 ( .A1(n451), .A2(n524), .ZN(n452) );
  INV_X1 U508 ( .A(n567), .ZN(n453) );
  NOR2_X1 U509 ( .A1(n453), .A2(n534), .ZN(n456) );
  XOR2_X1 U510 ( .A(KEYINPUT34), .B(KEYINPUT95), .Z(n476) );
  AND2_X1 U511 ( .A1(n560), .A2(n582), .ZN(n487) );
  INV_X1 U512 ( .A(n461), .ZN(n513) );
  NAND2_X1 U513 ( .A1(n513), .A2(n524), .ZN(n457) );
  NAND2_X1 U514 ( .A1(n457), .A2(n467), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n458), .B(KEYINPUT25), .ZN(n459) );
  XOR2_X1 U516 ( .A(KEYINPUT93), .B(n459), .Z(n464) );
  NOR2_X1 U517 ( .A1(n524), .A2(n467), .ZN(n460) );
  XOR2_X1 U518 ( .A(KEYINPUT26), .B(n460), .Z(n575) );
  XNOR2_X1 U519 ( .A(KEYINPUT27), .B(KEYINPUT90), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(n461), .ZN(n468) );
  XNOR2_X1 U521 ( .A(n543), .B(KEYINPUT92), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n465), .B(KEYINPUT94), .ZN(n466) );
  XOR2_X1 U524 ( .A(n467), .B(KEYINPUT28), .Z(n519) );
  NOR2_X1 U525 ( .A1(n519), .A2(n468), .ZN(n469) );
  NAND2_X1 U526 ( .A1(n469), .A2(n542), .ZN(n523) );
  NOR2_X1 U527 ( .A1(n524), .A2(n523), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT91), .B(n470), .Z(n471) );
  NOR2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n484) );
  NOR2_X1 U530 ( .A1(n568), .A2(n585), .ZN(n473) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  NOR2_X1 U532 ( .A1(n484), .A2(n474), .ZN(n498) );
  AND2_X1 U533 ( .A1(n487), .A2(n498), .ZN(n482) );
  NAND2_X1 U534 ( .A1(n482), .A2(n542), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n482), .A2(n513), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(KEYINPUT96), .ZN(n479) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(n479), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .Z(n481) );
  NAND2_X1 U541 ( .A1(n482), .A2(n524), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NAND2_X1 U543 ( .A1(n482), .A2(n519), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U545 ( .A1(n485), .A2(n585), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT37), .B(n486), .ZN(n508) );
  NAND2_X1 U547 ( .A1(n487), .A2(n508), .ZN(n488) );
  NAND2_X1 U548 ( .A1(n496), .A2(n542), .ZN(n491) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(KEYINPUT97), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n496), .A2(n513), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT98), .B(KEYINPUT40), .Z(n494) );
  NAND2_X1 U555 ( .A1(n524), .A2(n496), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U557 ( .A(G43GAT), .B(n495), .Z(G1330GAT) );
  NAND2_X1 U558 ( .A1(n496), .A2(n519), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U560 ( .A(n550), .B(KEYINPUT99), .ZN(n562) );
  AND2_X1 U561 ( .A1(n578), .A2(n562), .ZN(n509) );
  AND2_X1 U562 ( .A1(n509), .A2(n498), .ZN(n505) );
  NAND2_X1 U563 ( .A1(n505), .A2(n542), .ZN(n499) );
  XNOR2_X1 U564 ( .A(KEYINPUT42), .B(n499), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n500), .ZN(G1332GAT) );
  NAND2_X1 U566 ( .A1(n505), .A2(n513), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n501), .B(KEYINPUT100), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  XOR2_X1 U569 ( .A(G71GAT), .B(KEYINPUT101), .Z(n504) );
  NAND2_X1 U570 ( .A1(n505), .A2(n524), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .Z(n507) );
  NAND2_X1 U573 ( .A1(n505), .A2(n519), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  XOR2_X1 U575 ( .A(G85GAT), .B(KEYINPUT103), .Z(n512) );
  NAND2_X1 U576 ( .A1(n509), .A2(n508), .ZN(n510) );
  XOR2_X1 U577 ( .A(KEYINPUT102), .B(n510), .Z(n518) );
  NAND2_X1 U578 ( .A1(n518), .A2(n542), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n518), .A2(n513), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(KEYINPUT104), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(n515), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT105), .Z(n517) );
  NAND2_X1 U584 ( .A1(n524), .A2(n518), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT106), .Z(n521) );
  NAND2_X1 U587 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U589 ( .A(G106GAT), .B(n522), .Z(G1339GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n528) );
  NOR2_X1 U591 ( .A1(n545), .A2(n523), .ZN(n525) );
  NAND2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U593 ( .A(KEYINPUT108), .B(n526), .Z(n537) );
  NAND2_X1 U594 ( .A1(n560), .A2(n537), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U598 ( .A1(n537), .A2(n562), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U600 ( .A(G120GAT), .B(n532), .Z(G1341GAT) );
  INV_X1 U601 ( .A(n537), .ZN(n533) );
  NOR2_X1 U602 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(n535), .Z(n536) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U606 ( .A1(n568), .A2(n537), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT112), .Z(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n558), .A2(n560), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT114), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n549) );
  XNOR2_X1 U616 ( .A(KEYINPUT115), .B(KEYINPUT53), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n554) );
  INV_X1 U618 ( .A(n558), .ZN(n555) );
  NOR2_X1 U619 ( .A1(n550), .A2(n555), .ZN(n552) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U622 ( .A(n554), .B(n553), .Z(G1345GAT) );
  OR2_X1 U623 ( .A1(n585), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT118), .ZN(n557) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n558), .A2(n568), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n567), .A2(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT57), .Z(n564) );
  NAND2_X1 U631 ( .A1(n562), .A2(n567), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n566) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n572) );
  XOR2_X1 U636 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n570) );
  NAND2_X1 U637 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U638 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(G1351GAT) );
  AND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n577) );
  INV_X1 U641 ( .A(n575), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n588) );
  NOR2_X1 U643 ( .A1(n578), .A2(n588), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n588), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n588), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(G218GAT), .B(n592), .Z(G1355GAT) );
endmodule

