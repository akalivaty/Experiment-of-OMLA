//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n192), .A2(KEYINPUT87), .A3(KEYINPUT88), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT88), .B1(new_n192), .B2(KEYINPUT87), .ZN(new_n194));
  XNOR2_X1  g008(.A(G125), .B(G140), .ZN(new_n195));
  OAI22_X1  g009(.A1(new_n193), .A2(new_n194), .B1(new_n191), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(KEYINPUT87), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT88), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n195), .A2(new_n191), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n192), .A2(KEYINPUT87), .A3(KEYINPUT88), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(G237), .A2(G953), .ZN(new_n203));
  AOI21_X1  g017(.A(G143), .B1(new_n203), .B2(G214), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(G143), .A3(G214), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n205), .A2(KEYINPUT18), .A3(G131), .A4(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT18), .A2(G131), .ZN(new_n208));
  INV_X1    g022(.A(new_n206), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(new_n204), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n196), .A2(new_n202), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT89), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT89), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n196), .A2(new_n202), .A3(new_n214), .A4(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n195), .A2(KEYINPUT16), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n188), .A2(KEYINPUT16), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(G146), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(G146), .B1(new_n217), .B2(new_n218), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(KEYINPUT17), .B(G131), .C1(new_n209), .C2(new_n204), .ZN(new_n223));
  OAI21_X1  g037(.A(G131), .B1(new_n209), .B2(new_n204), .ZN(new_n224));
  INV_X1    g038(.A(G131), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n205), .A2(new_n225), .A3(new_n206), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n222), .B(new_n223), .C1(KEYINPUT17), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n216), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G113), .B(G122), .ZN(new_n230));
  INV_X1    g044(.A(G104), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT93), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(G902), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n229), .A2(new_n234), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G475), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT90), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT90), .B1(new_n224), .B2(new_n226), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT19), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n188), .B(new_n190), .C1(KEYINPUT91), .C2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n243), .B(new_n191), .C1(new_n195), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n219), .ZN(new_n246));
  NOR3_X1   g060(.A1(new_n240), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n216), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT92), .A3(new_n233), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n247), .B1(new_n213), .B2(new_n215), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(new_n232), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n216), .A2(new_n232), .A3(new_n228), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT20), .ZN(new_n256));
  NOR2_X1   g070(.A1(G475), .A2(G902), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n256), .B1(new_n255), .B2(new_n257), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n239), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(G234), .A2(G237), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(G952), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(G902), .A3(G953), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT21), .B(G898), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G902), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT9), .B(G234), .ZN(new_n273));
  INV_X1    g087(.A(G217), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n273), .A2(new_n274), .A3(G953), .ZN(new_n275));
  XOR2_X1   g089(.A(G116), .B(G122), .Z(new_n276));
  OR2_X1    g090(.A1(new_n276), .A2(G107), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(G107), .ZN(new_n278));
  INV_X1    g092(.A(G134), .ZN(new_n279));
  XNOR2_X1  g093(.A(G128), .B(G143), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n277), .A2(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G143), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT13), .B1(new_n282), .B2(G128), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(G128), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(KEYINPUT94), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT13), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT95), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G128), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(G143), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT95), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT13), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(new_n287), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT94), .B1(new_n283), .B2(new_n284), .ZN(new_n293));
  OAI211_X1 g107(.A(KEYINPUT96), .B(G134), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT94), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n286), .B1(new_n288), .B2(G143), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n296), .B1(new_n297), .B2(new_n289), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n298), .A2(new_n285), .A3(new_n287), .A4(new_n291), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT96), .B1(new_n299), .B2(G134), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n281), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT97), .ZN(new_n302));
  OAI21_X1  g116(.A(G134), .B1(new_n292), .B2(new_n293), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT96), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n294), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT97), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(new_n281), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n280), .B(new_n279), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT14), .A3(G122), .ZN(new_n312));
  OAI211_X1 g126(.A(G107), .B(new_n312), .C1(new_n276), .C2(KEYINPUT14), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n277), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n275), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n314), .ZN(new_n316));
  INV_X1    g130(.A(new_n275), .ZN(new_n317));
  AOI211_X1 g131(.A(new_n316), .B(new_n317), .C1(new_n302), .C2(new_n308), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n272), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT98), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G478), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(KEYINPUT15), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT98), .B(new_n272), .C1(new_n315), .C2(new_n318), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n301), .A2(KEYINPUT97), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n307), .B1(new_n306), .B2(new_n281), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n314), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n317), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n309), .A2(new_n314), .A3(new_n275), .ZN(new_n330));
  AOI21_X1  g144(.A(G902), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n323), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT99), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n325), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n321), .A2(KEYINPUT99), .A3(new_n323), .A4(new_n324), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT100), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(KEYINPUT100), .A3(new_n335), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n271), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT11), .B1(new_n279), .B2(G137), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT11), .ZN(new_n342));
  INV_X1    g156(.A(G137), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(G134), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT65), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n343), .B2(G134), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n279), .A2(KEYINPUT65), .A3(G137), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G131), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT66), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n341), .A2(new_n344), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n352), .A2(new_n225), .A3(new_n347), .A4(new_n348), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(KEYINPUT0), .A2(G128), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n355), .A2(KEYINPUT64), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT0), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(new_n288), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n191), .A2(G143), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n282), .A2(G146), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n355), .A2(KEYINPUT64), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n356), .A2(new_n359), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT66), .B(G131), .C1(new_n345), .C2(new_n349), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n354), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G119), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G116), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n311), .A2(G119), .ZN(new_n371));
  INV_X1    g185(.A(G113), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n372), .A2(KEYINPUT2), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(KEYINPUT2), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n370), .B(new_n371), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n370), .A2(new_n371), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT2), .B(G113), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT1), .B1(new_n282), .B2(G146), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n362), .A2(G128), .A3(new_n381), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n360), .B(new_n361), .C1(KEYINPUT1), .C2(new_n288), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n279), .A2(G137), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n343), .A2(G134), .ZN(new_n386));
  OAI21_X1  g200(.A(G131), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n353), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n368), .A2(new_n380), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT67), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT67), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n368), .A2(new_n391), .A3(new_n380), .A4(new_n388), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n368), .A2(new_n388), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n379), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT28), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT28), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n400));
  NAND2_X1  g214(.A1(new_n203), .A2(G210), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT26), .B(G101), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(G902), .B1(new_n406), .B2(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n390), .A2(new_n392), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT30), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n368), .A2(new_n410), .A3(new_n388), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n368), .B2(new_n388), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n379), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT29), .B1(new_n414), .B2(new_n405), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT70), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n415), .B1(new_n406), .B2(new_n416), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n399), .A2(KEYINPUT70), .A3(new_n405), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n407), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G472), .ZN(new_n420));
  INV_X1    g234(.A(G472), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n413), .A2(new_n390), .A3(new_n392), .A4(new_n404), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n399), .A2(new_n405), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT31), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT69), .B1(new_n422), .B2(KEYINPUT31), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n393), .A2(KEYINPUT30), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n368), .A2(new_n410), .A3(new_n388), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n380), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(new_n408), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT69), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(new_n432), .A3(new_n425), .A4(new_n404), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n421), .B(new_n272), .C1(new_n426), .C2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(KEYINPUT32), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT32), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n427), .A2(new_n433), .ZN(new_n438));
  INV_X1    g252(.A(new_n398), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n395), .B2(KEYINPUT28), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n425), .B1(new_n440), .B2(new_n404), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n422), .ZN(new_n442));
  AOI21_X1  g256(.A(G902), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n437), .B1(new_n443), .B2(new_n421), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n420), .B1(new_n436), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n274), .B1(G234), .B2(new_n272), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT24), .B(G110), .Z(new_n447));
  NOR2_X1   g261(.A1(new_n369), .A2(G128), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n288), .A2(G119), .ZN(new_n449));
  OR3_X1    g263(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT71), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT71), .B1(new_n448), .B2(new_n449), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT72), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n448), .B1(new_n453), .B2(KEYINPUT23), .ZN(new_n454));
  INV_X1    g268(.A(G110), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT23), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT72), .B1(new_n369), .B2(G128), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n454), .B(new_n455), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n219), .B(new_n192), .C1(new_n452), .C2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G110), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n450), .A2(new_n451), .A3(new_n447), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n463), .B(new_n464), .C1(new_n220), .C2(new_n221), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT22), .B(G137), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n461), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n461), .B2(new_n465), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT25), .B1(new_n471), .B2(new_n272), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT25), .ZN(new_n473));
  NOR4_X1   g287(.A1(new_n469), .A2(new_n470), .A3(new_n473), .A4(G902), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n446), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n446), .A2(G902), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT73), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G214), .B1(G237), .B2(G902), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT80), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n370), .B2(KEYINPUT5), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT5), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT5), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n486), .A2(new_n369), .A3(KEYINPUT80), .A4(G116), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n484), .A2(new_n485), .A3(G113), .A4(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT3), .B1(new_n231), .B2(G107), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT3), .ZN(new_n490));
  INV_X1    g304(.A(G107), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(G104), .ZN(new_n492));
  INV_X1    g306(.A(G101), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n231), .A2(G107), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n489), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n231), .A2(G107), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n491), .A2(G104), .ZN(new_n497));
  OAI21_X1  g311(.A(G101), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n488), .A2(new_n375), .A3(new_n495), .A4(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT81), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n495), .A2(new_n498), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n502), .A2(KEYINPUT81), .A3(new_n375), .A4(new_n488), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n489), .A2(new_n492), .A3(new_n494), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G101), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n507), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT4), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n509), .A3(G101), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n379), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT79), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n507), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT79), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n379), .A4(new_n510), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n505), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(G110), .B(G122), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n505), .A2(new_n516), .A3(new_n518), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n364), .A2(new_n365), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G125), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n382), .A2(new_n383), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT82), .B1(new_n525), .B2(new_n189), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT82), .ZN(new_n527));
  AOI211_X1 g341(.A(new_n527), .B(G125), .C1(new_n382), .C2(new_n383), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n263), .A2(G224), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n529), .B(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT6), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n517), .A2(new_n533), .A3(new_n519), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n522), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n488), .A2(new_n375), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n495), .A2(new_n498), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT83), .A3(new_n499), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n518), .B(KEYINPUT8), .Z(new_n540));
  AOI22_X1  g354(.A1(new_n488), .A2(new_n375), .B1(new_n495), .B2(new_n498), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT83), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT84), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n539), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n529), .A2(new_n546), .A3(new_n531), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n544), .B1(new_n539), .B2(new_n543), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n504), .B1(new_n515), .B2(new_n512), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n527), .B1(new_n384), .B2(G125), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n525), .A2(KEYINPUT82), .A3(new_n189), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(KEYINPUT85), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT85), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n526), .B2(new_n528), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n555), .A3(new_n524), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT86), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n531), .B1(new_n557), .B2(new_n546), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n557), .B2(new_n546), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n550), .A2(new_n518), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(G902), .B1(new_n549), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n535), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(G210), .B1(G237), .B2(G902), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n535), .A2(new_n561), .A3(new_n563), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n482), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G469), .ZN(new_n569));
  XNOR2_X1  g383(.A(G110), .B(G140), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT75), .ZN(new_n571));
  INV_X1    g385(.A(G227), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(G953), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n571), .B(new_n573), .Z(new_n574));
  AND2_X1   g388(.A1(new_n354), .A2(new_n367), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n384), .A2(KEYINPUT76), .A3(new_n502), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT76), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n525), .B2(new_n537), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n366), .A2(new_n513), .A3(new_n510), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n525), .A2(new_n537), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT10), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n575), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT78), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n354), .A2(new_n367), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n510), .A2(new_n364), .A3(new_n365), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n588), .A2(new_n513), .B1(new_n582), .B2(KEYINPUT10), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT78), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n589), .A2(new_n590), .A3(new_n587), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n574), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n525), .A2(new_n537), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n576), .A2(new_n579), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n598), .A2(new_n575), .A3(KEYINPUT12), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT12), .B1(new_n598), .B2(new_n575), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n595), .A2(new_n574), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n569), .B(new_n272), .C1(new_n596), .C2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n569), .A2(new_n272), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT77), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n595), .A2(KEYINPUT77), .A3(new_n574), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n594), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n595), .B1(new_n599), .B2(new_n600), .ZN(new_n611));
  INV_X1    g425(.A(new_n574), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n613), .A3(G469), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n604), .A2(new_n606), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(G221), .B1(new_n273), .B2(G902), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT74), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n568), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n340), .A2(new_n445), .A3(new_n480), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  NAND3_X1  g436(.A1(new_n442), .A2(new_n427), .A3(new_n433), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n272), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(G472), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n435), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n615), .A2(new_n618), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n480), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n322), .A2(G902), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n635), .B(new_n636), .C1(new_n315), .C2(new_n318), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n329), .A2(new_n633), .A3(new_n634), .A4(new_n330), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n632), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n260), .B1(new_n630), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n535), .A2(new_n561), .A3(new_n563), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n563), .B1(new_n535), .B2(new_n561), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n481), .B(new_n270), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n629), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G104), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT102), .B(KEYINPUT34), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  AND3_X1   g462(.A1(new_n334), .A2(KEYINPUT100), .A3(new_n335), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT100), .B1(new_n334), .B2(new_n335), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n649), .A2(new_n650), .A3(new_n260), .ZN(new_n651));
  INV_X1    g465(.A(new_n643), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n629), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n443), .A2(new_n421), .ZN(new_n656));
  INV_X1    g470(.A(new_n435), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n461), .A2(new_n465), .ZN(new_n658));
  INV_X1    g472(.A(new_n468), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n658), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n478), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n475), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n656), .A2(new_n657), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n340), .A2(new_n620), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n265), .B1(new_n267), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n568), .A2(new_n619), .A3(new_n664), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n651), .A2(new_n445), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  NOR2_X1   g488(.A1(new_n649), .A2(new_n650), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n670), .B(KEYINPUT39), .Z(new_n676));
  NAND2_X1  g490(.A1(new_n627), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n675), .B(new_n260), .C1(KEYINPUT40), .C2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n565), .A2(new_n566), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT38), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n679), .A2(new_n481), .A3(new_n664), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n414), .A2(new_n404), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n395), .A2(new_n404), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(G902), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n421), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n435), .A2(KEYINPUT32), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n443), .A2(new_n437), .A3(new_n421), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OR3_X1    g503(.A1(new_n678), .A2(new_n682), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  NAND2_X1  g505(.A1(new_n637), .A2(new_n638), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n631), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n695), .A2(new_n260), .A3(new_n671), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n445), .A2(new_n672), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  NOR2_X1   g512(.A1(new_n591), .A2(new_n592), .ZN(new_n699));
  AOI211_X1 g513(.A(KEYINPUT78), .B(new_n587), .C1(new_n589), .C2(new_n590), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n595), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n603), .B1(new_n701), .B2(new_n612), .ZN(new_n702));
  OAI21_X1  g516(.A(G469), .B1(new_n702), .B2(G902), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n703), .A2(new_n618), .A3(new_n604), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n445), .A2(new_n480), .A3(new_n644), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  INV_X1    g521(.A(new_n480), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n687), .A2(new_n688), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n708), .B1(new_n709), .B2(new_n420), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n704), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n651), .A2(new_n652), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NAND3_X1  g528(.A1(new_n704), .A2(new_n567), .A3(new_n663), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n340), .A2(new_n445), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  NOR4_X1   g532(.A1(new_n649), .A2(new_n650), .A3(new_n568), .A4(new_n261), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n703), .A2(new_n604), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n720), .A2(new_n617), .A3(new_n269), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n435), .A2(KEYINPUT103), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n623), .A2(new_n723), .A3(new_n421), .A4(new_n272), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n625), .A2(new_n722), .A3(new_n480), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT104), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n725), .A2(KEYINPUT104), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n719), .B(new_n721), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  NAND3_X1  g544(.A1(new_n695), .A2(new_n260), .A3(new_n671), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n715), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n625), .A3(new_n724), .A4(new_n722), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n611), .A2(new_n735), .A3(new_n612), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n735), .B1(new_n611), .B2(new_n612), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n610), .B(G469), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n604), .A2(new_n606), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n617), .A2(new_n482), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n565), .A2(new_n566), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT106), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n740), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n641), .A2(new_n642), .A3(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n604), .A2(new_n606), .A3(new_n738), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n731), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n445), .A2(new_n748), .A3(new_n480), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n710), .A2(KEYINPUT42), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND4_X1  g568(.A1(new_n338), .A2(new_n339), .A3(new_n261), .A4(new_n671), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n739), .A2(new_n741), .A3(KEYINPUT106), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n710), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  AOI21_X1  g575(.A(KEYINPUT45), .B1(new_n610), .B2(new_n613), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n569), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n610), .B(KEYINPUT45), .C1(new_n736), .C2(new_n737), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n606), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n604), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n766), .A2(new_n767), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n618), .B(new_n676), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT107), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n261), .A2(new_n695), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT43), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n626), .A2(new_n663), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  OR3_X1    g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n776), .B1(new_n774), .B2(new_n775), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n565), .A2(new_n481), .A3(new_n566), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n772), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n343), .ZN(G39));
  OAI21_X1  g597(.A(new_n618), .B1(new_n769), .B2(new_n770), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT47), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(KEYINPUT47), .B(new_n618), .C1(new_n769), .C2(new_n770), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n445), .A2(new_n480), .A3(new_n731), .A4(new_n779), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  XNOR2_X1  g605(.A(new_n720), .B(KEYINPUT108), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT49), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(KEYINPUT49), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n681), .A2(new_n773), .A3(new_n708), .A4(new_n743), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n794), .A2(new_n795), .A3(new_n689), .A4(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n798));
  NOR2_X1   g612(.A1(new_n774), .A2(new_n264), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n741), .A2(new_n720), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT115), .ZN(new_n802));
  INV_X1    g616(.A(new_n710), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n798), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n480), .A2(new_n689), .A3(new_n265), .A4(new_n800), .ZN(new_n805));
  INV_X1    g619(.A(new_n640), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n804), .A2(G952), .A3(new_n263), .A4(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n725), .A2(KEYINPUT104), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n726), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n799), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n811), .A2(new_n568), .A3(new_n617), .A4(new_n720), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n802), .A2(new_n803), .A3(new_n798), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n808), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n625), .A2(new_n722), .A3(new_n663), .A4(new_n724), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n802), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n805), .A2(new_n261), .A3(new_n694), .A4(new_n693), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT51), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n811), .A2(new_n779), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n792), .A2(new_n617), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n786), .A2(new_n787), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n811), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n681), .A2(new_n481), .A3(new_n617), .A4(new_n720), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT50), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n823), .A2(KEYINPUT50), .A3(new_n824), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n816), .B(new_n822), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n816), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n788), .A2(KEYINPUT114), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n820), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n788), .A2(KEYINPUT114), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n819), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n817), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n814), .B(new_n827), .C1(KEYINPUT51), .C2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT110), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n663), .A2(new_n617), .A3(new_n670), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n746), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n746), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n689), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n836), .B1(new_n842), .B2(new_n719), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n338), .A2(new_n567), .A3(new_n339), .A4(new_n260), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n844), .A2(new_n689), .A3(new_n841), .A4(KEYINPUT111), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n445), .A2(new_n672), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n697), .B(new_n733), .C1(new_n847), .C2(new_n755), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT52), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n705), .B(new_n717), .C1(new_n711), .C2(new_n712), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n675), .A2(new_n567), .A3(new_n260), .A4(new_n721), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n809), .B2(new_n726), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT109), .B1(new_n640), .B2(new_n643), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT109), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n652), .A2(new_n854), .A3(new_n260), .A4(new_n695), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n652), .A2(new_n261), .A3(new_n334), .A4(new_n335), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n629), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n621), .A2(new_n858), .A3(new_n666), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n850), .A2(new_n852), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n848), .ZN(new_n861));
  INV_X1    g675(.A(new_n686), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(new_n436), .B2(new_n444), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n839), .A2(new_n840), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT111), .B1(new_n865), .B2(new_n844), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n842), .A2(new_n719), .A3(new_n836), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n861), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n696), .B1(new_n756), .B2(new_n757), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n687), .A2(new_n688), .B1(G472), .B2(new_n419), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n670), .B1(new_n475), .B2(new_n662), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n239), .B(new_n873), .C1(new_n258), .C2(new_n259), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n779), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n627), .A2(new_n875), .A3(new_n336), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n871), .A2(new_n815), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  AOI221_X4 g691(.A(new_n877), .B1(new_n759), .B2(new_n710), .C1(new_n751), .C2(new_n752), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n849), .A2(new_n860), .A3(new_n870), .A4(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n877), .ZN(new_n882));
  INV_X1    g696(.A(new_n752), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT42), .B1(new_n710), .B2(new_n748), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n760), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n848), .B1(new_n866), .B2(new_n867), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n886), .B2(new_n869), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n869), .B1(new_n673), .B2(new_n733), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n888), .A2(KEYINPUT53), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n887), .A2(new_n860), .A3(new_n849), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n849), .A2(new_n870), .A3(new_n878), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n705), .A2(new_n717), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n713), .A2(new_n729), .A3(new_n894), .A4(KEYINPUT112), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n888), .A2(new_n859), .A3(new_n880), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT112), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n850), .B2(new_n852), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  XOR2_X1   g714(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n881), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n835), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(G952), .A2(G953), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n797), .B1(new_n904), .B2(new_n905), .ZN(G75));
  NOR2_X1   g720(.A1(new_n263), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI22_X1  g722(.A1(new_n893), .A2(new_n899), .B1(new_n879), .B2(new_n880), .ZN(new_n909));
  INV_X1    g723(.A(G210), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n272), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n522), .A2(new_n534), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT117), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n532), .B(KEYINPUT55), .Z(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n915), .A2(KEYINPUT56), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n908), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n900), .A2(new_n881), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(G902), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n920), .B2(new_n910), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n911), .A2(KEYINPUT118), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n917), .B1(new_n924), .B2(new_n915), .ZN(G51));
  XNOR2_X1  g739(.A(new_n605), .B(KEYINPUT57), .ZN(new_n926));
  INV_X1    g740(.A(new_n902), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n909), .A2(new_n901), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n702), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n909), .A2(new_n272), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n764), .A3(new_n763), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n907), .B1(new_n931), .B2(new_n933), .ZN(G54));
  INV_X1    g748(.A(new_n255), .ZN(new_n935));
  NAND2_X1  g749(.A1(KEYINPUT58), .A2(G475), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n920), .B2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .A4(new_n255), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n908), .ZN(G60));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT59), .Z(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n892), .B2(new_n902), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n908), .B1(new_n942), .B2(new_n692), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n637), .B2(new_n638), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n927), .B2(new_n928), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT119), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT119), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n947), .B(new_n944), .C1(new_n927), .C2(new_n928), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n943), .B1(new_n946), .B2(new_n948), .ZN(G63));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT60), .ZN(new_n951));
  OAI22_X1  g765(.A1(new_n909), .A2(new_n951), .B1(new_n469), .B2(new_n470), .ZN(new_n952));
  INV_X1    g766(.A(new_n951), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n879), .A2(new_n880), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n849), .A2(new_n870), .A3(new_n878), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n661), .B(new_n953), .C1(new_n954), .C2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n952), .A2(new_n958), .A3(new_n908), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n958), .A2(KEYINPUT120), .A3(new_n908), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT61), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n951), .B1(new_n900), .B2(new_n881), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n907), .B1(new_n962), .B2(new_n661), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n963), .B(new_n952), .C1(KEYINPUT120), .C2(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n961), .A2(new_n965), .ZN(G66));
  INV_X1    g780(.A(new_n268), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n263), .B1(new_n967), .B2(G224), .ZN(new_n968));
  INV_X1    g782(.A(new_n860), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n969), .B2(new_n263), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n913), .B1(G898), .B2(new_n263), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(new_n971), .Z(G69));
  NOR2_X1   g786(.A1(new_n411), .A2(new_n412), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n195), .A2(new_n244), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(new_n243), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n973), .B(new_n975), .Z(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT122), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n848), .B(KEYINPUT121), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n690), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n978), .B1(new_n980), .B2(KEYINPUT62), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT123), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n640), .B1(new_n336), .B2(new_n260), .ZN(new_n983));
  AOI211_X1 g797(.A(new_n779), .B(new_n677), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n984), .B(new_n710), .C1(new_n982), .C2(new_n983), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n790), .B(new_n985), .C1(new_n772), .C2(new_n781), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n980), .B2(KEYINPUT62), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT62), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n979), .A2(KEYINPUT122), .A3(new_n988), .A4(new_n690), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n981), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n977), .B1(new_n990), .B2(G953), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n977), .B1(G900), .B2(G953), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n782), .B1(new_n788), .B2(new_n789), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n719), .A2(new_n710), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n753), .B(new_n760), .C1(new_n772), .C2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n993), .A2(new_n979), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n992), .B1(new_n997), .B2(G953), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n572), .B2(new_n669), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT124), .Z(new_n1000));
  AND3_X1   g814(.A1(new_n991), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1000), .B1(new_n991), .B2(new_n998), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1001), .A2(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(new_n990), .A2(new_n860), .ZN(new_n1004));
  XNOR2_X1  g818(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT126), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n683), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1008), .B1(new_n997), .B2(new_n969), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n414), .A2(new_n404), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n908), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1011), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1014), .A2(new_n683), .A3(new_n1007), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT127), .Z(new_n1016));
  AOI21_X1  g830(.A(new_n1016), .B1(new_n881), .B2(new_n890), .ZN(new_n1017));
  NOR3_X1   g831(.A1(new_n1009), .A2(new_n1013), .A3(new_n1017), .ZN(G57));
endmodule


