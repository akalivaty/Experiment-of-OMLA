//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1293, new_n1294, new_n1295, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  OR2_X1    g0012(.A1(KEYINPUT65), .A2(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(KEYINPUT65), .A2(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n212), .B1(new_n218), .B2(new_n219), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n216), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT65), .A2(G20), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT65), .A2(G20), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT8), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT8), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G150), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(new_n201), .B2(new_n206), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n248), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(KEYINPUT69), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(KEYINPUT69), .ZN(new_n265));
  INV_X1    g0065(.A(G13), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n266), .A2(new_n206), .A3(G1), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n248), .ZN(new_n268));
  INV_X1    g0068(.A(G50), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n205), .B2(G20), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n268), .A2(new_n270), .B1(new_n269), .B2(new_n267), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n264), .A2(new_n265), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT68), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT68), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n275), .B(new_n205), .C1(G41), .C2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n279), .A2(G274), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n279), .A2(new_n273), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(G226), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(G222), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n286), .B1(new_n202), .B2(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n216), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n283), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n272), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT72), .B(G200), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n303), .B2(new_n293), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n272), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n272), .A2(new_n305), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n299), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n284), .A2(G232), .A3(G1698), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n284), .A2(G226), .A3(new_n285), .ZN(new_n313));
  AND3_X1   g0113(.A1(KEYINPUT74), .A2(G33), .A3(G97), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT74), .B1(G33), .B2(G97), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n291), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n280), .A2(new_n277), .B1(new_n282), .B2(G238), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n320), .B1(new_n319), .B2(new_n321), .ZN(new_n323));
  OAI21_X1  g0123(.A(G200), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT13), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(G190), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n267), .ZN(new_n329));
  OR3_X1    g0129(.A1(new_n329), .A2(KEYINPUT12), .A3(G68), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT12), .B1(new_n329), .B2(G68), .ZN(new_n331));
  INV_X1    g0131(.A(G68), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n205), .B2(G20), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n330), .A2(new_n331), .B1(new_n268), .B2(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n252), .B2(new_n202), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n248), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT11), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(KEYINPUT11), .A3(new_n248), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n334), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n324), .A2(new_n328), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n324), .A2(new_n328), .A3(new_n342), .A4(KEYINPUT75), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n248), .ZN(new_n348));
  AOI22_X1  g0148(.A1(G77), .A2(new_n215), .B1(new_n257), .B2(new_n260), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT70), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(G33), .A3(new_n251), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT71), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n348), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n205), .A2(G20), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n268), .A2(G77), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(G77), .B2(new_n329), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n281), .B1(G244), .B2(new_n282), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n284), .A2(G232), .A3(new_n285), .ZN(new_n361));
  INV_X1    g0161(.A(G107), .ZN(new_n362));
  INV_X1    g0162(.A(G238), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n361), .B1(new_n362), .B2(new_n284), .C1(new_n287), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n291), .ZN(new_n365));
  AOI21_X1  g0165(.A(G169), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT73), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n360), .A2(new_n365), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n366), .A2(new_n367), .B1(new_n368), .B2(G179), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n360), .A2(new_n365), .A3(KEYINPUT73), .A4(new_n296), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n359), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n355), .A2(new_n358), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n303), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n372), .B(new_n373), .C1(new_n300), .C2(new_n368), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n347), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n268), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n257), .A2(new_n356), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n376), .A2(new_n377), .B1(new_n329), .B2(new_n257), .ZN(new_n378));
  INV_X1    g0178(.A(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT3), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT3), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G33), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(new_n251), .A3(KEYINPUT7), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n284), .A2(G20), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(KEYINPUT77), .C1(new_n385), .C2(KEYINPUT7), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT77), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n383), .A2(new_n251), .A3(new_n387), .A4(KEYINPUT7), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(G68), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g0189(.A(G58), .B(G68), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n390), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n383), .A2(new_n251), .A3(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n396), .B(G68), .C1(new_n385), .C2(new_n395), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n397), .A2(new_n391), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n348), .B1(new_n398), .B2(KEYINPUT16), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n378), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n380), .A2(new_n382), .A3(G226), .A4(G1698), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n380), .A2(new_n382), .A3(G223), .A4(new_n285), .ZN(new_n402));
  INV_X1    g0202(.A(G87), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n401), .B(new_n402), .C1(new_n379), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n291), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n280), .A2(new_n277), .B1(new_n282), .B2(G232), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n405), .A2(new_n406), .A3(G179), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n294), .B1(new_n405), .B2(new_n406), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT78), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G169), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n405), .A2(new_n406), .A3(G179), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT18), .B1(new_n400), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n378), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT16), .B1(new_n389), .B2(new_n391), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n397), .A2(new_n391), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n248), .B1(new_n419), .B2(new_n393), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n417), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n409), .A4(new_n414), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G200), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n405), .B2(new_n406), .ZN(new_n426));
  XOR2_X1   g0226(.A(KEYINPUT79), .B(G190), .Z(new_n427));
  AND2_X1   g0227(.A1(new_n405), .A2(new_n406), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n417), .C1(new_n418), .C2(new_n420), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n400), .A2(KEYINPUT17), .A3(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n424), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n322), .A2(new_n323), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT14), .B1(new_n436), .B2(new_n294), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT14), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n438), .B(G169), .C1(new_n322), .C2(new_n323), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT76), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n436), .B2(G179), .ZN(new_n441));
  NOR4_X1   g0241(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT76), .A4(new_n296), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n437), .B(new_n439), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n341), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n311), .A2(new_n375), .A3(new_n435), .A4(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT87), .B(KEYINPUT22), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n213), .A2(new_n380), .A3(new_n382), .A4(new_n214), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n447), .B2(new_n403), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT22), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(KEYINPUT87), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n251), .A2(new_n284), .A3(G87), .A4(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT23), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n215), .A2(new_n452), .A3(new_n362), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G116), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G20), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(KEYINPUT88), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT88), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT23), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n362), .A2(G20), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n448), .A2(new_n451), .A3(new_n453), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT24), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n461), .A2(new_n453), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(new_n451), .A4(new_n448), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n248), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n266), .A2(G1), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(G20), .A3(new_n362), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n470), .B(KEYINPUT25), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n205), .A2(G33), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n268), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(G107), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n380), .A2(new_n382), .A3(G257), .A4(G1698), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n380), .A2(new_n382), .A3(G250), .A4(new_n285), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G294), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n291), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n481), .A2(G274), .A3(new_n279), .A4(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n481), .A2(new_n483), .B1(new_n217), .B2(new_n278), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G264), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n480), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT89), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n479), .A2(new_n291), .B1(new_n485), .B2(G264), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT89), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(new_n484), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(G169), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n487), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G179), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n475), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(G190), .B1(new_n488), .B2(new_n491), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n493), .A2(G200), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n468), .B(new_n474), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n485), .A2(G257), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n484), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n380), .A2(new_n382), .A3(G250), .A4(G1698), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n380), .A2(new_n382), .A3(G244), .A4(new_n285), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n504), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n507), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT82), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n506), .A2(KEYINPUT82), .A3(new_n507), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT83), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n291), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n506), .A2(new_n507), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n505), .A2(new_n504), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n506), .A2(KEYINPUT82), .A3(new_n507), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT82), .B1(new_n506), .B2(new_n507), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n516), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(KEYINPUT83), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n503), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n294), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT6), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n524), .A2(G97), .A3(G107), .ZN(new_n525));
  INV_X1    g0325(.A(G97), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(KEYINPUT6), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n362), .A2(KEYINPUT80), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n362), .A2(KEYINPUT80), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n525), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g0330(.A(KEYINPUT80), .B(G107), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n526), .A2(new_n362), .A3(KEYINPUT6), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n524), .A2(G97), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(new_n534), .A3(new_n215), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n260), .A2(G77), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT81), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT81), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n539), .A3(new_n536), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n386), .A2(G107), .A3(new_n388), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n248), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n267), .A2(new_n526), .ZN(new_n544));
  INV_X1    g0344(.A(new_n473), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(new_n526), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n279), .B1(new_n520), .B2(KEYINPUT83), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n513), .A2(new_n514), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n296), .A3(new_n503), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n523), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n546), .B1(new_n542), .B2(new_n248), .ZN(new_n554));
  OAI211_X1 g0354(.A(G190), .B(new_n503), .C1(new_n515), .C2(new_n521), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n502), .B1(new_n549), .B2(new_n550), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n425), .ZN(new_n557));
  AND2_X1   g0357(.A1(KEYINPUT5), .A2(G41), .ZN(new_n558));
  NOR2_X1   g0358(.A1(KEYINPUT5), .A2(G41), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n483), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(KEYINPUT86), .A3(G270), .A4(new_n279), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n561), .A2(new_n484), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n381), .A2(G33), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n379), .A2(KEYINPUT3), .ZN(new_n564));
  OAI21_X1  g0364(.A(G303), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n380), .A2(new_n382), .A3(G264), .A4(G1698), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n380), .A2(new_n382), .A3(G257), .A4(new_n285), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n291), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n560), .A2(G270), .A3(new_n279), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT86), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n562), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G116), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n267), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n268), .A2(G116), .A3(new_n472), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n379), .A2(G97), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n213), .A2(new_n577), .A3(new_n214), .A4(new_n504), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n247), .A2(new_n216), .B1(G20), .B2(new_n574), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n578), .A2(KEYINPUT20), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT20), .B1(new_n578), .B2(new_n579), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n575), .B(new_n576), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n573), .A2(G169), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT21), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n572), .A2(new_n484), .A3(new_n561), .ZN(new_n586));
  INV_X1    g0386(.A(new_n569), .ZN(new_n587));
  OAI21_X1  g0387(.A(G200), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n582), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n562), .A2(new_n427), .A3(new_n569), .A4(new_n572), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n296), .B1(new_n568), .B2(new_n291), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n582), .A2(new_n572), .A3(new_n562), .A4(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n573), .A2(KEYINPUT21), .A3(G169), .A4(new_n582), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n585), .A2(new_n591), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n213), .A2(G33), .A3(G97), .A4(new_n214), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT19), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n251), .A2(new_n284), .A3(G68), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g0400(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n601));
  NAND2_X1  g0401(.A1(G33), .A2(G97), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT74), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(KEYINPUT74), .A2(G33), .A3(G97), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(KEYINPUT19), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n601), .B1(new_n606), .B2(new_n251), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n248), .B1(new_n600), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n351), .A2(new_n267), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n473), .A2(new_n352), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n380), .A2(new_n382), .A3(G238), .A4(new_n285), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n380), .A2(new_n382), .A3(G244), .A4(G1698), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n454), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n291), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n279), .A2(G274), .A3(new_n483), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n205), .A2(G45), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n617), .B(G250), .C1(new_n290), .C2(new_n216), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n615), .A2(new_n620), .A3(new_n296), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT84), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n615), .A2(new_n620), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n294), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n614), .B2(new_n291), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(KEYINPUT84), .A3(new_n296), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n611), .A2(new_n623), .A3(new_n625), .A4(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT85), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n626), .B2(G190), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(new_n629), .A3(G190), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n215), .B1(new_n316), .B2(KEYINPUT19), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n599), .B(new_n598), .C1(new_n634), .C2(new_n601), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n635), .A2(new_n248), .B1(new_n267), .B2(new_n351), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n624), .A2(new_n303), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n473), .A2(G87), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n628), .B1(new_n633), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n595), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n500), .A2(new_n553), .A3(new_n557), .A4(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n445), .A2(new_n642), .ZN(G372));
  INV_X1    g0443(.A(new_n343), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n371), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n434), .B1(new_n645), .B2(new_n444), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n411), .A2(new_n413), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n421), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT18), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n421), .A2(new_n422), .A3(new_n647), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n310), .B2(new_n309), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n299), .ZN(new_n654));
  INV_X1    g0454(.A(new_n445), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n553), .A2(new_n557), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n626), .A2(G190), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n636), .A2(new_n637), .A3(new_n638), .A4(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n611), .A2(new_n625), .A3(new_n621), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n468), .A2(new_n474), .B1(new_n492), .B2(new_n494), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n585), .A2(new_n593), .A3(new_n594), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n499), .B(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT26), .B1(new_n553), .B2(new_n640), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n659), .A2(KEYINPUT90), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT90), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n611), .A2(new_n667), .A3(new_n625), .A4(new_n621), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n660), .A2(new_n523), .A3(new_n552), .A4(new_n548), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT26), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n664), .A2(new_n665), .A3(new_n670), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n655), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n654), .A2(new_n674), .ZN(G369));
  NAND2_X1  g0475(.A1(new_n251), .A2(new_n469), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n589), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n662), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n595), .B2(new_n683), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G330), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n475), .A2(new_n681), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n500), .A2(new_n690), .B1(new_n661), .B2(new_n681), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n496), .A2(new_n499), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n662), .A2(new_n682), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n694), .A2(new_n695), .B1(new_n496), .B2(new_n681), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT91), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n209), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n601), .A2(new_n574), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n700), .A2(new_n205), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n219), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(new_n700), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT92), .Z(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n656), .A2(new_n663), .B1(KEYINPUT26), .B2(new_n671), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n665), .A2(new_n670), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n709), .A2(KEYINPUT29), .A3(new_n681), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n671), .A2(KEYINPUT26), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n554), .B1(new_n294), .B2(new_n522), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT26), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n611), .A2(new_n625), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n623), .A2(new_n627), .ZN(new_n715));
  INV_X1    g0515(.A(new_n632), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n630), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n608), .A2(new_n609), .A3(new_n638), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n626), .A2(new_n302), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n714), .A2(new_n715), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n712), .A2(new_n713), .A3(new_n721), .A4(new_n552), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n669), .A2(KEYINPUT94), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT94), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n666), .A2(new_n724), .A3(new_n668), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n711), .A2(new_n722), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT95), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n711), .A2(new_n722), .A3(new_n726), .A4(KEYINPUT95), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(new_n664), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n682), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n710), .B1(new_n732), .B2(KEYINPUT29), .ZN(new_n733));
  INV_X1    g0533(.A(new_n595), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(new_n496), .A3(new_n721), .A4(new_n499), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n656), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n569), .A2(G179), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT93), .B1(new_n738), .B2(new_n586), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT93), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n592), .A2(new_n562), .A3(new_n740), .A4(new_n572), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n489), .A2(new_n626), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n737), .B1(new_n522), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n741), .A2(new_n742), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n556), .A2(new_n745), .A3(KEYINPUT30), .A4(new_n739), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n493), .A2(G179), .A3(new_n626), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n522), .A2(new_n573), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n744), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n749), .A2(new_n681), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n736), .A2(new_n682), .B1(new_n750), .B2(KEYINPUT31), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n681), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT31), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n687), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n733), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n706), .B1(new_n758), .B2(G1), .ZN(G364));
  INV_X1    g0559(.A(new_n700), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n215), .A2(new_n266), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G45), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n760), .A2(G1), .A3(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT96), .Z(new_n764));
  NOR2_X1   g0564(.A1(new_n699), .A2(new_n383), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G355), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G116), .B2(new_n209), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n699), .A2(new_n284), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n482), .B2(new_n703), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n242), .A2(new_n482), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n216), .B1(G20), .B2(new_n294), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n764), .B1(new_n772), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n302), .A2(G179), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n206), .A2(new_n300), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n403), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n251), .A2(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n780), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n383), .B(new_n783), .C1(G107), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT97), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G179), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT32), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n251), .A2(new_n296), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n795), .A2(new_n300), .A3(G200), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n795), .A2(new_n425), .A3(new_n427), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n797), .A2(G68), .B1(new_n798), .B2(G58), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n251), .B1(G190), .B2(new_n789), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n526), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n795), .A2(G200), .A3(new_n427), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n792), .A2(new_n793), .B1(new_n269), .B2(new_n802), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n251), .A2(new_n296), .A3(G190), .A4(G200), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n801), .B(new_n803), .C1(G77), .C2(new_n804), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n788), .A2(new_n794), .A3(new_n799), .A4(new_n805), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n807));
  INV_X1    g0607(.A(new_n798), .ZN(new_n808));
  INV_X1    g0608(.A(G322), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  INV_X1    g0610(.A(new_n804), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n808), .A2(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT33), .B(G317), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(new_n797), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n786), .A2(G283), .ZN(new_n815));
  INV_X1    g0615(.A(new_n790), .ZN(new_n816));
  INV_X1    g0616(.A(new_n800), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n816), .A2(G329), .B1(new_n817), .B2(G294), .ZN(new_n818));
  INV_X1    g0618(.A(G303), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n383), .B1(new_n782), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n802), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(G326), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n814), .A2(new_n815), .A3(new_n818), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n807), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n779), .B1(new_n825), .B2(new_n776), .ZN(new_n826));
  INV_X1    g0626(.A(new_n775), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n685), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n686), .A2(new_n687), .ZN(new_n829));
  INV_X1    g0629(.A(new_n764), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n689), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  NAND2_X1  g0633(.A1(new_n673), .A2(new_n682), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n359), .A2(new_n681), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n371), .A2(new_n374), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n359), .A2(new_n369), .A3(new_n370), .A4(new_n681), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n834), .B(new_n838), .ZN(new_n839));
  OR3_X1    g0639(.A1(new_n839), .A2(KEYINPUT100), .A3(new_n755), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT100), .B1(new_n839), .B2(new_n755), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n764), .B1(new_n839), .B2(new_n755), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n776), .ZN(new_n844));
  INV_X1    g0644(.A(G294), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n808), .A2(new_n845), .B1(new_n819), .B2(new_n802), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G116), .B2(new_n804), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n284), .B(new_n801), .C1(new_n797), .C2(G283), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n786), .A2(G87), .ZN(new_n849));
  INV_X1    g0649(.A(new_n782), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n816), .A2(G311), .B1(new_n850), .B2(G107), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n847), .A2(new_n848), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n786), .A2(G68), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n253), .B2(new_n800), .C1(new_n854), .C2(new_n790), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n383), .B(new_n855), .C1(G50), .C2(new_n850), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n798), .A2(G143), .B1(G159), .B2(new_n804), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n857), .B1(new_n858), .B2(new_n802), .C1(new_n859), .C2(new_n796), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT34), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n860), .A2(new_n861), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n852), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n844), .B1(new_n865), .B2(KEYINPUT99), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(KEYINPUT99), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n776), .A2(new_n773), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n830), .B1(new_n202), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n867), .B(new_n869), .C1(new_n774), .C2(new_n838), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n843), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT101), .Z(G384));
  NAND2_X1  g0672(.A1(new_n530), .A2(new_n534), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT102), .Z(new_n874));
  AOI211_X1 g0674(.A(new_n574), .B(new_n218), .C1(new_n874), .C2(KEYINPUT35), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(KEYINPUT35), .B2(new_n874), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT36), .ZN(new_n877));
  OAI21_X1  g0677(.A(G77), .B1(new_n253), .B2(new_n332), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n878), .A2(new_n219), .B1(G50), .B2(new_n332), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(G1), .A3(new_n266), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT103), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT39), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT16), .B1(new_n397), .B2(new_n391), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n417), .B1(new_n420), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n679), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n424), .B2(new_n434), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n421), .A2(new_n409), .A3(new_n414), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n421), .A2(new_n886), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .A4(new_n430), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n885), .B1(new_n647), .B2(new_n886), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n893), .A2(new_n430), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n892), .B1(new_n894), .B2(new_n891), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n890), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n651), .B2(new_n434), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n648), .A2(new_n890), .A3(new_n430), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n892), .B1(new_n899), .B2(new_n891), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n883), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n888), .A2(new_n895), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n444), .A2(new_n681), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n902), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n341), .A2(new_n681), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n441), .A2(new_n442), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n437), .A2(new_n439), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n910), .B1(new_n913), .B2(new_n347), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n343), .A2(new_n910), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n443), .B2(new_n341), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n682), .B(new_n838), .C1(new_n707), .C2(new_n708), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n371), .A2(new_n681), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n917), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n905), .A2(new_n906), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n651), .A2(new_n679), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n909), .B1(new_n925), .B2(KEYINPUT104), .ZN(new_n926));
  INV_X1    g0726(.A(new_n924), .ZN(new_n927));
  AOI211_X1 g0727(.A(KEYINPUT104), .B(new_n927), .C1(new_n921), .C2(new_n922), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n654), .B1(new_n733), .B2(new_n445), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n896), .A2(new_n901), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n838), .B1(new_n914), .B2(new_n916), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT105), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n749), .B2(new_n681), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n749), .A2(new_n937), .A3(new_n681), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(new_n753), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n936), .B1(new_n751), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n933), .B1(new_n935), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT40), .B1(new_n905), .B2(new_n906), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n944), .A2(new_n942), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n642), .B2(new_n681), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n749), .A2(new_n937), .A3(new_n681), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n949), .A2(new_n938), .A3(KEYINPUT31), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n655), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n946), .A2(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(G330), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n932), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n205), .B2(new_n761), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n932), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n882), .B1(new_n956), .B2(new_n957), .ZN(G367));
  NAND2_X1  g0758(.A1(new_n718), .A2(new_n681), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n670), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(new_n660), .B2(new_n959), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT109), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n553), .B(new_n557), .C1(new_n554), .C2(new_n682), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n712), .A2(new_n552), .A3(new_n681), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n969), .A2(new_n500), .A3(new_n662), .A4(new_n682), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT42), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n553), .B1(new_n967), .B2(new_n496), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n682), .B1(new_n972), .B2(KEYINPUT107), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(KEYINPUT107), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT43), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n961), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT108), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n964), .A2(new_n965), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n966), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n965), .B(new_n964), .C1(new_n975), .C2(new_n978), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n981), .A2(new_n692), .A3(new_n969), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  INV_X1    g0784(.A(new_n969), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(new_n693), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n700), .B(KEYINPUT41), .Z(new_n987));
  NOR2_X1   g0787(.A1(new_n697), .A2(new_n969), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n697), .A2(new_n969), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n692), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n691), .A2(new_n695), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n694), .B2(new_n695), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(new_n689), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n757), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n989), .A2(new_n693), .A3(new_n992), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n994), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n987), .B1(new_n1000), .B2(new_n758), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n762), .A2(G1), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n983), .B(new_n986), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n961), .A2(new_n775), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n238), .A2(new_n769), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n778), .B1(new_n699), .B2(new_n352), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n830), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n850), .A2(G116), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT46), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1008), .A2(new_n1009), .B1(G303), .B2(new_n798), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n1009), .B2(new_n1008), .C1(new_n845), .C2(new_n796), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n786), .A2(G97), .B1(new_n817), .B2(G107), .ZN(new_n1012));
  INV_X1    g0812(.A(G317), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1012), .B(new_n383), .C1(new_n1013), .C2(new_n790), .ZN(new_n1014));
  INV_X1    g0814(.A(G283), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n811), .A2(new_n1015), .B1(new_n802), .B2(new_n810), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1011), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n798), .A2(G150), .B1(G50), .B2(new_n804), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n791), .B2(new_n796), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n850), .A2(G58), .B1(new_n817), .B2(G68), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n858), .B2(new_n790), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n821), .A2(G143), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n786), .A2(G77), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(new_n1023), .A3(new_n284), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1019), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1017), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT47), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1004), .B(new_n1007), .C1(new_n1027), .C2(new_n844), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1003), .A2(new_n1028), .ZN(G387));
  NAND2_X1  g0829(.A1(new_n757), .A2(new_n997), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1030), .A2(KEYINPUT114), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n998), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(KEYINPUT114), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1031), .A2(new_n700), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n257), .A2(new_n269), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT50), .Z(new_n1036));
  AOI211_X1 g0836(.A(G45), .B(new_n701), .C1(G68), .C2(G77), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n769), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n234), .B2(new_n482), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n765), .A2(new_n701), .B1(new_n362), .B2(new_n699), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n778), .B1(new_n1041), .B2(KEYINPUT110), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT110), .B2(new_n1041), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n764), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n798), .A2(G317), .B1(G303), .B2(new_n804), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n810), .B2(new_n796), .C1(new_n809), .C2(new_n802), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n782), .A2(new_n845), .B1(new_n800), .B2(new_n1015), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT111), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n284), .B1(new_n816), .B2(G326), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n574), .B2(new_n785), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT112), .Z(new_n1058));
  NAND3_X1  g0858(.A1(new_n1054), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n821), .A2(G159), .B1(G68), .B2(new_n804), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n269), .B2(new_n808), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n850), .A2(G77), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n817), .A2(new_n352), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n859), .C2(new_n790), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n284), .B1(new_n785), .B2(new_n526), .C1(new_n258), .C2(new_n796), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1061), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1044), .B1(new_n1068), .B2(new_n776), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1069), .A2(KEYINPUT113), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1069), .A2(KEYINPUT113), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n691), .C2(new_n775), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n997), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1072), .B1(new_n1002), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1034), .A2(new_n1074), .ZN(G393));
  AND2_X1   g0875(.A1(new_n1000), .A2(new_n700), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n994), .A2(new_n999), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n1032), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n994), .A2(new_n1002), .A3(new_n999), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n808), .A2(new_n810), .B1(new_n1013), .B2(new_n802), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n383), .B1(new_n785), .B2(new_n362), .C1(new_n811), .C2(new_n845), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G303), .B2(new_n797), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n782), .A2(new_n1015), .B1(new_n800), .B2(new_n574), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G322), .B2(new_n816), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1082), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n808), .A2(new_n791), .B1(new_n859), .B2(new_n802), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT51), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n849), .B(new_n284), .C1(new_n269), .C2(new_n796), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n257), .B2(new_n804), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n800), .A2(new_n202), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n782), .A2(new_n332), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(G143), .C2(new_n816), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1089), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n844), .B1(new_n1087), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n769), .A2(new_n245), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n778), .B(new_n1097), .C1(G97), .C2(new_n699), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n1096), .A2(new_n830), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n969), .B2(new_n827), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1080), .A2(KEYINPUT115), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT115), .B1(new_n1080), .B2(new_n1100), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1079), .B1(new_n1102), .B2(new_n1103), .ZN(G390));
  INV_X1    g0904(.A(new_n868), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n821), .A2(G283), .B1(G97), .B2(new_n804), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n362), .B2(new_n796), .C1(new_n574), .C2(new_n808), .ZN(new_n1107));
  NOR4_X1   g0907(.A1(new_n1107), .A2(new_n284), .A3(new_n783), .A4(new_n1092), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n853), .B1(new_n845), .B2(new_n790), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT122), .Z(new_n1110));
  INV_X1    g0910(.A(G128), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n808), .A2(new_n854), .B1(new_n1111), .B2(new_n802), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT121), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n850), .A2(G150), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT53), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n786), .A2(G50), .B1(new_n817), .B2(G159), .ZN(new_n1116));
  INV_X1    g0916(.A(G125), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n284), .C1(new_n1117), .C2(new_n790), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n811), .A2(new_n1119), .B1(new_n796), .B2(new_n858), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1115), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1108), .A2(new_n1110), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n764), .B1(new_n257), .B2(new_n1105), .C1(new_n1122), .C2(new_n844), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n902), .A2(new_n907), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n773), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT116), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n836), .A2(new_n837), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n656), .A2(new_n663), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n727), .B2(new_n728), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n681), .B(new_n1127), .C1(new_n1129), .C2(new_n730), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1126), .B1(new_n1130), .B2(new_n919), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n917), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n731), .A2(new_n682), .A3(new_n838), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(KEYINPUT116), .A3(new_n920), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n934), .A2(new_n908), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n921), .A2(new_n908), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1135), .A2(new_n1136), .B1(new_n1124), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(G330), .B1(new_n950), .B2(new_n948), .ZN(new_n1139));
  OAI21_X1  g0939(.A(KEYINPUT117), .B1(new_n1139), .B2(new_n936), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n687), .B1(new_n751), .B2(new_n941), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT117), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n910), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n345), .A2(new_n346), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n443), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n916), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1127), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1141), .A2(new_n1142), .A3(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1140), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1138), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1137), .A2(new_n1124), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n755), .A2(new_n838), .A3(new_n1132), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1125), .B1(new_n1155), .B2(new_n1002), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT120), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1139), .A2(new_n445), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1159), .B(new_n654), .C1(new_n733), .C2(new_n445), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1161));
  OAI211_X1 g0961(.A(G330), .B(new_n838), .C1(new_n950), .C2(new_n948), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n917), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(KEYINPUT118), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT118), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1162), .A2(new_n1165), .A3(new_n917), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1166), .A2(new_n1153), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1161), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n754), .ZN(new_n1169));
  OAI211_X1 g0969(.A(G330), .B(new_n838), .C1(new_n948), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n917), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1140), .A2(new_n1148), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n918), .A2(new_n920), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI211_X1 g0974(.A(KEYINPUT119), .B(new_n1160), .C1(new_n1168), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT119), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1133), .A2(KEYINPUT116), .A3(new_n920), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT116), .B1(new_n1133), .B2(new_n920), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1164), .A2(new_n1153), .A3(new_n1166), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1174), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1160), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1176), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1157), .B1(new_n1175), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1166), .A2(new_n1153), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1165), .B1(new_n1162), .B2(new_n917), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1187), .A2(new_n1161), .B1(new_n1173), .B2(new_n1172), .ZN(new_n1188));
  OAI21_X1  g0988(.A(KEYINPUT119), .B1(new_n1188), .B2(new_n1160), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1181), .A2(new_n1176), .A3(new_n1182), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(KEYINPUT120), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1155), .B1(new_n1184), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1175), .A2(new_n1183), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1138), .A2(new_n1153), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n700), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1156), .B1(new_n1192), .B2(new_n1196), .ZN(G378));
  OAI21_X1  g0997(.A(new_n1182), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n272), .A2(new_n886), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n311), .B(new_n1199), .Z(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1200), .B(new_n1201), .Z(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(G330), .B1(new_n943), .B2(new_n945), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n926), .B2(new_n929), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n927), .B1(new_n921), .B2(new_n922), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT104), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n908), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1206), .A2(new_n1207), .B1(new_n1208), .B2(new_n1124), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1147), .B1(new_n950), .B2(new_n948), .ZN(new_n1210));
  OAI21_X1  g1010(.A(KEYINPUT40), .B1(new_n1210), .B2(new_n934), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n942), .A2(new_n933), .A3(new_n922), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n687), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1209), .A2(new_n1213), .A3(new_n928), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1203), .B1(new_n1205), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n926), .A2(new_n1204), .A3(new_n929), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1213), .B1(new_n1209), .B2(new_n928), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1217), .A3(new_n1202), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1160), .B1(new_n1221), .B2(new_n1155), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(KEYINPUT57), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n700), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1002), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1202), .A2(new_n773), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n764), .B1(G50), .B2(new_n1105), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n797), .A2(G97), .B1(new_n821), .B2(G116), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n362), .B2(new_n808), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1062), .B1(new_n253), .B2(new_n785), .C1(new_n1015), .C2(new_n790), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n284), .A2(G41), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n800), .B2(new_n332), .C1(new_n811), .C2(new_n351), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1231), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT58), .Z(new_n1236));
  OAI22_X1  g1036(.A1(new_n808), .A2(new_n1111), .B1(new_n858), .B2(new_n811), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1119), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n850), .A2(new_n1238), .B1(new_n817), .B2(G150), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1117), .B2(new_n802), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1237), .B(new_n1240), .C1(G132), .C2(new_n797), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n816), .A2(G124), .ZN(new_n1245));
  AOI211_X1 g1045(.A(G33), .B(G41), .C1(new_n786), .C2(G159), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n269), .B1(G33), .B2(G41), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1236), .B(new_n1247), .C1(new_n1233), .C2(new_n1248), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1249), .A2(KEYINPUT123), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n844), .B1(new_n1249), .B2(KEYINPUT123), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1229), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1228), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1227), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1225), .A2(new_n1255), .ZN(G375));
  OAI22_X1  g1056(.A1(new_n790), .A2(new_n1111), .B1(new_n782), .B2(new_n791), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G50), .B2(new_n817), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n284), .B1(new_n785), .B2(new_n253), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G137), .B2(new_n798), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n804), .A2(G150), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n797), .A2(new_n1238), .B1(new_n821), .B2(G132), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1258), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n821), .A2(G294), .B1(G107), .B2(new_n804), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1015), .B2(new_n808), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1063), .B1(new_n782), .B2(new_n526), .C1(new_n819), .C2(new_n790), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1023), .B(new_n383), .C1(new_n574), .C2(new_n796), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT124), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1263), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1268), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(KEYINPUT124), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n776), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n830), .B1(new_n332), .B2(new_n868), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1273), .B(new_n1274), .C1(new_n1132), .C2(new_n774), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1188), .B2(new_n1226), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1184), .A2(new_n1191), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1160), .B(new_n1174), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1281), .A2(new_n987), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1277), .B1(new_n1279), .B2(new_n1282), .ZN(G381));
  INV_X1    g1083(.A(G375), .ZN(new_n1284));
  INV_X1    g1084(.A(G378), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1103), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1286), .A2(new_n1101), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n871), .B(KEYINPUT101), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(G393), .A2(G396), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(G381), .A2(G387), .A3(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1284), .A2(new_n1285), .A3(new_n1291), .ZN(G407));
  NAND2_X1  g1092(.A1(new_n680), .A2(G213), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1284), .A2(new_n1285), .A3(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(G407), .A2(new_n1295), .A3(G213), .ZN(G409));
  AOI21_X1  g1096(.A(new_n832), .B1(new_n1034), .B2(new_n1074), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1289), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(G390), .B1(new_n1003), .B2(new_n1028), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(G387), .A2(new_n1287), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G387), .A2(new_n1287), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(G390), .A2(new_n1003), .A3(new_n1028), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1298), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(G378), .B(new_n1255), .C1(new_n1220), .C2(new_n1224), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1175), .A2(new_n1183), .A3(new_n1157), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT120), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1195), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n760), .B1(new_n1221), .B2(new_n1155), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1219), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1222), .A2(new_n987), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT125), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1227), .B2(new_n1254), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1216), .A2(new_n1217), .A3(new_n1202), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1202), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1002), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1319), .A2(KEYINPUT125), .A3(new_n1253), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1316), .A2(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1312), .B(new_n1156), .C1(new_n1314), .C2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1307), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT62), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1189), .A2(new_n1190), .A3(new_n1280), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(KEYINPUT60), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n700), .B1(new_n1281), .B2(KEYINPUT60), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(G384), .A3(new_n1277), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1327), .B1(new_n1325), .B2(KEYINPUT60), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1288), .B1(new_n1331), .B2(new_n1276), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1323), .A2(new_n1324), .A3(new_n1293), .A4(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT61), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1294), .B1(new_n1307), .B2(new_n1322), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1294), .A2(KEYINPUT126), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1330), .A2(new_n1332), .A3(new_n1338), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1294), .A2(G2897), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1339), .B(new_n1340), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1335), .B(new_n1336), .C1(new_n1337), .C2(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1324), .B1(new_n1337), .B2(new_n1334), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1306), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  OR2_X1    g1144(.A1(new_n1341), .A2(new_n1337), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1302), .A2(new_n1336), .A3(new_n1305), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1346), .B(KEYINPUT127), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1337), .A2(new_n1334), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT63), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1337), .A2(KEYINPUT63), .A3(new_n1334), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1345), .A2(new_n1347), .A3(new_n1350), .A4(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1344), .A2(new_n1352), .ZN(G405));
  NAND2_X1  g1153(.A1(G375), .A2(new_n1285), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1354), .A2(new_n1307), .A3(new_n1333), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1333), .B1(new_n1354), .B2(new_n1307), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1306), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1354), .A2(new_n1307), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1334), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1360), .A2(new_n1305), .A3(new_n1302), .A4(new_n1355), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1358), .A2(new_n1361), .ZN(G402));
endmodule


