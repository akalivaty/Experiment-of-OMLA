

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777;

  NOR2_X1 U377 ( .A1(n472), .A2(n471), .ZN(n544) );
  NAND2_X1 U378 ( .A1(n597), .A2(n596), .ZN(n642) );
  XNOR2_X1 U379 ( .A(n520), .B(n519), .ZN(n628) );
  XNOR2_X1 U380 ( .A(n469), .B(n468), .ZN(n705) );
  INV_X2 U381 ( .A(G953), .ZN(n754) );
  XNOR2_X1 U382 ( .A(KEYINPUT66), .B(n658), .ZN(n355) );
  AND2_X1 U383 ( .A1(n401), .A2(n400), .ZN(n356) );
  XNOR2_X2 U384 ( .A(G140), .B(KEYINPUT10), .ZN(n441) );
  AND2_X1 U385 ( .A1(n688), .A2(n610), .ZN(n612) );
  XNOR2_X1 U386 ( .A(n395), .B(n402), .ZN(n688) );
  AND2_X2 U387 ( .A1(n544), .A2(n363), .ZN(n634) );
  AND2_X2 U388 ( .A1(n536), .A2(n588), .ZN(n629) );
  XNOR2_X2 U389 ( .A(n573), .B(KEYINPUT1), .ZN(n601) );
  XNOR2_X1 U390 ( .A(n411), .B(n488), .ZN(n394) );
  XNOR2_X2 U391 ( .A(G122), .B(G116), .ZN(n490) );
  INV_X2 U392 ( .A(G131), .ZN(n419) );
  NOR2_X1 U393 ( .A1(G953), .A2(G237), .ZN(n476) );
  INV_X1 U394 ( .A(KEYINPUT64), .ZN(n358) );
  NAND2_X1 U395 ( .A1(n396), .A2(n365), .ZN(n395) );
  NOR2_X1 U396 ( .A1(n638), .A2(n637), .ZN(n645) );
  NAND2_X1 U397 ( .A1(n389), .A2(n388), .ZN(n594) );
  XNOR2_X1 U398 ( .A(n590), .B(n369), .ZN(n611) );
  AND2_X1 U399 ( .A1(n567), .A2(n366), .ZN(n590) );
  AND2_X1 U400 ( .A1(n390), .A2(n392), .ZN(n389) );
  XNOR2_X1 U401 ( .A(n628), .B(n521), .ZN(n378) );
  NAND2_X2 U402 ( .A1(n397), .A2(n356), .ZN(n573) );
  XNOR2_X1 U403 ( .A(n541), .B(KEYINPUT38), .ZN(n549) );
  AND2_X1 U404 ( .A1(n564), .A2(n537), .ZN(n434) );
  XNOR2_X1 U405 ( .A(n484), .B(n483), .ZN(n547) );
  XNOR2_X1 U406 ( .A(n473), .B(n420), .ZN(n411) );
  XNOR2_X1 U407 ( .A(n380), .B(n428), .ZN(n503) );
  XNOR2_X1 U408 ( .A(n509), .B(n421), .ZN(n488) );
  XNOR2_X1 U409 ( .A(n412), .B(KEYINPUT3), .ZN(n380) );
  XNOR2_X1 U410 ( .A(n507), .B(n441), .ZN(n767) );
  XNOR2_X1 U411 ( .A(n490), .B(n489), .ZN(n500) );
  XNOR2_X1 U412 ( .A(KEYINPUT4), .B(G137), .ZN(n420) );
  NAND2_X1 U413 ( .A1(n717), .A2(n601), .ZN(n602) );
  NOR2_X4 U414 ( .A1(n357), .A2(n715), .ZN(n692) );
  XNOR2_X2 U415 ( .A(n359), .B(n358), .ZN(n357) );
  NAND2_X1 U416 ( .A1(n360), .A2(n355), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n655), .B(n361), .ZN(n360) );
  INV_X1 U418 ( .A(KEYINPUT85), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n404), .B(n403), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n404), .B(n403), .ZN(n606) );
  XNOR2_X1 U421 ( .A(n591), .B(n512), .ZN(n683) );
  AND2_X1 U422 ( .A1(n608), .A2(n518), .ZN(n363) );
  NOR2_X2 U423 ( .A1(n679), .A2(n708), .ZN(n681) );
  BUF_X1 U424 ( .A(n543), .Z(n541) );
  NOR2_X2 U425 ( .A1(n686), .A2(n708), .ZN(n687) );
  XNOR2_X1 U426 ( .A(n517), .B(n516), .ZN(n543) );
  NOR2_X2 U427 ( .A1(n673), .A2(n708), .ZN(n674) );
  NOR2_X2 U428 ( .A1(n543), .A2(n739), .ZN(n520) );
  INV_X1 U429 ( .A(n652), .ZN(n408) );
  XNOR2_X1 U430 ( .A(G902), .B(KEYINPUT91), .ZN(n436) );
  INV_X1 U431 ( .A(KEYINPUT102), .ZN(n413) );
  XNOR2_X1 U432 ( .A(G113), .B(G116), .ZN(n425) );
  XOR2_X1 U433 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n423) );
  AND2_X1 U434 ( .A1(n659), .A2(n368), .ZN(n666) );
  NOR2_X1 U435 ( .A1(n664), .A2(n376), .ZN(n375) );
  NAND2_X1 U436 ( .A1(n549), .A2(n537), .ZN(n377) );
  NAND2_X1 U437 ( .A1(n399), .A2(n495), .ZN(n398) );
  INV_X1 U438 ( .A(KEYINPUT0), .ZN(n403) );
  BUF_X1 U439 ( .A(n601), .Z(n718) );
  AND2_X1 U440 ( .A1(n407), .A2(n513), .ZN(n406) );
  NAND2_X1 U441 ( .A1(n408), .A2(KEYINPUT76), .ZN(n407) );
  NOR2_X1 U442 ( .A1(n613), .A2(KEYINPUT44), .ZN(n614) );
  INV_X1 U443 ( .A(n661), .ZN(n376) );
  INV_X1 U444 ( .A(G469), .ZN(n399) );
  NAND2_X1 U445 ( .A1(G902), .A2(G469), .ZN(n400) );
  INV_X1 U446 ( .A(n549), .ZN(n740) );
  XOR2_X1 U447 ( .A(n515), .B(KEYINPUT93), .Z(n516) );
  NOR2_X1 U448 ( .A1(G902), .A2(n670), .ZN(n484) );
  XNOR2_X1 U449 ( .A(n469), .B(n430), .ZN(n676) );
  INV_X1 U450 ( .A(G107), .ZN(n489) );
  XNOR2_X1 U451 ( .A(G119), .B(G137), .ZN(n447) );
  XNOR2_X1 U452 ( .A(n473), .B(n474), .ZN(n475) );
  XNOR2_X1 U453 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n474) );
  XOR2_X1 U454 ( .A(G122), .B(KEYINPUT99), .Z(n478) );
  XNOR2_X1 U455 ( .A(G107), .B(G104), .ZN(n462) );
  XNOR2_X1 U456 ( .A(G101), .B(G110), .ZN(n463) );
  INV_X1 U457 ( .A(G140), .ZN(n464) );
  XNOR2_X1 U458 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n504) );
  XNOR2_X1 U459 ( .A(KEYINPUT89), .B(KEYINPUT4), .ZN(n508) );
  XNOR2_X1 U460 ( .A(n383), .B(n382), .ZN(n715) );
  INV_X1 U461 ( .A(KEYINPUT77), .ZN(n382) );
  NOR2_X1 U462 ( .A1(n377), .A2(n738), .ZN(n550) );
  XNOR2_X1 U463 ( .A(n385), .B(n384), .ZN(n555) );
  INV_X1 U464 ( .A(KEYINPUT39), .ZN(n384) );
  NAND2_X1 U465 ( .A1(n730), .A2(n370), .ZN(n392) );
  XNOR2_X1 U466 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U467 ( .A1(n386), .A2(n568), .ZN(n393) );
  XNOR2_X1 U468 ( .A(n577), .B(KEYINPUT97), .ZN(n386) );
  BUF_X1 U469 ( .A(n554), .Z(n596) );
  XNOR2_X1 U470 ( .A(n440), .B(n439), .ZN(n454) );
  AND2_X1 U471 ( .A1(n693), .A2(n495), .ZN(n453) );
  XNOR2_X1 U472 ( .A(n438), .B(KEYINPUT25), .ZN(n439) );
  INV_X1 U473 ( .A(KEYINPUT22), .ZN(n379) );
  BUF_X1 U474 ( .A(n692), .Z(n701) );
  NOR2_X1 U475 ( .A1(n754), .A2(G952), .ZN(n708) );
  XNOR2_X1 U476 ( .A(n630), .B(n631), .ZN(n374) );
  INV_X1 U477 ( .A(KEYINPUT35), .ZN(n402) );
  INV_X1 U478 ( .A(n393), .ZN(n595) );
  AND2_X1 U479 ( .A1(n652), .A2(n653), .ZN(n364) );
  XNOR2_X1 U480 ( .A(KEYINPUT79), .B(n609), .ZN(n365) );
  INV_X1 U481 ( .A(G902), .ZN(n495) );
  AND2_X1 U482 ( .A1(n514), .A2(G214), .ZN(n739) );
  AND2_X1 U483 ( .A1(n589), .A2(n603), .ZN(n366) );
  AND2_X1 U484 ( .A1(n598), .A2(n603), .ZN(n367) );
  AND2_X1 U485 ( .A1(n660), .A2(KEYINPUT2), .ZN(n368) );
  XNOR2_X1 U486 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n369) );
  XNOR2_X1 U487 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n370) );
  XOR2_X1 U488 ( .A(KEYINPUT80), .B(KEYINPUT34), .Z(n371) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n656) );
  XOR2_X1 U490 ( .A(G119), .B(KEYINPUT127), .Z(n372) );
  NAND2_X1 U491 ( .A1(n373), .A2(n364), .ZN(n409) );
  NOR2_X1 U492 ( .A1(n373), .A2(n653), .ZN(n410) );
  AND2_X2 U493 ( .A1(n373), .A2(n652), .ZN(n659) );
  AND2_X1 U494 ( .A1(n373), .A2(n375), .ZN(n665) );
  XNOR2_X2 U495 ( .A(n650), .B(KEYINPUT48), .ZN(n373) );
  XNOR2_X1 U496 ( .A(n437), .B(KEYINPUT20), .ZN(n455) );
  AND2_X1 U497 ( .A1(n378), .A2(n527), .ZN(n763) );
  XNOR2_X2 U498 ( .A(n605), .B(n604), .ZN(n752) );
  XNOR2_X1 U499 ( .A(n547), .B(KEYINPUT100), .ZN(n532) );
  NAND2_X1 U500 ( .A1(n374), .A2(n718), .ZN(n632) );
  NOR2_X2 U501 ( .A1(n603), .A2(n602), .ZN(n605) );
  NOR2_X1 U502 ( .A1(n736), .A2(n377), .ZN(n737) );
  NAND2_X1 U503 ( .A1(n378), .A2(n418), .ZN(n404) );
  AND2_X1 U504 ( .A1(n567), .A2(n367), .ZN(n624) );
  XNOR2_X2 U505 ( .A(n563), .B(n379), .ZN(n567) );
  XNOR2_X2 U506 ( .A(n381), .B(KEYINPUT45), .ZN(n667) );
  NAND2_X1 U507 ( .A1(n617), .A2(n616), .ZN(n381) );
  NAND2_X1 U508 ( .A1(n362), .A2(n391), .ZN(n388) );
  NAND2_X1 U509 ( .A1(n409), .A2(n406), .ZN(n405) );
  XNOR2_X1 U510 ( .A(n607), .B(n371), .ZN(n396) );
  NOR2_X1 U511 ( .A1(n669), .A2(n668), .ZN(n383) );
  NAND2_X1 U512 ( .A1(n544), .A2(n549), .ZN(n385) );
  NAND2_X1 U513 ( .A1(n570), .A2(n370), .ZN(n390) );
  NAND2_X1 U514 ( .A1(n416), .A2(n415), .ZN(n414) );
  NOR2_X2 U515 ( .A1(n523), .A2(n522), .ZN(n533) );
  NOR2_X1 U516 ( .A1(n410), .A2(n405), .ZN(n654) );
  NAND2_X1 U517 ( .A1(n387), .A2(n393), .ZN(n417) );
  INV_X1 U518 ( .A(n594), .ZN(n387) );
  NOR2_X1 U519 ( .A1(n730), .A2(n370), .ZN(n391) );
  XNOR2_X1 U520 ( .A(n611), .B(n372), .ZN(G21) );
  XNOR2_X2 U521 ( .A(n394), .B(G146), .ZN(n469) );
  XNOR2_X1 U522 ( .A(n394), .B(n769), .ZN(n772) );
  OR2_X1 U523 ( .A1(n705), .A2(n398), .ZN(n397) );
  NAND2_X1 U524 ( .A1(n705), .A2(G469), .ZN(n401) );
  XNOR2_X2 U525 ( .A(G119), .B(KEYINPUT92), .ZN(n412) );
  XNOR2_X1 U526 ( .A(n414), .B(n413), .ZN(n600) );
  INV_X1 U527 ( .A(n624), .ZN(n415) );
  NAND2_X1 U528 ( .A1(n417), .A2(n642), .ZN(n416) );
  AND2_X1 U529 ( .A1(n600), .A2(n599), .ZN(n617) );
  BUF_X1 U530 ( .A(n688), .Z(n689) );
  AND2_X1 U531 ( .A1(n749), .A2(n560), .ZN(n418) );
  INV_X1 U532 ( .A(KEYINPUT74), .ZN(n424) );
  XNOR2_X1 U533 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U534 ( .A(n427), .B(n426), .ZN(n429) );
  INV_X1 U535 ( .A(KEYINPUT87), .ZN(n519) );
  INV_X1 U536 ( .A(KEYINPUT19), .ZN(n521) );
  BUF_X1 U537 ( .A(n667), .Z(n710) );
  XNOR2_X2 U538 ( .A(n419), .B(KEYINPUT68), .ZN(n473) );
  XNOR2_X2 U539 ( .A(G128), .B(G143), .ZN(n509) );
  INV_X1 U540 ( .A(G134), .ZN(n421) );
  NAND2_X1 U541 ( .A1(n476), .A2(G210), .ZN(n422) );
  XNOR2_X1 U542 ( .A(n423), .B(n422), .ZN(n427) );
  XNOR2_X1 U543 ( .A(G101), .B(KEYINPUT70), .ZN(n428) );
  XNOR2_X1 U544 ( .A(n503), .B(n429), .ZN(n430) );
  NAND2_X1 U545 ( .A1(n676), .A2(n495), .ZN(n431) );
  XNOR2_X2 U546 ( .A(n431), .B(G472), .ZN(n564) );
  NOR2_X1 U547 ( .A1(G902), .A2(G237), .ZN(n432) );
  XNOR2_X1 U548 ( .A(n432), .B(KEYINPUT73), .ZN(n514) );
  INV_X1 U549 ( .A(n739), .ZN(n537) );
  INV_X1 U550 ( .A(KEYINPUT30), .ZN(n433) );
  XNOR2_X1 U551 ( .A(n434), .B(n433), .ZN(n472) );
  INV_X1 U552 ( .A(KEYINPUT15), .ZN(n435) );
  NAND2_X1 U553 ( .A1(n656), .A2(G234), .ZN(n437) );
  NAND2_X1 U554 ( .A1(n455), .A2(G217), .ZN(n440) );
  XOR2_X1 U555 ( .A(KEYINPUT96), .B(KEYINPUT78), .Z(n438) );
  XNOR2_X2 U556 ( .A(G146), .B(G125), .ZN(n507) );
  XOR2_X1 U557 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n443) );
  XNOR2_X1 U558 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n442) );
  XNOR2_X1 U559 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U560 ( .A(n767), .B(n444), .ZN(n452) );
  NAND2_X1 U561 ( .A1(n754), .A2(G234), .ZN(n446) );
  INV_X1 U562 ( .A(KEYINPUT8), .ZN(n445) );
  XNOR2_X1 U563 ( .A(n446), .B(n445), .ZN(n485) );
  NAND2_X1 U564 ( .A1(n485), .A2(G221), .ZN(n450) );
  XOR2_X1 U565 ( .A(G110), .B(G128), .Z(n448) );
  XNOR2_X1 U566 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U567 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U568 ( .A(n452), .B(n451), .ZN(n693) );
  XNOR2_X2 U569 ( .A(n454), .B(n453), .ZN(n721) );
  INV_X1 U570 ( .A(n721), .ZN(n586) );
  AND2_X1 U571 ( .A1(n455), .A2(G221), .ZN(n456) );
  XNOR2_X1 U572 ( .A(n456), .B(KEYINPUT21), .ZN(n561) );
  NAND2_X1 U573 ( .A1(n586), .A2(n561), .ZN(n574) );
  NAND2_X1 U574 ( .A1(G234), .A2(G237), .ZN(n457) );
  XNOR2_X1 U575 ( .A(n457), .B(KEYINPUT14), .ZN(n749) );
  NAND2_X1 U576 ( .A1(n754), .A2(G952), .ZN(n459) );
  NAND2_X1 U577 ( .A1(G953), .A2(G902), .ZN(n458) );
  NAND2_X1 U578 ( .A1(n459), .A2(n458), .ZN(n559) );
  NAND2_X1 U579 ( .A1(G953), .A2(G900), .ZN(n460) );
  AND2_X1 U580 ( .A1(n559), .A2(n460), .ZN(n461) );
  NAND2_X1 U581 ( .A1(n749), .A2(n461), .ZN(n523) );
  NOR2_X1 U582 ( .A1(n574), .A2(n523), .ZN(n470) );
  XNOR2_X1 U583 ( .A(n463), .B(n462), .ZN(n467) );
  NAND2_X1 U584 ( .A1(n754), .A2(G227), .ZN(n465) );
  XNOR2_X1 U585 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U586 ( .A(n467), .B(n466), .ZN(n468) );
  NAND2_X1 U587 ( .A1(n470), .A2(n573), .ZN(n471) );
  XNOR2_X1 U588 ( .A(n475), .B(n767), .ZN(n482) );
  NAND2_X1 U589 ( .A1(G214), .A2(n476), .ZN(n477) );
  XNOR2_X1 U590 ( .A(n478), .B(n477), .ZN(n480) );
  XNOR2_X2 U591 ( .A(G113), .B(G104), .ZN(n499) );
  XNOR2_X1 U592 ( .A(n499), .B(G143), .ZN(n479) );
  XNOR2_X1 U593 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U594 ( .A(n482), .B(n481), .ZN(n670) );
  XNOR2_X1 U595 ( .A(KEYINPUT13), .B(G475), .ZN(n483) );
  XOR2_X1 U596 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n487) );
  NAND2_X1 U597 ( .A1(G217), .A2(n485), .ZN(n486) );
  XNOR2_X1 U598 ( .A(n487), .B(n486), .ZN(n494) );
  INV_X1 U599 ( .A(n488), .ZN(n492) );
  INV_X1 U600 ( .A(n500), .ZN(n491) );
  XNOR2_X1 U601 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U602 ( .A(n494), .B(n493), .ZN(n697) );
  NAND2_X1 U603 ( .A1(n697), .A2(n495), .ZN(n497) );
  INV_X1 U604 ( .A(G478), .ZN(n496) );
  XNOR2_X1 U605 ( .A(n497), .B(n496), .ZN(n531) );
  INV_X1 U606 ( .A(n531), .ZN(n546) );
  AND2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n608) );
  XNOR2_X1 U608 ( .A(KEYINPUT16), .B(G110), .ZN(n498) );
  XNOR2_X1 U609 ( .A(n499), .B(n498), .ZN(n501) );
  XNOR2_X1 U610 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n502), .B(n503), .ZN(n591) );
  NAND2_X1 U612 ( .A1(n754), .A2(G224), .ZN(n505) );
  XNOR2_X1 U613 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U614 ( .A(n506), .B(n507), .ZN(n511) );
  XNOR2_X1 U615 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U616 ( .A(n511), .B(n510), .ZN(n512) );
  INV_X1 U617 ( .A(n656), .ZN(n513) );
  NOR2_X1 U618 ( .A1(n683), .A2(n513), .ZN(n517) );
  AND2_X1 U619 ( .A1(n514), .A2(G210), .ZN(n515) );
  INV_X1 U620 ( .A(n541), .ZN(n518) );
  XOR2_X1 U621 ( .A(n634), .B(G143), .Z(G45) );
  NAND2_X1 U622 ( .A1(n721), .A2(n561), .ZN(n522) );
  NAND2_X1 U623 ( .A1(n533), .A2(n564), .ZN(n525) );
  XNOR2_X1 U624 ( .A(KEYINPUT103), .B(KEYINPUT28), .ZN(n524) );
  NAND2_X1 U625 ( .A1(n526), .A2(n573), .ZN(n551) );
  INV_X1 U626 ( .A(n551), .ZN(n527) );
  INV_X1 U627 ( .A(n532), .ZN(n528) );
  NAND2_X1 U628 ( .A1(n528), .A2(n546), .ZN(n597) );
  INV_X1 U629 ( .A(n597), .ZN(n578) );
  NAND2_X1 U630 ( .A1(n763), .A2(n578), .ZN(n530) );
  XOR2_X1 U631 ( .A(G128), .B(KEYINPUT29), .Z(n529) );
  XNOR2_X1 U632 ( .A(n530), .B(n529), .ZN(G30) );
  NAND2_X1 U633 ( .A1(n532), .A2(n531), .ZN(n554) );
  INV_X1 U634 ( .A(n554), .ZN(n534) );
  AND2_X1 U635 ( .A1(n534), .A2(n533), .ZN(n536) );
  INV_X1 U636 ( .A(KEYINPUT6), .ZN(n535) );
  XNOR2_X1 U637 ( .A(n564), .B(n535), .ZN(n588) );
  INV_X1 U638 ( .A(n629), .ZN(n539) );
  INV_X1 U639 ( .A(n718), .ZN(n587) );
  NAND2_X1 U640 ( .A1(n587), .A2(n537), .ZN(n538) );
  NOR2_X1 U641 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U642 ( .A(KEYINPUT43), .B(n540), .Z(n542) );
  NAND2_X1 U643 ( .A1(n542), .A2(n541), .ZN(n661) );
  XNOR2_X1 U644 ( .A(n661), .B(G140), .ZN(G42) );
  XNOR2_X1 U645 ( .A(G134), .B(KEYINPUT112), .ZN(n545) );
  NOR2_X1 U646 ( .A1(n555), .A2(n597), .ZN(n651) );
  XOR2_X1 U647 ( .A(n545), .B(n651), .Z(G36) );
  NOR2_X1 U648 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U649 ( .A(n548), .B(KEYINPUT101), .ZN(n738) );
  XNOR2_X1 U650 ( .A(n550), .B(KEYINPUT41), .ZN(n733) );
  NOR2_X1 U651 ( .A1(n733), .A2(n551), .ZN(n553) );
  XNOR2_X1 U652 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n552) );
  XNOR2_X1 U653 ( .A(n553), .B(n552), .ZN(n625) );
  XNOR2_X1 U654 ( .A(n625), .B(G137), .ZN(G39) );
  NOR2_X1 U655 ( .A1(n555), .A2(n596), .ZN(n557) );
  XOR2_X1 U656 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n556) );
  XNOR2_X1 U657 ( .A(n557), .B(n556), .ZN(n626) );
  XNOR2_X1 U658 ( .A(n626), .B(G131), .ZN(G33) );
  NAND2_X1 U659 ( .A1(G953), .A2(G898), .ZN(n558) );
  AND2_X1 U660 ( .A1(n559), .A2(n558), .ZN(n560) );
  INV_X1 U661 ( .A(n561), .ZN(n722) );
  NOR2_X1 U662 ( .A1(n738), .A2(n722), .ZN(n562) );
  NAND2_X1 U663 ( .A1(n606), .A2(n562), .ZN(n563) );
  INV_X1 U664 ( .A(n564), .ZN(n568) );
  NAND2_X1 U665 ( .A1(n568), .A2(n721), .ZN(n565) );
  NOR2_X1 U666 ( .A1(n718), .A2(n565), .ZN(n566) );
  NAND2_X1 U667 ( .A1(n567), .A2(n566), .ZN(n610) );
  XNOR2_X1 U668 ( .A(n610), .B(G110), .ZN(G12) );
  INV_X1 U669 ( .A(n362), .ZN(n570) );
  INV_X1 U670 ( .A(n574), .ZN(n717) );
  INV_X1 U671 ( .A(n568), .ZN(n727) );
  AND2_X1 U672 ( .A1(n717), .A2(n727), .ZN(n569) );
  NAND2_X1 U673 ( .A1(n718), .A2(n569), .ZN(n730) );
  INV_X1 U674 ( .A(n596), .ZN(n762) );
  NAND2_X1 U675 ( .A1(n594), .A2(n762), .ZN(n571) );
  XNOR2_X1 U676 ( .A(n571), .B(G113), .ZN(G15) );
  NAND2_X1 U677 ( .A1(n594), .A2(n578), .ZN(n572) );
  XNOR2_X1 U678 ( .A(n572), .B(G116), .ZN(G18) );
  INV_X1 U679 ( .A(n573), .ZN(n575) );
  NOR2_X1 U680 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U681 ( .A1(n362), .A2(n576), .ZN(n577) );
  NAND2_X1 U682 ( .A1(n595), .A2(n578), .ZN(n583) );
  XOR2_X1 U683 ( .A(KEYINPUT27), .B(KEYINPUT109), .Z(n580) );
  XNOR2_X1 U684 ( .A(G107), .B(KEYINPUT26), .ZN(n579) );
  XNOR2_X1 U685 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U686 ( .A(KEYINPUT108), .B(n581), .Z(n582) );
  XNOR2_X1 U687 ( .A(n583), .B(n582), .ZN(G9) );
  NAND2_X1 U688 ( .A1(n595), .A2(n762), .ZN(n585) );
  XOR2_X1 U689 ( .A(G104), .B(KEYINPUT107), .Z(n584) );
  XNOR2_X1 U690 ( .A(n585), .B(n584), .ZN(G6) );
  NOR2_X1 U691 ( .A1(n587), .A2(n586), .ZN(n589) );
  INV_X1 U692 ( .A(n588), .ZN(n603) );
  INV_X1 U693 ( .A(G898), .ZN(n592) );
  NAND2_X1 U694 ( .A1(n592), .A2(G953), .ZN(n593) );
  NAND2_X1 U695 ( .A1(n591), .A2(n593), .ZN(n623) );
  INV_X1 U696 ( .A(n642), .ZN(n736) );
  NOR2_X1 U697 ( .A1(n718), .A2(n721), .ZN(n598) );
  INV_X1 U698 ( .A(KEYINPUT72), .ZN(n613) );
  NAND2_X1 U699 ( .A1(n613), .A2(KEYINPUT44), .ZN(n599) );
  XNOR2_X1 U700 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n604) );
  NAND2_X1 U701 ( .A1(n752), .A2(n606), .ZN(n607) );
  INV_X1 U702 ( .A(n608), .ZN(n609) );
  NAND2_X1 U703 ( .A1(n612), .A2(n611), .ZN(n615) );
  XNOR2_X1 U704 ( .A(n615), .B(n614), .ZN(n616) );
  NAND2_X1 U705 ( .A1(n710), .A2(n754), .ZN(n621) );
  NAND2_X1 U706 ( .A1(G953), .A2(G224), .ZN(n618) );
  XNOR2_X1 U707 ( .A(KEYINPUT61), .B(n618), .ZN(n619) );
  NAND2_X1 U708 ( .A1(n619), .A2(G898), .ZN(n620) );
  NAND2_X1 U709 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U710 ( .A(n623), .B(n622), .Z(G69) );
  XOR2_X1 U711 ( .A(G101), .B(n624), .Z(G3) );
  NAND2_X1 U712 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U713 ( .A(n627), .B(KEYINPUT46), .ZN(n649) );
  INV_X1 U714 ( .A(KEYINPUT36), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U716 ( .A(KEYINPUT106), .B(n632), .Z(n691) );
  INV_X1 U717 ( .A(KEYINPUT47), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n642), .A2(n636), .ZN(n633) );
  NOR2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U720 ( .A(n635), .B(KEYINPUT83), .ZN(n638) );
  NOR2_X1 U721 ( .A1(n763), .A2(n636), .ZN(n637) );
  NOR2_X1 U722 ( .A1(KEYINPUT47), .A2(KEYINPUT67), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n763), .A2(n639), .ZN(n641) );
  NAND2_X1 U724 ( .A1(KEYINPUT67), .A2(KEYINPUT47), .ZN(n640) );
  NAND2_X1 U725 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U728 ( .A1(n691), .A2(n646), .ZN(n647) );
  XNOR2_X1 U729 ( .A(n647), .B(KEYINPUT69), .ZN(n648) );
  NOR2_X2 U730 ( .A1(n649), .A2(n648), .ZN(n650) );
  INV_X1 U731 ( .A(n651), .ZN(n662) );
  AND2_X1 U732 ( .A1(n661), .A2(n662), .ZN(n652) );
  INV_X1 U733 ( .A(KEYINPUT76), .ZN(n653) );
  NAND2_X1 U734 ( .A1(n654), .A2(n667), .ZN(n655) );
  XOR2_X1 U735 ( .A(n656), .B(KEYINPUT86), .Z(n657) );
  NAND2_X1 U736 ( .A1(n657), .A2(KEYINPUT2), .ZN(n658) );
  INV_X1 U737 ( .A(KEYINPUT81), .ZN(n660) );
  NAND2_X1 U738 ( .A1(n662), .A2(KEYINPUT2), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n663), .A2(KEYINPUT81), .ZN(n664) );
  NOR2_X1 U740 ( .A1(n666), .A2(n665), .ZN(n669) );
  INV_X1 U741 ( .A(n667), .ZN(n668) );
  NAND2_X1 U742 ( .A1(n692), .A2(G475), .ZN(n672) );
  XOR2_X1 U743 ( .A(KEYINPUT59), .B(n670), .Z(n671) );
  XNOR2_X1 U744 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U745 ( .A(n674), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U746 ( .A1(n692), .A2(G472), .ZN(n678) );
  XOR2_X1 U747 ( .A(KEYINPUT90), .B(KEYINPUT62), .Z(n675) );
  XNOR2_X1 U748 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n678), .B(n677), .ZN(n679) );
  XOR2_X1 U750 ( .A(KEYINPUT88), .B(KEYINPUT63), .Z(n680) );
  XNOR2_X1 U751 ( .A(n681), .B(n680), .ZN(G57) );
  NAND2_X1 U752 ( .A1(n692), .A2(G210), .ZN(n685) );
  XOR2_X1 U753 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n682) );
  XNOR2_X1 U754 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U756 ( .A(n687), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U757 ( .A(n689), .B(G122), .ZN(G24) );
  XNOR2_X1 U758 ( .A(G125), .B(KEYINPUT37), .ZN(n690) );
  XNOR2_X1 U759 ( .A(n691), .B(n690), .ZN(G27) );
  NAND2_X1 U760 ( .A1(n701), .A2(G217), .ZN(n695) );
  XOR2_X1 U761 ( .A(KEYINPUT122), .B(n693), .Z(n694) );
  XNOR2_X1 U762 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n696), .A2(n708), .ZN(G66) );
  NAND2_X1 U764 ( .A1(n701), .A2(G478), .ZN(n699) );
  XNOR2_X1 U765 ( .A(n697), .B(KEYINPUT121), .ZN(n698) );
  XNOR2_X1 U766 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U767 ( .A1(n700), .A2(n708), .ZN(G63) );
  NAND2_X1 U768 ( .A1(n701), .A2(G469), .ZN(n707) );
  XNOR2_X1 U769 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n703) );
  XNOR2_X1 U770 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n702) );
  XNOR2_X1 U771 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U772 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U773 ( .A(n707), .B(n706), .ZN(n709) );
  NOR2_X1 U774 ( .A1(n709), .A2(n708), .ZN(G54) );
  NOR2_X1 U775 ( .A1(n710), .A2(KEYINPUT2), .ZN(n711) );
  XNOR2_X1 U776 ( .A(n711), .B(KEYINPUT84), .ZN(n713) );
  NOR2_X1 U777 ( .A1(n659), .A2(KEYINPUT2), .ZN(n712) );
  NOR2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U779 ( .A(KEYINPUT82), .B(n714), .Z(n716) );
  OR2_X1 U780 ( .A1(n716), .A2(n715), .ZN(n759) );
  NOR2_X1 U781 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U782 ( .A(n719), .B(KEYINPUT115), .ZN(n720) );
  XNOR2_X1 U783 ( .A(n720), .B(KEYINPUT50), .ZN(n729) );
  XOR2_X1 U784 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n724) );
  NAND2_X1 U785 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U786 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U787 ( .A(n725), .B(KEYINPUT113), .ZN(n726) );
  NOR2_X1 U788 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U789 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U790 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U791 ( .A(KEYINPUT51), .B(n732), .Z(n734) );
  INV_X1 U792 ( .A(n733), .ZN(n753) );
  NAND2_X1 U793 ( .A1(n734), .A2(n753), .ZN(n735) );
  XNOR2_X1 U794 ( .A(n735), .B(KEYINPUT116), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n737), .B(KEYINPUT117), .ZN(n744) );
  INV_X1 U796 ( .A(n738), .ZN(n742) );
  NAND2_X1 U797 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U798 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U799 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U800 ( .A1(n745), .A2(n752), .ZN(n746) );
  NAND2_X1 U801 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U802 ( .A(KEYINPUT52), .B(n748), .Z(n751) );
  NAND2_X1 U803 ( .A1(G952), .A2(n749), .ZN(n750) );
  NOR2_X1 U804 ( .A1(n751), .A2(n750), .ZN(n757) );
  NAND2_X1 U805 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U806 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U807 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U808 ( .A1(n759), .A2(n758), .ZN(n761) );
  XOR2_X1 U809 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n760) );
  XNOR2_X1 U810 ( .A(n761), .B(n760), .ZN(G75) );
  NAND2_X1 U811 ( .A1(n763), .A2(n762), .ZN(n765) );
  XOR2_X1 U812 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n764) );
  XNOR2_X1 U813 ( .A(n765), .B(n764), .ZN(n766) );
  XNOR2_X1 U814 ( .A(G146), .B(n766), .ZN(G48) );
  XOR2_X1 U815 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n768) );
  XOR2_X1 U816 ( .A(n768), .B(n767), .Z(n769) );
  XNOR2_X1 U817 ( .A(n659), .B(n772), .ZN(n770) );
  NOR2_X1 U818 ( .A1(n770), .A2(G953), .ZN(n771) );
  XNOR2_X1 U819 ( .A(KEYINPUT125), .B(n771), .ZN(n777) );
  XNOR2_X1 U820 ( .A(G227), .B(n772), .ZN(n773) );
  NAND2_X1 U821 ( .A1(n773), .A2(G900), .ZN(n774) );
  NAND2_X1 U822 ( .A1(n774), .A2(G953), .ZN(n775) );
  XNOR2_X1 U823 ( .A(KEYINPUT126), .B(n775), .ZN(n776) );
  NAND2_X1 U824 ( .A1(n777), .A2(n776), .ZN(G72) );
endmodule

