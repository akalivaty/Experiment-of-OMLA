//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(G125), .A2(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  AOI211_X1 g008(.A(new_n188), .B(new_n190), .C1(new_n194), .C2(KEYINPUT16), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(KEYINPUT16), .ZN(new_n196));
  INV_X1    g010(.A(new_n190), .ZN(new_n197));
  AOI21_X1  g011(.A(G146), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(G237), .A2(G953), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G214), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT93), .A2(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n200), .B(G214), .C1(KEYINPUT93), .C2(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G131), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT17), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n203), .A2(new_n204), .A3(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n208), .B1(new_n203), .B2(new_n204), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT17), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n199), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G113), .B(G122), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n214), .B(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n194), .B(new_n188), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT18), .A2(G131), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n203), .A2(new_n204), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n217), .B(new_n219), .C1(new_n206), .C2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n213), .A2(new_n216), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n216), .B1(new_n213), .B2(new_n221), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n187), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(KEYINPUT94), .B(G475), .Z(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n196), .A2(G146), .A3(new_n197), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT19), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n194), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n192), .A2(KEYINPUT19), .A3(new_n193), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n188), .A3(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n203), .A2(new_n204), .A3(new_n208), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n229), .B(new_n233), .C1(new_n234), .C2(new_n211), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n221), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n216), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(G475), .B1(new_n222), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT20), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n239), .A2(new_n240), .A3(new_n187), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n239), .B2(new_n187), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n228), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT95), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT66), .A2(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT66), .A2(G128), .ZN(new_n246));
  OAI21_X1  g060(.A(G143), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT13), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n252), .A3(G134), .ZN(new_n253));
  XOR2_X1   g067(.A(G116), .B(G122), .Z(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G107), .ZN(new_n255));
  XNOR2_X1  g069(.A(G116), .B(G122), .ZN(new_n256));
  INV_X1    g070(.A(G107), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G134), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n247), .B(new_n249), .C1(new_n251), .C2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n253), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G116), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT14), .A3(G122), .ZN(new_n264));
  OAI211_X1 g078(.A(G107), .B(new_n264), .C1(new_n254), .C2(KEYINPUT14), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n247), .A2(new_n260), .A3(new_n249), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n260), .B1(new_n247), .B2(new_n249), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n265), .B(new_n258), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n244), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT9), .B(G234), .Z(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(G217), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n262), .A2(new_n268), .A3(new_n244), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n270), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n275), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n273), .B1(new_n277), .B2(new_n269), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(new_n278), .A3(new_n187), .ZN(new_n279));
  INV_X1    g093(.A(G478), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(KEYINPUT15), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n281), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n276), .A2(new_n278), .A3(new_n187), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n243), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(G234), .A2(G237), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(G952), .A3(new_n272), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT21), .B(G898), .Z(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(G902), .A3(G953), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n289), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n286), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT96), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n286), .A2(KEYINPUT96), .A3(new_n295), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n272), .A2(G227), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(new_n191), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT82), .ZN(new_n303));
  XOR2_X1   g117(.A(new_n303), .B(G110), .Z(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n248), .A2(G146), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n188), .A2(G143), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n307), .A2(new_n308), .A3(G128), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT64), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n248), .B2(G146), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n188), .A2(KEYINPUT64), .A3(G143), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT1), .B1(new_n248), .B2(G146), .ZN(new_n314));
  OR2_X1    g128(.A1(KEYINPUT66), .A2(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT66), .A2(G128), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n306), .A2(new_n309), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT10), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n257), .A3(G104), .ZN(new_n322));
  INV_X1    g136(.A(G101), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n215), .A2(G107), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n320), .A2(new_n322), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n257), .A2(G104), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n215), .A2(G107), .ZN(new_n327));
  OAI21_X1  g141(.A(G101), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n318), .A2(new_n319), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G101), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT83), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT4), .A4(new_n325), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n332), .A2(KEYINPUT4), .A3(new_n325), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT83), .B1(new_n332), .B2(KEYINPUT4), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(KEYINPUT0), .A2(G128), .ZN(new_n338));
  NOR2_X1   g152(.A1(KEYINPUT0), .A2(G128), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n313), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n307), .A2(new_n308), .A3(new_n338), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT65), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n307), .A2(new_n308), .A3(new_n338), .A4(KEYINPUT65), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n330), .B1(new_n337), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT11), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n260), .B2(G137), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n260), .A2(G137), .ZN(new_n350));
  INV_X1    g164(.A(G137), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT11), .A3(G134), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G131), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n349), .A2(new_n352), .A3(new_n208), .A4(new_n350), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n307), .A2(new_n308), .A3(new_n306), .A4(G128), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n314), .A2(G128), .B1(new_n307), .B2(new_n308), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n325), .B(new_n328), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n319), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n347), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n357), .B1(new_n347), .B2(new_n362), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n305), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT12), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n313), .A2(new_n317), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n329), .A2(new_n368), .A3(new_n358), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n361), .A3(KEYINPUT85), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n356), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT85), .B1(new_n369), .B2(new_n361), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n367), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT86), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(KEYINPUT86), .B(new_n367), .C1(new_n371), .C2(new_n372), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n369), .A2(new_n361), .ZN(new_n377));
  XOR2_X1   g191(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n378));
  NOR2_X1   g192(.A1(new_n357), .A2(new_n378), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n375), .A2(new_n376), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n363), .A2(new_n304), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n366), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G469), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n187), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n305), .B1(new_n380), .B2(new_n364), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n381), .A2(new_n365), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(G469), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(G469), .A2(G902), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n271), .ZN(new_n390));
  OAI21_X1  g204(.A(G221), .B1(new_n390), .B2(G902), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT81), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G214), .B1(G237), .B2(G902), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G210), .B1(G237), .B2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G119), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G116), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n263), .A2(G119), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT5), .ZN(new_n402));
  OAI21_X1  g216(.A(G113), .B1(new_n400), .B2(KEYINPUT5), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT87), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n400), .A2(new_n401), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT2), .B(G113), .Z(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n402), .B2(new_n403), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n405), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n329), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n406), .A2(KEYINPUT68), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(new_n407), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n412), .B1(new_n415), .B2(new_n337), .ZN(new_n416));
  XOR2_X1   g230(.A(G110), .B(G122), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  OR3_X1    g232(.A1(new_n416), .A2(KEYINPUT6), .A3(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n415), .A2(new_n337), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n417), .B1(new_n420), .B2(new_n412), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n415), .A2(new_n337), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n422), .B(new_n418), .C1(new_n329), .C2(new_n411), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT88), .B1(new_n346), .B2(new_n189), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n318), .A2(new_n189), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(G125), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n272), .A2(G224), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT89), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n430), .B(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n419), .A2(new_n424), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n430), .A2(new_n433), .ZN(new_n436));
  AOI22_X1  g250(.A1(KEYINPUT7), .A2(new_n436), .B1(new_n416), .B2(new_n418), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n411), .A2(new_n329), .ZN(new_n438));
  INV_X1    g252(.A(new_n404), .ZN(new_n439));
  INV_X1    g253(.A(new_n329), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n408), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT91), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT91), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n439), .A2(new_n440), .A3(new_n443), .A4(new_n408), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n438), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT90), .B(KEYINPUT8), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n417), .B(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT7), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n430), .B1(new_n449), .B2(new_n433), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(G902), .B1(new_n437), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n435), .B1(new_n452), .B2(KEYINPUT92), .ZN(new_n453));
  INV_X1    g267(.A(new_n430), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT7), .A3(new_n432), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n455), .A2(new_n423), .A3(new_n448), .A4(new_n450), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(KEYINPUT92), .A3(new_n187), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n398), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n187), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT92), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n462), .A2(new_n397), .A3(new_n457), .A4(new_n435), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n396), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n300), .A2(new_n394), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n194), .A2(new_n188), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT23), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n399), .B2(G128), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n399), .A2(G128), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n315), .A2(new_n316), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(G119), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n468), .B1(new_n471), .B2(new_n467), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G110), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT24), .B(G110), .Z(new_n474));
  NOR2_X1   g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n229), .B(new_n466), .C1(new_n473), .C2(new_n475), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n195), .A2(new_n198), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n472), .A2(G110), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(new_n474), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT78), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n471), .A2(KEYINPUT78), .A3(new_n474), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n477), .A2(new_n478), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT22), .B(G137), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT79), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n486));
  XOR2_X1   g300(.A(new_n485), .B(new_n486), .Z(new_n487));
  AND3_X1   g301(.A1(new_n476), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n476), .B2(new_n483), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n187), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT25), .ZN(new_n491));
  INV_X1    g305(.A(G217), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(G234), .B2(new_n187), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT25), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n494), .B(new_n187), .C1(new_n488), .C2(new_n489), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n493), .A2(G902), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n488), .B2(new_n489), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT80), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT80), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(new_n501), .A3(new_n498), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT77), .ZN(new_n504));
  INV_X1    g318(.A(G472), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT28), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n351), .A2(G134), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n260), .A2(G137), .ZN(new_n508));
  OAI21_X1  g322(.A(G131), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n355), .A2(new_n509), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n357), .A2(new_n427), .B1(new_n318), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n506), .B1(new_n415), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n346), .A2(new_n356), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT69), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n318), .A2(new_n515), .A3(new_n510), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n368), .A2(new_n358), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n355), .A2(new_n509), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT69), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n514), .B(new_n414), .C1(new_n516), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT70), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n515), .B1(new_n318), .B2(new_n510), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(KEYINPUT69), .A3(new_n518), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT70), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n514), .A4(new_n414), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT76), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n522), .A2(new_n523), .B1(new_n356), .B2(new_n346), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(new_n414), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n521), .A2(KEYINPUT76), .A3(new_n526), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n513), .B1(new_n534), .B2(KEYINPUT28), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(G101), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n200), .A2(G210), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT29), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(G902), .B1(new_n535), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n521), .A2(new_n526), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n346), .A2(new_n356), .B1(new_n517), .B2(new_n518), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(new_n414), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n544), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n548), .A2(KEYINPUT75), .A3(new_n512), .A4(new_n539), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n521), .B2(new_n526), .ZN(new_n550));
  INV_X1    g364(.A(new_n544), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n512), .B(new_n539), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT75), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n530), .A2(KEYINPUT30), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n546), .A2(KEYINPUT67), .A3(KEYINPUT30), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT67), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT30), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n511), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n555), .B(new_n415), .C1(new_n556), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n527), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n540), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n549), .A2(new_n554), .A3(new_n541), .A4(new_n562), .ZN(new_n563));
  AOI211_X1 g377(.A(new_n504), .B(new_n505), .C1(new_n543), .C2(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n521), .A2(KEYINPUT76), .A3(new_n526), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT76), .B1(new_n521), .B2(new_n526), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n565), .A2(new_n566), .A3(new_n531), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n512), .B(new_n542), .C1(new_n567), .C2(new_n506), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n554), .A2(new_n562), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n541), .B1(new_n552), .B2(new_n553), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n187), .B(new_n568), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT77), .B1(new_n571), .B2(G472), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT74), .ZN(new_n574));
  NOR2_X1   g388(.A1(G472), .A2(G902), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT67), .B1(new_n546), .B2(KEYINPUT30), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n511), .A2(new_n557), .A3(new_n558), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n577), .A2(new_n578), .B1(KEYINPUT30), .B2(new_n530), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n579), .A2(new_n415), .B1(new_n526), .B2(new_n521), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n580), .A2(KEYINPUT71), .A3(KEYINPUT31), .A4(new_n539), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n560), .A2(KEYINPUT71), .A3(new_n527), .A4(new_n539), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT31), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n512), .B1(new_n550), .B2(new_n551), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n540), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n576), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT73), .B(KEYINPUT32), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n574), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(KEYINPUT32), .ZN(new_n591));
  INV_X1    g405(.A(new_n589), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n581), .A2(new_n584), .B1(new_n540), .B2(new_n586), .ZN(new_n593));
  OAI211_X1 g407(.A(KEYINPUT74), .B(new_n592), .C1(new_n593), .C2(new_n576), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n465), .B(new_n503), .C1(new_n573), .C2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT97), .B(G101), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G3));
  NAND2_X1  g412(.A1(new_n276), .A2(new_n278), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT33), .B1(new_n276), .B2(new_n278), .ZN(new_n602));
  OAI211_X1 g416(.A(G478), .B(new_n187), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n279), .A2(new_n280), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n243), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n464), .A2(new_n295), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT98), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n464), .A2(new_n611), .A3(new_n295), .A4(new_n608), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n585), .A2(new_n587), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n187), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n588), .B1(new_n616), .B2(G472), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n503), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n389), .A2(new_n393), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  AND3_X1   g438(.A1(new_n419), .A2(new_n424), .A3(new_n434), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT92), .B1(new_n456), .B2(new_n187), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n397), .B1(new_n627), .B2(new_n457), .ZN(new_n628));
  INV_X1    g442(.A(new_n463), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n395), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n294), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n239), .A2(new_n240), .A3(new_n187), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n632), .B1(new_n242), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n239), .A2(KEYINPUT99), .A3(new_n240), .A4(new_n187), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n634), .A2(new_n635), .B1(new_n225), .B2(new_n227), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n636), .A2(new_n285), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n621), .A2(new_n631), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NAND2_X1  g454(.A1(new_n476), .A2(new_n483), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n487), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n497), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n496), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n465), .A2(new_n617), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT37), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G110), .ZN(G12));
  OR2_X1    g462(.A1(new_n292), .A2(G900), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n288), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n636), .A2(new_n285), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n636), .A2(KEYINPUT100), .A3(new_n285), .A4(new_n650), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n394), .A2(new_n464), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n655), .B(new_n645), .C1(new_n573), .C2(new_n595), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  OAI21_X1  g471(.A(new_n187), .B1(new_n534), .B2(new_n539), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n561), .A2(new_n539), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n590), .A2(new_n591), .A3(new_n594), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT101), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n650), .B(KEYINPUT39), .Z(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n394), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n663), .B1(KEYINPUT40), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n668));
  INV_X1    g482(.A(new_n645), .ZN(new_n669));
  INV_X1    g483(.A(new_n285), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n607), .A2(new_n670), .ZN(new_n671));
  AND4_X1   g485(.A1(new_n395), .A2(new_n668), .A3(new_n669), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n459), .A2(new_n463), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT38), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n667), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT102), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n248), .ZN(G45));
  NAND3_X1  g491(.A1(new_n605), .A2(new_n243), .A3(new_n650), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n630), .A2(new_n620), .A3(new_n678), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n679), .B(new_n645), .C1(new_n573), .C2(new_n595), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  NAND2_X1  g495(.A1(new_n571), .A2(G472), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n504), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n571), .A2(KEYINPUT77), .A3(G472), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n619), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n384), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n383), .B1(new_n382), .B2(new_n187), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n688), .A2(new_n689), .A3(new_n392), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n614), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT41), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G113), .ZN(G15));
  AOI21_X1  g507(.A(new_n294), .B1(new_n500), .B2(new_n502), .ZN(new_n694));
  AND4_X1   g508(.A1(new_n464), .A2(new_n690), .A3(new_n694), .A4(new_n637), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n695), .B1(new_n573), .B2(new_n595), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  AND3_X1   g511(.A1(new_n300), .A2(new_n464), .A3(new_n690), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n698), .B(new_n645), .C1(new_n573), .C2(new_n595), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  XNOR2_X1  g514(.A(KEYINPUT104), .B(G472), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n616), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n499), .B(KEYINPUT105), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n585), .B1(new_n535), .B2(new_n539), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n575), .B(KEYINPUT103), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n690), .A2(new_n702), .A3(new_n703), .A4(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n631), .A3(new_n671), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  INV_X1    g523(.A(new_n678), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n702), .A2(new_n710), .A3(new_n645), .A4(new_n706), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n464), .A2(new_n690), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n189), .ZN(G27));
  INV_X1    g528(.A(KEYINPUT32), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n593), .B2(new_n576), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n593), .A2(new_n715), .A3(new_n576), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n716), .B1(new_n717), .B2(KEYINPUT108), .ZN(new_n718));
  OR3_X1    g532(.A1(new_n588), .A2(KEYINPUT108), .A3(KEYINPUT32), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n718), .B(new_n719), .C1(new_n564), .C2(new_n572), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n720), .A2(KEYINPUT42), .A3(new_n703), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n387), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n385), .A2(KEYINPUT106), .A3(G469), .A4(new_n386), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(new_n384), .A3(new_n388), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(KEYINPUT107), .A3(new_n393), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT107), .B1(new_n725), .B2(new_n393), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n459), .A2(new_n395), .A3(new_n463), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n727), .A2(new_n728), .A3(new_n678), .A4(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n721), .A2(KEYINPUT109), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n720), .A2(KEYINPUT42), .A3(new_n703), .ZN(new_n733));
  INV_X1    g547(.A(new_n728), .ZN(new_n734));
  INV_X1    g548(.A(new_n729), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n710), .A3(new_n726), .A4(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n732), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n687), .A2(new_n739), .A3(new_n710), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n731), .A2(new_n737), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n208), .ZN(G33));
  NAND4_X1  g556(.A1(new_n687), .A2(new_n739), .A3(new_n653), .A4(new_n654), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  NAND2_X1  g558(.A1(new_n385), .A2(new_n386), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(G469), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT46), .B1(new_n747), .B2(new_n388), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n688), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n388), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n392), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(new_n665), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n243), .B(KEYINPUT111), .Z(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n605), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n606), .A2(new_n243), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n754), .B(KEYINPUT43), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n756), .B2(KEYINPUT110), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n618), .A3(new_n645), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n729), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n752), .B(new_n762), .C1(new_n761), .C2(new_n760), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  XNOR2_X1  g578(.A(new_n751), .B(KEYINPUT47), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n503), .A2(new_n678), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n685), .A2(new_n686), .A3(new_n735), .A4(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT112), .Z(new_n768));
  AOI21_X1  g582(.A(KEYINPUT113), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n765), .A2(KEYINPUT113), .A3(new_n768), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  AND3_X1   g587(.A1(new_n757), .A2(new_n289), .A3(new_n759), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n674), .A2(new_n395), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n707), .A3(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n776), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT50), .B1(new_n776), .B2(KEYINPUT116), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n702), .A2(new_n706), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n774), .A2(new_n703), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n688), .A2(new_n689), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n393), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n735), .B(new_n781), .C1(new_n765), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n690), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n729), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n663), .A2(new_n503), .A3(new_n289), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n606), .A2(new_n607), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n774), .A2(new_n787), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n780), .A2(new_n645), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(KEYINPUT118), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n790), .B2(new_n794), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n779), .B(new_n785), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT51), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n801));
  INV_X1    g615(.A(new_n779), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(new_n802), .B2(new_n795), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n779), .A2(KEYINPUT117), .A3(new_n794), .A4(new_n790), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n785), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n800), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n740), .A2(new_n738), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT109), .B1(new_n721), .B2(new_n730), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n733), .A2(new_n736), .A3(new_n732), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n503), .B1(new_n573), .B2(new_n595), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n813), .A2(new_n613), .A3(new_n786), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n617), .A2(new_n503), .ZN(new_n815));
  INV_X1    g629(.A(new_n608), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n670), .B2(new_n243), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n394), .A3(new_n631), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n596), .A2(new_n818), .A3(new_n646), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n699), .A2(new_n708), .A3(new_n696), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n814), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n730), .A2(new_n793), .ZN(new_n822));
  INV_X1    g636(.A(new_n650), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n285), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n735), .A2(KEYINPUT115), .A3(new_n636), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n459), .A2(new_n395), .A3(new_n463), .A4(new_n636), .ZN(new_n827));
  INV_X1    g641(.A(new_n824), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n620), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n669), .B1(new_n685), .B2(new_n686), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n743), .A2(new_n822), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n812), .A2(new_n821), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n713), .B1(new_n831), .B2(new_n655), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n464), .A2(new_n671), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n725), .A2(new_n393), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n645), .A2(new_n823), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n837), .A2(new_n662), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n835), .A2(new_n836), .A3(new_n680), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n713), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n656), .A2(new_n680), .A3(new_n843), .A4(new_n841), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n808), .B1(new_n834), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n596), .A2(new_n646), .A3(new_n818), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n699), .A2(new_n696), .A3(new_n708), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n691), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n743), .A2(new_n822), .A3(new_n832), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n842), .A2(new_n845), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n853), .A3(KEYINPUT53), .A4(new_n812), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n847), .A2(KEYINPUT54), .A3(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n807), .B(new_n859), .C1(new_n816), .C2(new_n788), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n720), .A2(new_n703), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n791), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT48), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n781), .A2(new_n464), .A3(new_n690), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(G952), .A3(new_n272), .A4(new_n864), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n860), .A2(new_n865), .B1(G952), .B2(G953), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n703), .B1(new_n783), .B2(KEYINPUT49), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n674), .A2(new_n396), .A3(new_n867), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n392), .B(new_n754), .C1(KEYINPUT49), .C2(new_n783), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n663), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT114), .Z(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n871), .ZN(G75));
  NOR2_X1   g686(.A1(new_n272), .A2(G952), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n187), .B1(new_n847), .B2(new_n854), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT56), .B1(new_n875), .B2(G210), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n419), .A2(new_n424), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n434), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n882), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n878), .B1(new_n883), .B2(new_n884), .ZN(G51));
  XNOR2_X1  g699(.A(new_n388), .B(KEYINPUT57), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n382), .B1(new_n859), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n875), .A2(G469), .A3(new_n746), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n873), .B1(new_n887), .B2(new_n888), .ZN(G54));
  NAND3_X1  g703(.A1(new_n875), .A2(KEYINPUT58), .A3(G475), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n222), .A2(new_n238), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n890), .A2(new_n892), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n893), .A2(new_n894), .A3(new_n873), .ZN(G60));
  NAND2_X1  g709(.A1(G478), .A2(G902), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT59), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n857), .A2(new_n858), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n601), .A2(new_n602), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n900), .A2(new_n901), .A3(new_n873), .ZN(G63));
  XNOR2_X1  g716(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n492), .A2(new_n187), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n741), .A2(new_n850), .A3(new_n851), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT53), .B1(new_n906), .B2(new_n853), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n814), .A2(new_n820), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n833), .A2(new_n908), .A3(new_n848), .ZN(new_n909));
  NOR4_X1   g723(.A1(new_n909), .A2(new_n846), .A3(new_n741), .A4(new_n808), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n905), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n488), .A2(new_n489), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n873), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n914));
  AND4_X1   g728(.A1(new_n914), .A2(new_n855), .A3(new_n643), .A4(new_n905), .ZN(new_n915));
  INV_X1    g729(.A(new_n905), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n847), .B2(new_n854), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n917), .B2(new_n643), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n913), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT61), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n855), .A2(new_n643), .A3(new_n905), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT121), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n917), .A2(new_n914), .A3(new_n643), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n920), .A2(KEYINPUT61), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n920), .A2(KEYINPUT61), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .A4(new_n913), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n921), .A2(new_n928), .ZN(G66));
  INV_X1    g743(.A(G224), .ZN(new_n930));
  OAI21_X1  g744(.A(G953), .B1(new_n291), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n821), .B2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n880), .B1(G898), .B2(new_n272), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(G69));
  NAND2_X1  g748(.A1(new_n231), .A2(new_n232), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n579), .B(new_n935), .Z(new_n936));
  NAND3_X1  g750(.A1(new_n752), .A2(new_n861), .A3(new_n837), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n771), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n743), .B(new_n939), .C1(new_n940), .C2(new_n769), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n937), .A2(new_n938), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n656), .A2(new_n680), .A3(new_n843), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n942), .A2(new_n812), .A3(new_n763), .A4(new_n945), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n941), .A2(new_n946), .A3(G953), .ZN(new_n947));
  INV_X1    g761(.A(G227), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n272), .B1(new_n948), .B2(G900), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n936), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n945), .A2(new_n675), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT124), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(KEYINPUT62), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n951), .B(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n687), .A2(new_n394), .A3(new_n665), .A4(new_n817), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n763), .B1(new_n729), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n763), .B(new_n958), .C1(new_n729), .C2(new_n955), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI22_X1  g774(.A1(new_n770), .A2(new_n771), .B1(new_n952), .B2(KEYINPUT62), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n954), .A2(new_n960), .A3(new_n961), .A4(new_n272), .ZN(new_n962));
  INV_X1    g776(.A(new_n936), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n949), .A2(G900), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n950), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n950), .B2(new_n965), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(G72));
  NOR3_X1   g783(.A1(new_n941), .A2(new_n946), .A3(new_n850), .ZN(new_n970));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n540), .B(new_n580), .C1(new_n970), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n580), .A2(new_n539), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n562), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n855), .A2(new_n972), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n974), .A2(new_n874), .A3(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n954), .A2(new_n960), .A3(new_n961), .A4(new_n821), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n659), .B1(new_n979), .B2(new_n972), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n978), .A2(new_n980), .ZN(G57));
endmodule


