//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G116), .ZN(new_n192));
  OAI21_X1  g006(.A(G113), .B1(new_n192), .B2(KEYINPUT5), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n191), .A2(G116), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n194), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G119), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n192), .A2(new_n199), .A3(KEYINPUT65), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n193), .B1(new_n201), .B2(KEYINPUT5), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT79), .B1(new_n203), .B2(G107), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT79), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G101), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n206), .A3(G104), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n211), .A2(new_n213), .A3(new_n214), .A4(new_n208), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n217));
  AND3_X1   g031(.A1(KEYINPUT64), .A2(KEYINPUT2), .A3(G113), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT64), .B1(KEYINPUT2), .B2(G113), .ZN(new_n219));
  OAI22_X1  g033(.A1(new_n218), .A2(new_n219), .B1(KEYINPUT2), .B2(G113), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n192), .A2(new_n199), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR4_X1   g036(.A1(new_n202), .A2(new_n216), .A3(new_n217), .A4(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n192), .A2(new_n199), .A3(KEYINPUT65), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT65), .B1(new_n192), .B2(new_n199), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT5), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n193), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n222), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n216), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT82), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n220), .A2(new_n221), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n198), .A2(new_n220), .A3(new_n200), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n211), .A2(new_n213), .A3(new_n208), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT77), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT77), .A4(new_n208), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n237), .A2(new_n238), .A3(G101), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(G101), .A3(new_n239), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n215), .A2(KEYINPUT4), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT78), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n242), .A2(KEYINPUT78), .A3(new_n243), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n241), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n190), .B1(new_n231), .B2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n234), .A2(new_n240), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n242), .A2(KEYINPUT78), .A3(new_n243), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT78), .B1(new_n242), .B2(new_n243), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT5), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n198), .B2(new_n200), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n232), .B1(new_n255), .B2(new_n193), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n217), .B1(new_n256), .B2(new_n216), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n228), .A2(KEYINPUT82), .A3(new_n229), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n253), .A2(new_n259), .A3(new_n189), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n249), .A2(KEYINPUT6), .A3(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G143), .B(G146), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(G128), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  INV_X1    g079(.A(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G143), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n265), .B1(new_n267), .B2(KEYINPUT1), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n264), .B1(new_n268), .B2(new_n262), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G125), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G146), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT0), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(new_n265), .ZN(new_n277));
  NOR2_X1   g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n262), .B1(new_n276), .B2(new_n265), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(G125), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G224), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n282), .B(new_n284), .Z(new_n285));
  NAND2_X1  g099(.A1(new_n253), .A2(new_n259), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n189), .A2(KEYINPUT6), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT83), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT83), .ZN(new_n289));
  INV_X1    g103(.A(new_n287), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n289), .B(new_n290), .C1(new_n253), .C2(new_n259), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n261), .B(new_n285), .C1(new_n288), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT84), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n286), .A2(new_n287), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n289), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n286), .A2(KEYINPUT83), .A3(new_n287), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n298), .A2(KEYINPUT84), .A3(new_n261), .A4(new_n285), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n282), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n281), .A2(KEYINPUT85), .B1(KEYINPUT7), .B2(new_n284), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n228), .A2(new_n216), .ZN(new_n305));
  XOR2_X1   g119(.A(new_n189), .B(KEYINPUT8), .Z(new_n306));
  OAI21_X1  g120(.A(new_n227), .B1(new_n254), .B2(new_n221), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n232), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n306), .B1(new_n308), .B2(new_n229), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n303), .A2(new_n304), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(G902), .B1(new_n310), .B2(new_n260), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n300), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G210), .B1(G237), .B2(G902), .ZN(new_n313));
  XOR2_X1   g127(.A(new_n313), .B(KEYINPUT86), .Z(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n300), .A2(new_n313), .A3(new_n311), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n188), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT11), .ZN(new_n318));
  INV_X1    g132(.A(G134), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(G137), .ZN(new_n320));
  INV_X1    g134(.A(G137), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT11), .A3(G134), .ZN(new_n322));
  INV_X1    g136(.A(G131), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(G137), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n320), .A2(new_n322), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n319), .A2(G137), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n321), .A2(G134), .ZN(new_n327));
  OAI21_X1  g141(.A(G131), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n270), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G131), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n325), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n279), .A2(new_n280), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n330), .A2(new_n336), .A3(KEYINPUT30), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n329), .A2(KEYINPUT66), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT66), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n325), .A2(new_n328), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n341), .A3(new_n269), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n338), .B1(new_n342), .B2(new_n335), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n234), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(G237), .A2(G953), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G210), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT27), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT26), .B(G101), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n234), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n342), .A2(new_n350), .A3(new_n335), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n344), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT31), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT31), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n344), .A2(new_n354), .A3(new_n349), .A4(new_n351), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n234), .B1(new_n330), .B2(new_n336), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n351), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT28), .ZN(new_n358));
  INV_X1    g172(.A(new_n351), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT67), .B1(new_n359), .B2(KEYINPUT28), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT67), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n351), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n358), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n353), .B(new_n355), .C1(new_n364), .C2(new_n349), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT32), .ZN(new_n366));
  NOR2_X1   g180(.A1(G472), .A2(G902), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n365), .B2(new_n367), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n360), .A2(new_n363), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n350), .B1(new_n342), .B2(new_n335), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n351), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT68), .A3(KEYINPUT28), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT28), .B1(new_n359), .B2(new_n372), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT68), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n371), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT29), .A3(new_n349), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n344), .A2(new_n351), .ZN(new_n381));
  INV_X1    g195(.A(new_n349), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n358), .A2(new_n360), .A3(new_n349), .A4(new_n363), .ZN(new_n384));
  AOI21_X1  g198(.A(G902), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G472), .ZN(new_n387));
  OAI22_X1  g201(.A1(new_n369), .A2(new_n370), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n265), .A2(KEYINPUT23), .A3(G119), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n191), .A2(G128), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n191), .A2(G128), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n389), .B(new_n390), .C1(new_n391), .C2(KEYINPUT23), .ZN(new_n392));
  XOR2_X1   g206(.A(KEYINPUT24), .B(G110), .Z(new_n393));
  XNOR2_X1  g207(.A(G119), .B(G128), .ZN(new_n394));
  OAI22_X1  g208(.A1(new_n392), .A2(G110), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G125), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n271), .A2(G140), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT16), .ZN(new_n399));
  OR3_X1    g213(.A1(new_n271), .A2(KEYINPUT16), .A3(G140), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(G146), .ZN(new_n401));
  XNOR2_X1  g215(.A(G125), .B(G140), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n266), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n395), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n392), .A2(G110), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n265), .A2(G119), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n390), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT24), .B(G110), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT69), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT69), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n393), .B2(new_n394), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n406), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n399), .A2(G146), .A3(new_n400), .ZN(new_n414));
  AOI21_X1  g228(.A(G146), .B1(new_n399), .B2(new_n400), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT70), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n393), .A2(new_n394), .A3(new_n411), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT69), .B1(new_n408), .B2(new_n409), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n418), .A2(new_n419), .B1(G110), .B2(new_n392), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n399), .A2(new_n400), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n266), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n401), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT70), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n405), .B1(new_n417), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT22), .B(G137), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT71), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n420), .A2(new_n423), .A3(new_n424), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n424), .B1(new_n420), .B2(new_n423), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n404), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT71), .ZN(new_n434));
  INV_X1    g248(.A(new_n429), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n404), .B(new_n429), .C1(new_n431), .C2(new_n432), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT72), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n426), .A2(KEYINPUT72), .A3(new_n429), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n430), .A2(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G217), .ZN(new_n442));
  INV_X1    g256(.A(G902), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(G234), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(G902), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n430), .A2(new_n436), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n439), .A2(new_n440), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n443), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT25), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT73), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT25), .A4(new_n443), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT74), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n441), .A2(KEYINPUT74), .A3(KEYINPUT25), .A4(new_n443), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT73), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n449), .A2(new_n457), .A3(new_n450), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n452), .A2(new_n455), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n446), .B1(new_n459), .B2(new_n444), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT9), .B(G234), .ZN(new_n461));
  OAI21_X1  g275(.A(G221), .B1(new_n461), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(G469), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n283), .A2(G227), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT75), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G140), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT10), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n270), .A2(new_n216), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT81), .ZN(new_n470));
  AND4_X1   g284(.A1(new_n263), .A2(new_n267), .A3(new_n274), .A4(G128), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT1), .B1(new_n273), .B2(G146), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT80), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n267), .A2(KEYINPUT80), .A3(KEYINPUT1), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(G128), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n471), .B1(new_n476), .B2(new_n275), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(new_n216), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n470), .B1(new_n478), .B2(KEYINPUT10), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT81), .B(new_n468), .C1(new_n477), .C2(new_n216), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n469), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n334), .B(new_n240), .C1(new_n251), .C2(new_n252), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n333), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n480), .ZN(new_n485));
  INV_X1    g299(.A(new_n333), .ZN(new_n486));
  INV_X1    g300(.A(new_n469), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n482), .A4(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n467), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n229), .A2(new_n269), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n333), .B1(new_n490), .B2(new_n478), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT12), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(KEYINPUT12), .B(new_n333), .C1(new_n490), .C2(new_n478), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n488), .A2(new_n495), .A3(new_n467), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n463), .B(new_n443), .C1(new_n489), .C2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n488), .A2(new_n495), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n467), .B(KEYINPUT76), .Z(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n486), .B1(new_n481), .B2(new_n482), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n488), .A2(new_n467), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n463), .B1(new_n504), .B2(new_n443), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n462), .B1(new_n498), .B2(new_n505), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n461), .A2(new_n442), .A3(G953), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT91), .B1(new_n195), .B2(G122), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n510));
  INV_X1    g324(.A(G122), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(G116), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n195), .A2(G122), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n513), .A2(KEYINPUT92), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT92), .B1(new_n513), .B2(new_n514), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n206), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n514), .A2(KEYINPUT14), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n514), .A2(KEYINPUT14), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n273), .A2(G128), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n273), .A2(G128), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n319), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n523), .ZN(new_n525));
  OAI21_X1  g339(.A(G134), .B1(new_n525), .B2(new_n521), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n520), .A2(G107), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n508), .B1(new_n517), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n517), .A2(new_n508), .A3(new_n527), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT13), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n523), .A2(KEYINPUT93), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT93), .B1(new_n523), .B2(new_n532), .ZN(new_n535));
  OAI221_X1 g349(.A(new_n522), .B1(new_n532), .B2(new_n523), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G134), .ZN(new_n537));
  INV_X1    g351(.A(new_n516), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n513), .A2(KEYINPUT92), .A3(new_n514), .ZN(new_n539));
  AOI21_X1  g353(.A(G107), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n515), .A2(new_n516), .A3(new_n206), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n524), .B(new_n537), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n507), .B1(new_n531), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n530), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n542), .B(new_n507), .C1(new_n544), .C2(new_n528), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n443), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G478), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(KEYINPUT15), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  OAI221_X1 g364(.A(new_n443), .B1(KEYINPUT15), .B2(new_n548), .C1(new_n546), .C2(new_n543), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G952), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(G953), .ZN(new_n555));
  NAND2_X1  g369(.A1(G234), .A2(G237), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT21), .B(G898), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(G902), .A3(G953), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G237), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n283), .A3(G214), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(KEYINPUT87), .A3(new_n273), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n273), .A2(KEYINPUT87), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(G214), .A3(new_n345), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(KEYINPUT18), .A3(G131), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n397), .A2(new_n398), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G146), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n403), .ZN(new_n571));
  NAND2_X1  g385(.A1(KEYINPUT18), .A2(G131), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n564), .A2(new_n572), .A3(new_n566), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n568), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n567), .A2(G131), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n323), .B1(new_n564), .B2(new_n566), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n575), .A2(KEYINPUT17), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(KEYINPUT17), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n416), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n574), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g394(.A(G113), .B(G122), .Z(new_n581));
  XOR2_X1   g395(.A(KEYINPUT88), .B(G104), .Z(new_n582));
  XOR2_X1   g396(.A(new_n581), .B(new_n582), .Z(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n583), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n585), .B(new_n574), .C1(new_n577), .C2(new_n579), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n443), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(G475), .ZN(new_n589));
  NOR2_X1   g403(.A1(G475), .A2(G902), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n402), .A2(KEYINPUT19), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n402), .A2(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n266), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n593), .B(new_n401), .C1(new_n575), .C2(new_n576), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n574), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n583), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT89), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n596), .A2(new_n597), .A3(new_n586), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n596), .B2(new_n586), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n590), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT20), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(new_n586), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT20), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n590), .A2(KEYINPUT90), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n590), .A2(KEYINPUT90), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n602), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n589), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n553), .A2(new_n561), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n506), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n317), .A2(new_n388), .A3(new_n460), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  NAND2_X1  g425(.A1(new_n365), .A2(new_n443), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G472), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n365), .A2(new_n367), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n506), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n616), .A2(new_n460), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n300), .A2(KEYINPUT95), .A3(new_n313), .A4(new_n311), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n187), .ZN(new_n619));
  INV_X1    g433(.A(new_n313), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n312), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n311), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n294), .B2(new_n299), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT95), .B1(new_n623), .B2(new_n313), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n619), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n547), .A2(new_n548), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n543), .A2(KEYINPUT97), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n542), .B1(new_n544), .B2(new_n528), .ZN(new_n628));
  INV_X1    g442(.A(new_n507), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n627), .A2(new_n632), .A3(KEYINPUT33), .A4(new_n545), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT96), .B(KEYINPUT33), .Z(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(new_n543), .B2(new_n546), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n443), .A2(G478), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n626), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n601), .A2(new_n606), .ZN(new_n639));
  INV_X1    g453(.A(new_n589), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n561), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n617), .A2(new_n625), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  OAI211_X1 g461(.A(new_n603), .B(new_n590), .C1(new_n598), .C2(new_n599), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n589), .B1(new_n601), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(new_n561), .A3(new_n552), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT98), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n617), .A2(new_n625), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT99), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n435), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n426), .B(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n657), .A2(G902), .A3(new_n444), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n459), .B2(new_n444), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n608), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n317), .A3(new_n616), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  NAND2_X1  g477(.A1(new_n459), .A2(new_n444), .ZN(new_n664));
  INV_X1    g478(.A(new_n658), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n462), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n503), .A2(new_n502), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n499), .B2(new_n500), .ZN(new_n669));
  OAI21_X1  g483(.A(G469), .B1(new_n669), .B2(G902), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n667), .B1(new_n670), .B2(new_n497), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n666), .A2(new_n388), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n621), .A2(new_n624), .ZN(new_n673));
  AOI211_X1 g487(.A(new_n620), .B(new_n622), .C1(new_n294), .C2(new_n299), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n188), .B1(new_n674), .B2(KEYINPUT95), .ZN(new_n675));
  INV_X1    g489(.A(new_n649), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n283), .A2(G900), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(G902), .A3(new_n556), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n680), .A2(new_n557), .A3(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n676), .A2(new_n553), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n673), .A2(new_n675), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n673), .A2(new_n675), .A3(KEYINPUT101), .A4(new_n683), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n672), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n265), .ZN(G30));
  XNOR2_X1  g503(.A(new_n682), .B(KEYINPUT39), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n506), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT104), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT40), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n691), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n674), .B1(new_n314), .B2(new_n312), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n374), .A2(new_n382), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT103), .Z(new_n702));
  AOI21_X1  g516(.A(G902), .B1(new_n702), .B2(new_n352), .ZN(new_n703));
  OAI22_X1  g517(.A1(new_n369), .A2(new_n370), .B1(new_n703), .B2(new_n387), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n553), .A2(new_n607), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n659), .A3(new_n187), .A4(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n694), .A2(new_n697), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT105), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n694), .A2(new_n697), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n273), .ZN(G45));
  INV_X1    g527(.A(new_n682), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n638), .A2(new_n641), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n666), .A2(new_n388), .A3(new_n671), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n673), .A2(new_n675), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT106), .B(G146), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G48));
  NAND3_X1  g534(.A1(new_n673), .A2(new_n675), .A3(new_n644), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n443), .B1(new_n489), .B2(new_n496), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(G469), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n462), .A3(new_n497), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT107), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n723), .A2(new_n726), .A3(new_n462), .A4(new_n497), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n725), .A2(new_n388), .A3(new_n460), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT41), .B(G113), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND3_X1  g545(.A1(new_n651), .A2(new_n673), .A3(new_n675), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n728), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n195), .ZN(G18));
  NAND4_X1  g548(.A1(new_n673), .A2(new_n675), .A3(new_n727), .A4(new_n725), .ZN(new_n735));
  INV_X1    g549(.A(new_n608), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n666), .A2(new_n388), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n191), .ZN(G21));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n740));
  INV_X1    g554(.A(new_n444), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n449), .A2(new_n457), .A3(new_n450), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n457), .B1(new_n449), .B2(new_n450), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n455), .A2(new_n456), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT109), .B1(new_n746), .B2(new_n446), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n748));
  INV_X1    g562(.A(new_n446), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n664), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n725), .A2(new_n561), .A3(new_n727), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n353), .B1(new_n379), .B2(new_n349), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT108), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(new_n353), .C1(new_n379), .C2(new_n349), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n355), .A3(new_n756), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n757), .A2(new_n367), .B1(G472), .B2(new_n612), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n751), .A2(new_n752), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n625), .A2(new_n705), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n740), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n758), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n747), .B2(new_n750), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n673), .A2(new_n675), .A3(new_n705), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(new_n764), .A3(KEYINPUT110), .A4(new_n752), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT111), .B(G122), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G24));
  NAND3_X1  g582(.A1(new_n758), .A2(new_n666), .A3(new_n715), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n735), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n271), .ZN(G27));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  INV_X1    g586(.A(new_n388), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n747), .B2(new_n750), .ZN(new_n774));
  INV_X1    g588(.A(new_n314), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n316), .B(new_n187), .C1(new_n775), .C2(new_n623), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n638), .A2(new_n641), .A3(new_n714), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n776), .A2(new_n506), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n772), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n388), .A2(new_n460), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n715), .A2(new_n772), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n780), .A2(new_n781), .A3(new_n776), .A4(new_n506), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  INV_X1    g598(.A(new_n683), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n780), .A2(new_n776), .A3(new_n785), .A4(new_n506), .ZN(new_n786));
  XOR2_X1   g600(.A(KEYINPUT112), .B(G134), .Z(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(G36));
  NAND2_X1  g602(.A1(new_n638), .A2(new_n607), .ZN(new_n789));
  AND2_X1   g603(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n790));
  NOR2_X1   g604(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n789), .B2(new_n791), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n615), .A3(new_n666), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n776), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n463), .B1(new_n504), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n797), .B2(new_n504), .ZN(new_n799));
  NAND2_X1  g613(.A1(G469), .A2(G902), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT46), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n498), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n800), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n667), .B(new_n690), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n796), .B(new_n804), .C1(new_n795), .C2(new_n794), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  AOI21_X1  g620(.A(new_n667), .B1(new_n802), .B2(new_n803), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT47), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n776), .A2(new_n388), .A3(new_n460), .A4(new_n777), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  NAND2_X1  g625(.A1(new_n723), .A2(new_n497), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n812), .A2(KEYINPUT49), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(KEYINPUT49), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n638), .A2(new_n187), .A3(new_n607), .A4(new_n462), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n813), .A2(new_n814), .A3(new_n704), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n700), .A2(new_n751), .A3(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n725), .A2(new_n727), .ZN(new_n818));
  INV_X1    g632(.A(new_n776), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n460), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n820), .A2(new_n821), .A3(new_n557), .A4(new_n704), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n823), .A2(new_n641), .A3(new_n638), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n793), .A2(new_n556), .A3(new_n555), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n818), .A3(new_n819), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT118), .Z(new_n827));
  NOR2_X1   g641(.A1(new_n762), .A2(new_n659), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n825), .A2(new_n763), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n776), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n812), .A2(new_n462), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n831), .B1(new_n808), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n700), .A2(new_n188), .A3(new_n818), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT117), .B1(new_n834), .B2(new_n830), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT50), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n829), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  OAI221_X1 g654(.A(new_n555), .B1(new_n735), .B2(new_n830), .C1(new_n823), .C2(new_n642), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n827), .A2(new_n774), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT48), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(KEYINPUT48), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n839), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n847));
  INV_X1    g661(.A(new_n672), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT101), .B1(new_n625), .B2(new_n683), .ZN(new_n849));
  INV_X1    g663(.A(new_n687), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n735), .A2(new_n769), .B1(new_n716), .B2(new_n717), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n682), .B(KEYINPUT115), .Z(new_n854));
  NAND3_X1  g668(.A1(new_n659), .A2(new_n671), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n659), .A2(new_n671), .A3(KEYINPUT116), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n704), .A3(new_n764), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n851), .A2(new_n853), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n686), .A2(new_n687), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n852), .B1(new_n864), .B2(new_n848), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(KEYINPUT52), .A3(new_n860), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n641), .B(new_n626), .C1(new_n636), .C2(new_n637), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n553), .A2(new_n607), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n868), .A2(new_n869), .A3(new_n561), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n317), .A2(new_n870), .A3(new_n460), .A4(new_n616), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n610), .A3(new_n661), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n728), .B1(new_n732), .B2(new_n721), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n872), .A2(new_n873), .A3(new_n738), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n779), .A2(new_n782), .A3(new_n786), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n676), .A2(new_n552), .A3(new_n682), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n819), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT114), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n672), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n819), .A2(KEYINPUT114), .A3(new_n876), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n879), .A2(new_n880), .B1(new_n828), .B2(new_n778), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n766), .A2(new_n874), .A3(new_n875), .A4(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n867), .A2(KEYINPUT53), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n867), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n847), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT52), .B1(new_n865), .B2(new_n860), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n673), .A2(new_n675), .A3(new_n704), .A4(new_n705), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n857), .B2(new_n858), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n688), .A2(new_n889), .A3(new_n852), .A4(new_n862), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n766), .A2(new_n874), .A3(new_n875), .A4(new_n881), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n867), .A2(new_n882), .A3(KEYINPUT53), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(KEYINPUT54), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n846), .B1(new_n885), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n554), .A2(new_n283), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT119), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n817), .B1(new_n896), .B2(new_n898), .ZN(G75));
  NOR2_X1   g713(.A1(new_n283), .A2(G952), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n443), .B1(new_n893), .B2(new_n894), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n902), .A2(new_n314), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n298), .A2(new_n261), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n285), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT55), .Z(new_n906));
  OR2_X1    g720(.A1(new_n906), .A2(KEYINPUT56), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n901), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n902), .A2(G210), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n906), .B1(new_n909), .B2(KEYINPUT56), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(KEYINPUT120), .B(new_n906), .C1(new_n909), .C2(KEYINPUT56), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(G51));
  NOR2_X1   g728(.A1(new_n489), .A2(new_n496), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n800), .B(KEYINPUT57), .Z(new_n916));
  NAND3_X1  g730(.A1(new_n885), .A2(new_n895), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n918), .B2(new_n917), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n902), .B(new_n798), .C1(new_n797), .C2(new_n504), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n900), .B1(new_n920), .B2(new_n921), .ZN(G54));
  NAND3_X1  g736(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n598), .A2(new_n599), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n900), .ZN(G60));
  INV_X1    g741(.A(new_n636), .ZN(new_n928));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT59), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n885), .A2(new_n928), .A3(new_n895), .A4(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n931), .A2(KEYINPUT122), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(KEYINPUT122), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n901), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n885), .A2(new_n895), .A3(new_n930), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n935), .A2(new_n936), .A3(new_n636), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n935), .B2(new_n636), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n934), .A2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(new_n893), .A2(new_n894), .ZN(new_n941));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT60), .Z(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n944), .A2(new_n657), .ZN(new_n945));
  INV_X1    g759(.A(new_n441), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n901), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n945), .A2(KEYINPUT61), .A3(new_n901), .A4(new_n947), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(G66));
  AOI21_X1  g766(.A(new_n283), .B1(new_n559), .B2(G224), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n766), .A2(new_n874), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n953), .B1(new_n955), .B2(new_n283), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n904), .B1(G898), .B2(new_n283), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(new_n957), .Z(G69));
  XOR2_X1   g772(.A(new_n875), .B(KEYINPUT126), .Z(new_n959));
  NAND3_X1  g773(.A1(new_n804), .A2(new_n764), .A3(new_n774), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n810), .A2(new_n805), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n961), .A3(new_n865), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n677), .B1(new_n962), .B2(new_n283), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n337), .A2(new_n343), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n591), .A2(new_n592), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n966), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n709), .A2(new_n711), .A3(new_n865), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n970));
  AND4_X1   g784(.A1(new_n388), .A2(new_n460), .A3(new_n869), .A4(new_n868), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n692), .A2(new_n819), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n805), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n805), .A2(KEYINPUT124), .A3(new_n972), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n709), .A2(new_n711), .A3(new_n978), .A4(new_n865), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n970), .A2(new_n810), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n968), .B1(new_n980), .B2(new_n283), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n967), .A2(new_n981), .A3(KEYINPUT125), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n283), .B1(G227), .B2(G900), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n980), .B2(new_n955), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n349), .A3(new_n381), .ZN(new_n989));
  INV_X1    g803(.A(new_n352), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n349), .B1(new_n344), .B2(new_n351), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n941), .B(new_n987), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n987), .B1(new_n962), .B2(new_n955), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n381), .A2(new_n349), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n900), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n989), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT127), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT127), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n989), .A2(new_n998), .A3(new_n992), .A4(new_n995), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(G57));
endmodule


