

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(G543), .A2(G651), .ZN(n680) );
  XOR2_X1 U550 ( .A(KEYINPUT1), .B(n551), .Z(n679) );
  NOR2_X2 U551 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  NOR2_X1 U552 ( .A1(n784), .A2(KEYINPUT33), .ZN(n785) );
  NOR2_X1 U553 ( .A1(G2105), .A2(n568), .ZN(n717) );
  INV_X1 U554 ( .A(KEYINPUT89), .ZN(n567) );
  NOR2_X1 U555 ( .A1(n746), .A2(G299), .ZN(n745) );
  AND2_X1 U556 ( .A1(n773), .A2(n769), .ZN(n521) );
  AND2_X1 U557 ( .A1(n528), .A2(n526), .ZN(n524) );
  NAND2_X1 U558 ( .A1(n525), .A2(KEYINPUT101), .ZN(n523) );
  NOR2_X1 U559 ( .A1(G164), .A2(G1384), .ZN(n830) );
  XNOR2_X1 U560 ( .A(n518), .B(n563), .ZN(n638) );
  NOR2_X1 U561 ( .A1(n566), .A2(n567), .ZN(n548) );
  NAND2_X1 U562 ( .A1(n566), .A2(n567), .ZN(n543) );
  XNOR2_X1 U563 ( .A(n719), .B(n718), .ZN(n721) );
  INV_X1 U564 ( .A(KEYINPUT23), .ZN(n718) );
  INV_X1 U565 ( .A(KEYINPUT65), .ZN(n722) );
  NOR2_X1 U566 ( .A1(n758), .A2(n947), .ZN(n742) );
  NAND2_X1 U567 ( .A1(n534), .A2(n513), .ZN(n533) );
  XNOR2_X1 U568 ( .A(KEYINPUT28), .B(KEYINPUT97), .ZN(n747) );
  AND2_X1 U569 ( .A1(n1003), .A2(n531), .ZN(n529) );
  NAND2_X1 U570 ( .A1(n772), .A2(n520), .ZN(n519) );
  XNOR2_X1 U571 ( .A(n522), .B(n530), .ZN(n784) );
  INV_X1 U572 ( .A(KEYINPUT64), .ZN(n530) );
  OR2_X1 U573 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U574 ( .A1(n614), .A2(n613), .ZN(n616) );
  NOR2_X1 U575 ( .A1(n555), .A2(G651), .ZN(n686) );
  NAND2_X1 U576 ( .A1(n543), .A2(n550), .ZN(n542) );
  NAND2_X1 U577 ( .A1(n546), .A2(n545), .ZN(n544) );
  NOR2_X1 U578 ( .A1(n725), .A2(n724), .ZN(G160) );
  XOR2_X1 U579 ( .A(n748), .B(n747), .Z(n513) );
  XOR2_X1 U580 ( .A(KEYINPUT103), .B(n794), .Z(n514) );
  OR2_X1 U581 ( .A1(n740), .A2(n739), .ZN(n515) );
  NOR2_X1 U582 ( .A1(n789), .A2(n788), .ZN(n516) );
  NOR2_X1 U583 ( .A1(n796), .A2(n783), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n519), .B(KEYINPUT32), .ZN(n781) );
  NAND2_X1 U585 ( .A1(n774), .A2(n521), .ZN(n520) );
  NAND2_X1 U586 ( .A1(n524), .A2(n523), .ZN(n522) );
  INV_X1 U587 ( .A(n790), .ZN(n525) );
  AND2_X1 U588 ( .A1(n527), .A2(n517), .ZN(n526) );
  OR2_X1 U589 ( .A1(n1003), .A2(n531), .ZN(n527) );
  NAND2_X1 U590 ( .A1(n790), .A2(n529), .ZN(n528) );
  INV_X1 U591 ( .A(KEYINPUT101), .ZN(n531) );
  XNOR2_X1 U592 ( .A(n533), .B(n532), .ZN(n753) );
  INV_X1 U593 ( .A(KEYINPUT29), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n515), .A2(n535), .ZN(n534) );
  XNOR2_X1 U595 ( .A(n745), .B(n536), .ZN(n535) );
  INV_X1 U596 ( .A(KEYINPUT98), .ZN(n536) );
  XNOR2_X1 U597 ( .A(n538), .B(n537), .ZN(n800) );
  INV_X1 U598 ( .A(KEYINPUT104), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n539), .A2(n514), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n540), .A2(n516), .ZN(n539) );
  XNOR2_X1 U601 ( .A(n785), .B(n541), .ZN(n540) );
  INV_X1 U602 ( .A(KEYINPUT102), .ZN(n541) );
  XNOR2_X1 U603 ( .A(n565), .B(n564), .ZN(n549) );
  INV_X1 U604 ( .A(n549), .ZN(n547) );
  NOR2_X2 U605 ( .A1(n544), .A2(n542), .ZN(G164) );
  NAND2_X1 U606 ( .A1(n549), .A2(n567), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n546) );
  BUF_X1 U608 ( .A(n638), .Z(n884) );
  NAND2_X2 U609 ( .A1(n727), .A2(n830), .ZN(n758) );
  AND2_X1 U610 ( .A1(n570), .A2(n569), .ZN(n550) );
  INV_X1 U611 ( .A(KEYINPUT99), .ZN(n760) );
  XNOR2_X1 U612 ( .A(n760), .B(KEYINPUT30), .ZN(n761) );
  INV_X1 U613 ( .A(KEYINPUT31), .ZN(n767) );
  NOR2_X1 U614 ( .A1(n796), .A2(G1966), .ZN(n777) );
  INV_X1 U615 ( .A(n829), .ZN(n727) );
  INV_X1 U616 ( .A(KEYINPUT17), .ZN(n563) );
  INV_X1 U617 ( .A(KEYINPUT13), .ZN(n611) );
  INV_X1 U618 ( .A(KEYINPUT78), .ZN(n577) );
  INV_X1 U619 ( .A(KEYINPUT105), .ZN(n835) );
  XNOR2_X1 U620 ( .A(n577), .B(KEYINPUT5), .ZN(n578) );
  XNOR2_X1 U621 ( .A(n579), .B(n578), .ZN(n580) );
  NAND2_X1 U622 ( .A1(n616), .A2(n615), .ZN(n996) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U624 ( .A(KEYINPUT7), .B(n582), .Z(G168) );
  INV_X1 U625 ( .A(G651), .ZN(n556) );
  NOR2_X1 U626 ( .A1(G543), .A2(n556), .ZN(n551) );
  NAND2_X1 U627 ( .A1(G65), .A2(n679), .ZN(n553) );
  XOR2_X1 U628 ( .A(KEYINPUT0), .B(G543), .Z(n555) );
  NAND2_X1 U629 ( .A1(G53), .A2(n686), .ZN(n552) );
  NAND2_X1 U630 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U631 ( .A(KEYINPUT71), .B(n554), .ZN(n561) );
  NAND2_X1 U632 ( .A1(G91), .A2(n680), .ZN(n559) );
  XNOR2_X2 U633 ( .A(n557), .B(KEYINPUT67), .ZN(n676) );
  NAND2_X1 U634 ( .A1(G78), .A2(n676), .ZN(n558) );
  AND2_X1 U635 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U636 ( .A1(n561), .A2(n560), .ZN(G299) );
  INV_X1 U637 ( .A(G2104), .ZN(n568) );
  NAND2_X1 U638 ( .A1(n717), .A2(G102), .ZN(n562) );
  XNOR2_X1 U639 ( .A(KEYINPUT87), .B(n562), .ZN(n566) );
  NAND2_X1 U640 ( .A1(n638), .A2(G138), .ZN(n565) );
  INV_X1 U641 ( .A(KEYINPUT88), .ZN(n564) );
  AND2_X1 U642 ( .A1(n568), .A2(G2105), .ZN(n879) );
  NAND2_X1 U643 ( .A1(G126), .A2(n879), .ZN(n570) );
  AND2_X1 U644 ( .A1(G2104), .A2(G2105), .ZN(n880) );
  NAND2_X1 U645 ( .A1(G114), .A2(n880), .ZN(n569) );
  NAND2_X1 U646 ( .A1(G63), .A2(n679), .ZN(n572) );
  NAND2_X1 U647 ( .A1(G51), .A2(n686), .ZN(n571) );
  NAND2_X1 U648 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U649 ( .A(KEYINPUT6), .B(n573), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n680), .A2(G89), .ZN(n574) );
  XNOR2_X1 U651 ( .A(n574), .B(KEYINPUT4), .ZN(n576) );
  NAND2_X1 U652 ( .A1(G76), .A2(n676), .ZN(n575) );
  NAND2_X1 U653 ( .A1(n576), .A2(n575), .ZN(n579) );
  NOR2_X1 U654 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U655 ( .A1(n680), .A2(G90), .ZN(n583) );
  XOR2_X1 U656 ( .A(KEYINPUT69), .B(n583), .Z(n585) );
  NAND2_X1 U657 ( .A1(n676), .A2(G77), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n586), .B(KEYINPUT9), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G64), .A2(n679), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n686), .A2(G52), .ZN(n589) );
  XOR2_X1 U663 ( .A(KEYINPUT68), .B(n589), .Z(n590) );
  NOR2_X1 U664 ( .A1(n591), .A2(n590), .ZN(G171) );
  XOR2_X1 U665 ( .A(G2446), .B(G2430), .Z(n593) );
  XNOR2_X1 U666 ( .A(G2451), .B(G2454), .ZN(n592) );
  XNOR2_X1 U667 ( .A(n593), .B(n592), .ZN(n594) );
  XOR2_X1 U668 ( .A(n594), .B(G2427), .Z(n596) );
  XNOR2_X1 U669 ( .A(G1341), .B(G1348), .ZN(n595) );
  XNOR2_X1 U670 ( .A(n596), .B(n595), .ZN(n600) );
  XOR2_X1 U671 ( .A(G2443), .B(KEYINPUT108), .Z(n598) );
  XNOR2_X1 U672 ( .A(G2438), .B(G2435), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n598), .B(n597), .ZN(n599) );
  XOR2_X1 U674 ( .A(n600), .B(n599), .Z(n601) );
  AND2_X1 U675 ( .A1(G14), .A2(n601), .ZN(G401) );
  INV_X1 U676 ( .A(G57), .ZN(G237) );
  INV_X1 U677 ( .A(G82), .ZN(G220) );
  NAND2_X1 U678 ( .A1(G94), .A2(G452), .ZN(n602) );
  XOR2_X1 U679 ( .A(KEYINPUT70), .B(n602), .Z(G173) );
  NAND2_X1 U680 ( .A1(G7), .A2(G661), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n603), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U682 ( .A(G223), .ZN(n853) );
  NAND2_X1 U683 ( .A1(n853), .A2(G567), .ZN(n604) );
  XNOR2_X1 U684 ( .A(n604), .B(KEYINPUT73), .ZN(n605) );
  XNOR2_X1 U685 ( .A(KEYINPUT11), .B(n605), .ZN(G234) );
  NAND2_X1 U686 ( .A1(G56), .A2(n679), .ZN(n606) );
  XOR2_X1 U687 ( .A(KEYINPUT14), .B(n606), .Z(n614) );
  NAND2_X1 U688 ( .A1(G81), .A2(n680), .ZN(n607) );
  XNOR2_X1 U689 ( .A(n607), .B(KEYINPUT74), .ZN(n608) );
  XNOR2_X1 U690 ( .A(n608), .B(KEYINPUT12), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n676), .A2(G68), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n610), .A2(n609), .ZN(n612) );
  XNOR2_X1 U693 ( .A(n612), .B(n611), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n686), .A2(G43), .ZN(n615) );
  INV_X1 U695 ( .A(G860), .ZN(n631) );
  OR2_X1 U696 ( .A1(n996), .A2(n631), .ZN(G153) );
  NAND2_X1 U697 ( .A1(G868), .A2(G171), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G54), .A2(n686), .ZN(n617) );
  XNOR2_X1 U699 ( .A(n617), .B(KEYINPUT76), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G92), .A2(n680), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G79), .A2(n676), .ZN(n618) );
  NAND2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G66), .A2(n679), .ZN(n620) );
  XNOR2_X1 U704 ( .A(KEYINPUT75), .B(n620), .ZN(n621) );
  NOR2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U707 ( .A(KEYINPUT15), .B(n625), .Z(n738) );
  INV_X1 U708 ( .A(n738), .ZN(n986) );
  INV_X1 U709 ( .A(G868), .ZN(n698) );
  NAND2_X1 U710 ( .A1(n986), .A2(n698), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U712 ( .A(n628), .B(KEYINPUT77), .ZN(G284) );
  NOR2_X1 U713 ( .A1(G286), .A2(n698), .ZN(n630) );
  NOR2_X1 U714 ( .A1(G868), .A2(G299), .ZN(n629) );
  NOR2_X1 U715 ( .A1(n630), .A2(n629), .ZN(G297) );
  NAND2_X1 U716 ( .A1(n631), .A2(G559), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n632), .A2(n986), .ZN(n633) );
  XNOR2_X1 U718 ( .A(n633), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U719 ( .A1(G868), .A2(n996), .ZN(n636) );
  NAND2_X1 U720 ( .A1(G868), .A2(n986), .ZN(n634) );
  NOR2_X1 U721 ( .A1(G559), .A2(n634), .ZN(n635) );
  NOR2_X1 U722 ( .A1(n636), .A2(n635), .ZN(G282) );
  NAND2_X1 U723 ( .A1(G123), .A2(n879), .ZN(n637) );
  XNOR2_X1 U724 ( .A(n637), .B(KEYINPUT18), .ZN(n645) );
  BUF_X1 U725 ( .A(n717), .Z(n883) );
  NAND2_X1 U726 ( .A1(G99), .A2(n883), .ZN(n640) );
  NAND2_X1 U727 ( .A1(G135), .A2(n884), .ZN(n639) );
  NAND2_X1 U728 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U729 ( .A1(G111), .A2(n880), .ZN(n641) );
  XNOR2_X1 U730 ( .A(KEYINPUT79), .B(n641), .ZN(n642) );
  NOR2_X1 U731 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n645), .A2(n644), .ZN(n873) );
  INV_X1 U733 ( .A(n873), .ZN(n939) );
  XOR2_X1 U734 ( .A(G2096), .B(n939), .Z(n646) );
  NOR2_X1 U735 ( .A1(G2100), .A2(n646), .ZN(n647) );
  XOR2_X1 U736 ( .A(KEYINPUT80), .B(n647), .Z(G156) );
  NAND2_X1 U737 ( .A1(G67), .A2(n679), .ZN(n649) );
  NAND2_X1 U738 ( .A1(G93), .A2(n680), .ZN(n648) );
  NAND2_X1 U739 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U740 ( .A1(G55), .A2(n686), .ZN(n650) );
  XNOR2_X1 U741 ( .A(KEYINPUT81), .B(n650), .ZN(n651) );
  NOR2_X1 U742 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U743 ( .A1(n676), .A2(G80), .ZN(n653) );
  NAND2_X1 U744 ( .A1(n654), .A2(n653), .ZN(n699) );
  NAND2_X1 U745 ( .A1(n986), .A2(G559), .ZN(n696) );
  XNOR2_X1 U746 ( .A(n996), .B(n696), .ZN(n655) );
  NOR2_X1 U747 ( .A1(G860), .A2(n655), .ZN(n656) );
  XOR2_X1 U748 ( .A(n699), .B(n656), .Z(G145) );
  NAND2_X1 U749 ( .A1(G49), .A2(n686), .ZN(n658) );
  NAND2_X1 U750 ( .A1(G74), .A2(G651), .ZN(n657) );
  NAND2_X1 U751 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U752 ( .A1(n679), .A2(n659), .ZN(n661) );
  NAND2_X1 U753 ( .A1(n555), .A2(G87), .ZN(n660) );
  NAND2_X1 U754 ( .A1(n661), .A2(n660), .ZN(G288) );
  NAND2_X1 U755 ( .A1(G62), .A2(n679), .ZN(n663) );
  NAND2_X1 U756 ( .A1(G50), .A2(n686), .ZN(n662) );
  NAND2_X1 U757 ( .A1(n663), .A2(n662), .ZN(n669) );
  NAND2_X1 U758 ( .A1(n680), .A2(G88), .ZN(n664) );
  XNOR2_X1 U759 ( .A(n664), .B(KEYINPUT84), .ZN(n666) );
  NAND2_X1 U760 ( .A1(G75), .A2(n676), .ZN(n665) );
  NAND2_X1 U761 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U762 ( .A(KEYINPUT85), .B(n667), .Z(n668) );
  NOR2_X1 U763 ( .A1(n669), .A2(n668), .ZN(G166) );
  AND2_X1 U764 ( .A1(n680), .A2(G85), .ZN(n673) );
  NAND2_X1 U765 ( .A1(G60), .A2(n679), .ZN(n671) );
  NAND2_X1 U766 ( .A1(G47), .A2(n686), .ZN(n670) );
  NAND2_X1 U767 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U768 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U769 ( .A1(n676), .A2(G72), .ZN(n674) );
  NAND2_X1 U770 ( .A1(n675), .A2(n674), .ZN(G290) );
  XOR2_X1 U771 ( .A(KEYINPUT2), .B(KEYINPUT82), .Z(n678) );
  NAND2_X1 U772 ( .A1(G73), .A2(n676), .ZN(n677) );
  XNOR2_X1 U773 ( .A(n678), .B(n677), .ZN(n684) );
  NAND2_X1 U774 ( .A1(G61), .A2(n679), .ZN(n682) );
  NAND2_X1 U775 ( .A1(G86), .A2(n680), .ZN(n681) );
  NAND2_X1 U776 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U777 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U778 ( .A(KEYINPUT83), .B(n685), .Z(n688) );
  NAND2_X1 U779 ( .A1(n686), .A2(G48), .ZN(n687) );
  NAND2_X1 U780 ( .A1(n688), .A2(n687), .ZN(G305) );
  XOR2_X1 U781 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n689) );
  XNOR2_X1 U782 ( .A(G299), .B(n689), .ZN(n690) );
  XNOR2_X1 U783 ( .A(n690), .B(G288), .ZN(n693) );
  XOR2_X1 U784 ( .A(G166), .B(G290), .Z(n691) );
  XNOR2_X1 U785 ( .A(n699), .B(n691), .ZN(n692) );
  XNOR2_X1 U786 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(G305), .ZN(n695) );
  XNOR2_X1 U788 ( .A(n695), .B(n996), .ZN(n900) );
  XNOR2_X1 U789 ( .A(n900), .B(n696), .ZN(n697) );
  NOR2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n701) );
  NOR2_X1 U791 ( .A1(G868), .A2(n699), .ZN(n700) );
  NOR2_X1 U792 ( .A1(n701), .A2(n700), .ZN(G295) );
  NAND2_X1 U793 ( .A1(G2078), .A2(G2084), .ZN(n702) );
  XOR2_X1 U794 ( .A(KEYINPUT20), .B(n702), .Z(n703) );
  NAND2_X1 U795 ( .A1(G2090), .A2(n703), .ZN(n704) );
  XNOR2_X1 U796 ( .A(KEYINPUT21), .B(n704), .ZN(n705) );
  NAND2_X1 U797 ( .A1(n705), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U798 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U799 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  NOR2_X1 U800 ( .A1(G219), .A2(G220), .ZN(n706) );
  XOR2_X1 U801 ( .A(KEYINPUT22), .B(n706), .Z(n707) );
  NOR2_X1 U802 ( .A1(G218), .A2(n707), .ZN(n708) );
  NAND2_X1 U803 ( .A1(G96), .A2(n708), .ZN(n933) );
  NAND2_X1 U804 ( .A1(n933), .A2(G2106), .ZN(n712) );
  NAND2_X1 U805 ( .A1(G69), .A2(G120), .ZN(n709) );
  NOR2_X1 U806 ( .A1(G237), .A2(n709), .ZN(n710) );
  NAND2_X1 U807 ( .A1(G108), .A2(n710), .ZN(n934) );
  NAND2_X1 U808 ( .A1(n934), .A2(G567), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n935) );
  NAND2_X1 U810 ( .A1(G661), .A2(G483), .ZN(n713) );
  NOR2_X1 U811 ( .A1(n935), .A2(n713), .ZN(n856) );
  NAND2_X1 U812 ( .A1(n856), .A2(G36), .ZN(G176) );
  XOR2_X1 U813 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  NAND2_X1 U814 ( .A1(n880), .A2(G113), .ZN(n715) );
  NAND2_X1 U815 ( .A1(n638), .A2(G137), .ZN(n714) );
  NAND2_X1 U816 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U817 ( .A(KEYINPUT66), .B(n716), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n717), .A2(G101), .ZN(n719) );
  NAND2_X1 U819 ( .A1(n879), .A2(G125), .ZN(n720) );
  NAND2_X1 U820 ( .A1(n721), .A2(n720), .ZN(n723) );
  XNOR2_X1 U821 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U822 ( .A1(G160), .A2(G40), .ZN(n829) );
  NAND2_X1 U823 ( .A1(G1348), .A2(n758), .ZN(n729) );
  INV_X1 U824 ( .A(n758), .ZN(n749) );
  NAND2_X1 U825 ( .A1(G2067), .A2(n749), .ZN(n728) );
  NAND2_X1 U826 ( .A1(n729), .A2(n728), .ZN(n737) );
  NOR2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n736) );
  INV_X1 U828 ( .A(n996), .ZN(n731) );
  NAND2_X1 U829 ( .A1(n758), .A2(G1341), .ZN(n730) );
  NAND2_X1 U830 ( .A1(n731), .A2(n730), .ZN(n734) );
  INV_X1 U831 ( .A(G1996), .ZN(n960) );
  NOR2_X1 U832 ( .A1(n758), .A2(n960), .ZN(n732) );
  XNOR2_X1 U833 ( .A(n732), .B(KEYINPUT26), .ZN(n733) );
  NOR2_X1 U834 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U835 ( .A1(n736), .A2(n735), .ZN(n740) );
  AND2_X1 U836 ( .A1(n738), .A2(n737), .ZN(n739) );
  INV_X1 U837 ( .A(G2072), .ZN(n947) );
  XNOR2_X1 U838 ( .A(KEYINPUT96), .B(KEYINPUT27), .ZN(n741) );
  XNOR2_X1 U839 ( .A(n742), .B(n741), .ZN(n744) );
  NAND2_X1 U840 ( .A1(n758), .A2(G1956), .ZN(n743) );
  NAND2_X1 U841 ( .A1(n744), .A2(n743), .ZN(n746) );
  NAND2_X1 U842 ( .A1(n746), .A2(G299), .ZN(n748) );
  INV_X1 U843 ( .A(G1961), .ZN(n1008) );
  NAND2_X1 U844 ( .A1(n758), .A2(n1008), .ZN(n751) );
  XNOR2_X1 U845 ( .A(G2078), .B(KEYINPUT25), .ZN(n962) );
  NAND2_X1 U846 ( .A1(n749), .A2(n962), .ZN(n750) );
  NAND2_X1 U847 ( .A1(n751), .A2(n750), .ZN(n764) );
  NAND2_X1 U848 ( .A1(G171), .A2(n764), .ZN(n752) );
  NAND2_X1 U849 ( .A1(n753), .A2(n752), .ZN(n774) );
  NAND2_X2 U850 ( .A1(n758), .A2(G8), .ZN(n796) );
  NOR2_X1 U851 ( .A1(G1971), .A2(n796), .ZN(n755) );
  NOR2_X1 U852 ( .A1(G2090), .A2(n758), .ZN(n754) );
  NOR2_X1 U853 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U854 ( .A1(G303), .A2(n756), .ZN(n757) );
  XNOR2_X1 U855 ( .A(n757), .B(KEYINPUT100), .ZN(n769) );
  NOR2_X1 U856 ( .A1(G2084), .A2(n758), .ZN(n775) );
  NOR2_X1 U857 ( .A1(n777), .A2(n775), .ZN(n759) );
  NAND2_X1 U858 ( .A1(G8), .A2(n759), .ZN(n762) );
  XNOR2_X1 U859 ( .A(n762), .B(n761), .ZN(n763) );
  NOR2_X1 U860 ( .A1(G168), .A2(n763), .ZN(n766) );
  NOR2_X1 U861 ( .A1(G171), .A2(n764), .ZN(n765) );
  NOR2_X1 U862 ( .A1(n766), .A2(n765), .ZN(n768) );
  XNOR2_X1 U863 ( .A(n768), .B(n767), .ZN(n773) );
  INV_X1 U864 ( .A(n769), .ZN(n770) );
  OR2_X1 U865 ( .A1(n770), .A2(G286), .ZN(n771) );
  AND2_X1 U866 ( .A1(G8), .A2(n771), .ZN(n772) );
  AND2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n779) );
  AND2_X1 U868 ( .A1(G8), .A2(n775), .ZN(n776) );
  OR2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n778) );
  OR2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n790) );
  NOR2_X1 U872 ( .A1(G1976), .A2(G288), .ZN(n786) );
  NOR2_X1 U873 ( .A1(G303), .A2(G1971), .ZN(n782) );
  NOR2_X1 U874 ( .A1(n786), .A2(n782), .ZN(n1003) );
  NAND2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n984) );
  INV_X1 U876 ( .A(n984), .ZN(n783) );
  XOR2_X1 U877 ( .A(G1981), .B(G305), .Z(n993) );
  INV_X1 U878 ( .A(n993), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n786), .A2(KEYINPUT33), .ZN(n787) );
  NOR2_X1 U880 ( .A1(n796), .A2(n787), .ZN(n788) );
  NOR2_X1 U881 ( .A1(G2090), .A2(G303), .ZN(n791) );
  NAND2_X1 U882 ( .A1(G8), .A2(n791), .ZN(n792) );
  NAND2_X1 U883 ( .A1(n790), .A2(n792), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n796), .A2(n793), .ZN(n794) );
  NOR2_X1 U885 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XNOR2_X1 U886 ( .A(n795), .B(KEYINPUT24), .ZN(n798) );
  INV_X1 U887 ( .A(n796), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n834) );
  XOR2_X1 U890 ( .A(G1986), .B(G290), .Z(n985) );
  XOR2_X1 U891 ( .A(G2067), .B(KEYINPUT37), .Z(n837) );
  XNOR2_X1 U892 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G128), .A2(n879), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G116), .A2(n880), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U896 ( .A(n803), .B(KEYINPUT35), .ZN(n804) );
  XNOR2_X1 U897 ( .A(n805), .B(n804), .ZN(n811) );
  NAND2_X1 U898 ( .A1(G104), .A2(n883), .ZN(n807) );
  NAND2_X1 U899 ( .A1(G140), .A2(n884), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U901 ( .A(n808), .B(KEYINPUT34), .ZN(n809) );
  XNOR2_X1 U902 ( .A(KEYINPUT92), .B(n809), .ZN(n810) );
  NOR2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U904 ( .A(KEYINPUT36), .B(n812), .Z(n876) );
  AND2_X1 U905 ( .A1(n837), .A2(n876), .ZN(n845) );
  NAND2_X1 U906 ( .A1(G119), .A2(n879), .ZN(n814) );
  NAND2_X1 U907 ( .A1(G131), .A2(n884), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n818) );
  NAND2_X1 U909 ( .A1(G95), .A2(n883), .ZN(n816) );
  NAND2_X1 U910 ( .A1(G107), .A2(n880), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n817) );
  OR2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n890) );
  NAND2_X1 U913 ( .A1(G1991), .A2(n890), .ZN(n828) );
  NAND2_X1 U914 ( .A1(G105), .A2(n883), .ZN(n819) );
  XOR2_X1 U915 ( .A(KEYINPUT38), .B(n819), .Z(n824) );
  NAND2_X1 U916 ( .A1(G129), .A2(n879), .ZN(n821) );
  NAND2_X1 U917 ( .A1(G117), .A2(n880), .ZN(n820) );
  NAND2_X1 U918 ( .A1(n821), .A2(n820), .ZN(n822) );
  XOR2_X1 U919 ( .A(KEYINPUT95), .B(n822), .Z(n823) );
  NOR2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n884), .A2(G141), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n872) );
  NAND2_X1 U923 ( .A1(G1996), .A2(n872), .ZN(n827) );
  NAND2_X1 U924 ( .A1(n828), .A2(n827), .ZN(n841) );
  NOR2_X1 U925 ( .A1(n845), .A2(n841), .ZN(n942) );
  NAND2_X1 U926 ( .A1(n985), .A2(n942), .ZN(n832) );
  NOR2_X1 U927 ( .A1(n830), .A2(n829), .ZN(n831) );
  XOR2_X1 U928 ( .A(KEYINPUT91), .B(n831), .Z(n848) );
  NAND2_X1 U929 ( .A1(n832), .A2(n848), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n834), .A2(n833), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n836), .B(n835), .ZN(n851) );
  NOR2_X1 U932 ( .A1(n837), .A2(n876), .ZN(n956) );
  NOR2_X1 U933 ( .A1(G1996), .A2(n872), .ZN(n838) );
  XNOR2_X1 U934 ( .A(KEYINPUT106), .B(n838), .ZN(n937) );
  NOR2_X1 U935 ( .A1(G1991), .A2(n890), .ZN(n940) );
  NOR2_X1 U936 ( .A1(G1986), .A2(G290), .ZN(n839) );
  NOR2_X1 U937 ( .A1(n940), .A2(n839), .ZN(n840) );
  NOR2_X1 U938 ( .A1(n841), .A2(n840), .ZN(n842) );
  NOR2_X1 U939 ( .A1(n937), .A2(n842), .ZN(n843) );
  XOR2_X1 U940 ( .A(KEYINPUT39), .B(n843), .Z(n844) );
  NOR2_X1 U941 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U942 ( .A1(n956), .A2(n846), .ZN(n847) );
  XNOR2_X1 U943 ( .A(KEYINPUT107), .B(n847), .ZN(n849) );
  NAND2_X1 U944 ( .A1(n849), .A2(n848), .ZN(n850) );
  NAND2_X1 U945 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U946 ( .A(n852), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U947 ( .A1(G2106), .A2(n853), .ZN(G217) );
  AND2_X1 U948 ( .A1(G15), .A2(G2), .ZN(n854) );
  NAND2_X1 U949 ( .A1(G661), .A2(n854), .ZN(G259) );
  NAND2_X1 U950 ( .A1(G3), .A2(G1), .ZN(n855) );
  NAND2_X1 U951 ( .A1(n856), .A2(n855), .ZN(G188) );
  NAND2_X1 U952 ( .A1(G124), .A2(n879), .ZN(n857) );
  XNOR2_X1 U953 ( .A(n857), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U954 ( .A1(G136), .A2(n884), .ZN(n858) );
  XOR2_X1 U955 ( .A(KEYINPUT111), .B(n858), .Z(n859) );
  NAND2_X1 U956 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U957 ( .A1(G100), .A2(n883), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G112), .A2(n880), .ZN(n861) );
  NAND2_X1 U959 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U960 ( .A1(n864), .A2(n863), .ZN(G162) );
  NAND2_X1 U961 ( .A1(G103), .A2(n883), .ZN(n866) );
  NAND2_X1 U962 ( .A1(G139), .A2(n884), .ZN(n865) );
  NAND2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n871) );
  NAND2_X1 U964 ( .A1(G127), .A2(n879), .ZN(n868) );
  NAND2_X1 U965 ( .A1(G115), .A2(n880), .ZN(n867) );
  NAND2_X1 U966 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U967 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n946) );
  XOR2_X1 U969 ( .A(G162), .B(n946), .Z(n878) );
  XNOR2_X1 U970 ( .A(G160), .B(n872), .ZN(n874) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U973 ( .A(n878), .B(n877), .ZN(n897) );
  NAND2_X1 U974 ( .A1(G130), .A2(n879), .ZN(n882) );
  NAND2_X1 U975 ( .A1(G118), .A2(n880), .ZN(n881) );
  NAND2_X1 U976 ( .A1(n882), .A2(n881), .ZN(n889) );
  NAND2_X1 U977 ( .A1(G106), .A2(n883), .ZN(n886) );
  NAND2_X1 U978 ( .A1(G142), .A2(n884), .ZN(n885) );
  NAND2_X1 U979 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U980 ( .A(n887), .B(KEYINPUT45), .Z(n888) );
  NOR2_X1 U981 ( .A1(n889), .A2(n888), .ZN(n891) );
  XNOR2_X1 U982 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U983 ( .A(n892), .B(KEYINPUT48), .Z(n894) );
  XNOR2_X1 U984 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n893) );
  XNOR2_X1 U985 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U986 ( .A(G164), .B(n895), .ZN(n896) );
  XNOR2_X1 U987 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U988 ( .A1(G37), .A2(n898), .ZN(n899) );
  XOR2_X1 U989 ( .A(KEYINPUT113), .B(n899), .Z(G395) );
  XOR2_X1 U990 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n902) );
  XNOR2_X1 U991 ( .A(n986), .B(n900), .ZN(n901) );
  XNOR2_X1 U992 ( .A(n902), .B(n901), .ZN(n904) );
  XOR2_X1 U993 ( .A(G286), .B(G171), .Z(n903) );
  XNOR2_X1 U994 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U995 ( .A1(G37), .A2(n905), .ZN(n906) );
  XNOR2_X1 U996 ( .A(KEYINPUT116), .B(n906), .ZN(G397) );
  XOR2_X1 U997 ( .A(G2100), .B(G2096), .Z(n908) );
  XNOR2_X1 U998 ( .A(KEYINPUT42), .B(G2678), .ZN(n907) );
  XNOR2_X1 U999 ( .A(n908), .B(n907), .ZN(n912) );
  XOR2_X1 U1000 ( .A(KEYINPUT43), .B(G2090), .Z(n910) );
  XNOR2_X1 U1001 ( .A(G2067), .B(G2072), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1003 ( .A(n912), .B(n911), .Z(n914) );
  XNOR2_X1 U1004 ( .A(G2078), .B(G2084), .ZN(n913) );
  XNOR2_X1 U1005 ( .A(n914), .B(n913), .ZN(G227) );
  XOR2_X1 U1006 ( .A(KEYINPUT110), .B(G1956), .Z(n916) );
  XNOR2_X1 U1007 ( .A(G1996), .B(G1991), .ZN(n915) );
  XNOR2_X1 U1008 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1009 ( .A(n917), .B(KEYINPUT41), .Z(n919) );
  XNOR2_X1 U1010 ( .A(G1981), .B(G1966), .ZN(n918) );
  XNOR2_X1 U1011 ( .A(n919), .B(n918), .ZN(n923) );
  XOR2_X1 U1012 ( .A(G1961), .B(G1971), .Z(n921) );
  XNOR2_X1 U1013 ( .A(G1986), .B(G1976), .ZN(n920) );
  XNOR2_X1 U1014 ( .A(n921), .B(n920), .ZN(n922) );
  XOR2_X1 U1015 ( .A(n923), .B(n922), .Z(n925) );
  XNOR2_X1 U1016 ( .A(G2474), .B(KEYINPUT109), .ZN(n924) );
  XNOR2_X1 U1017 ( .A(n925), .B(n924), .ZN(G229) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n926) );
  XNOR2_X1 U1019 ( .A(KEYINPUT118), .B(n926), .ZN(n932) );
  NOR2_X1 U1020 ( .A1(n935), .A2(G401), .ZN(n927) );
  XNOR2_X1 U1021 ( .A(n927), .B(KEYINPUT117), .ZN(n930) );
  NOR2_X1 U1022 ( .A1(G227), .A2(G229), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(KEYINPUT49), .B(n928), .ZN(n929) );
  NOR2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(G225) );
  XNOR2_X1 U1026 ( .A(KEYINPUT119), .B(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(G120), .ZN(G236) );
  INV_X1 U1029 ( .A(G96), .ZN(G221) );
  INV_X1 U1030 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(G325) );
  INV_X1 U1032 ( .A(G325), .ZN(G261) );
  INV_X1 U1033 ( .A(G171), .ZN(G301) );
  INV_X1 U1034 ( .A(n935), .ZN(G319) );
  INV_X1 U1035 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1038 ( .A(KEYINPUT51), .B(n938), .Z(n954) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n944) );
  XOR2_X1 U1041 ( .A(G2084), .B(G160), .Z(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1043 ( .A(KEYINPUT120), .B(n945), .Z(n952) );
  XOR2_X1 U1044 ( .A(G164), .B(G2078), .Z(n949) );
  XNOR2_X1 U1045 ( .A(n947), .B(n946), .ZN(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1047 ( .A(KEYINPUT50), .B(n950), .Z(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(KEYINPUT52), .B(n957), .ZN(n958) );
  INV_X1 U1052 ( .A(KEYINPUT55), .ZN(n980) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n980), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n959), .A2(G29), .ZN(n1038) );
  XOR2_X1 U1055 ( .A(G1991), .B(G25), .Z(n970) );
  XNOR2_X1 U1056 ( .A(G32), .B(n960), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(n961), .A2(G28), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(G27), .B(n962), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(G2067), .B(G26), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(G33), .B(G2072), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT53), .B(n971), .ZN(n973) );
  XOR2_X1 U1066 ( .A(G2090), .B(G35), .Z(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(KEYINPUT121), .B(n974), .ZN(n978) );
  XOR2_X1 U1069 ( .A(KEYINPUT122), .B(G34), .Z(n976) );
  XNOR2_X1 U1070 ( .A(G2084), .B(KEYINPUT54), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(n976), .B(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(n980), .B(n979), .ZN(n982) );
  INV_X1 U1074 ( .A(G29), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1076 ( .A1(G11), .A2(n983), .ZN(n1036) );
  XNOR2_X1 U1077 ( .A(G16), .B(KEYINPUT56), .ZN(n1007) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(G1348), .B(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(G1971), .A2(G303), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n992) );
  XOR2_X1 U1083 ( .A(G1956), .B(G299), .Z(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n1002) );
  XNOR2_X1 U1085 ( .A(G1966), .B(G168), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n995), .B(KEYINPUT57), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(G301), .B(G1961), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(n996), .B(G1341), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(KEYINPUT123), .B(n1005), .Z(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1034) );
  INV_X1 U1096 ( .A(G16), .ZN(n1032) );
  XNOR2_X1 U1097 ( .A(G5), .B(n1008), .ZN(n1025) );
  XOR2_X1 U1098 ( .A(G1348), .B(KEYINPUT59), .Z(n1009) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(G20), .B(G1956), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G1981), .B(G6), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(G19), .B(G1341), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(n1016), .B(KEYINPUT60), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(G1976), .B(G23), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(G1971), .B(G22), .ZN(n1017) );
  NOR2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1110 ( .A(G1986), .B(G24), .Z(n1019) );
  NAND2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1112 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(G21), .B(G1966), .ZN(n1026) );
  XNOR2_X1 U1116 ( .A(KEYINPUT124), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1117 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1118 ( .A(n1029), .B(KEYINPUT125), .Z(n1030) );
  XNOR2_X1 U1119 ( .A(KEYINPUT61), .B(n1030), .ZN(n1031) );
  NAND2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1121 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NOR2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1124 ( .A(n1039), .B(KEYINPUT62), .ZN(n1040) );
  XNOR2_X1 U1125 ( .A(KEYINPUT126), .B(n1040), .ZN(G150) );
  INV_X1 U1126 ( .A(G150), .ZN(G311) );
endmodule

