//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n605, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G69), .Z(G235));
  XNOR2_X1  g013(.A(KEYINPUT68), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT69), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G236), .A3(G237), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT70), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT73), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT72), .B(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(new_n460), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT72), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(KEYINPUT72), .ZN(new_n469));
  OAI211_X1 g044(.A(new_n462), .B(KEYINPUT3), .C1(new_n467), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n465), .A2(G137), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NOR3_X1   g047(.A1(new_n467), .A2(new_n469), .A3(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT74), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT74), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n472), .A2(new_n477), .A3(new_n474), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G113), .ZN(new_n481));
  OR3_X1    g056(.A1(new_n481), .A2(new_n468), .A3(KEYINPUT71), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT71), .B1(new_n481), .B2(new_n468), .ZN(new_n483));
  INV_X1    g058(.A(G125), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n461), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n482), .B(new_n483), .C1(new_n484), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G160));
  NAND2_X1  g065(.A1(new_n465), .A2(new_n470), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(new_n471), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n491), .A2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  OR2_X1    g070(.A1(G100), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR4_X1   g075(.A1(new_n486), .A2(KEYINPUT4), .A3(new_n500), .A4(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n465), .A2(G138), .A3(new_n470), .A4(new_n471), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n465), .A2(G126), .A3(new_n470), .A4(G2105), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n471), .A2(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  OR3_X1    g081(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT75), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT75), .B1(new_n505), .B2(new_n506), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n503), .A2(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT76), .Z(new_n523));
  NAND2_X1  g098(.A1(new_n516), .A2(new_n520), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G88), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n523), .A2(KEYINPUT77), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(KEYINPUT77), .B1(new_n523), .B2(new_n526), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n519), .B1(new_n527), .B2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND3_X1  g105(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT78), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n520), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI221_X1 g112(.A(new_n534), .B1(new_n535), .B2(new_n536), .C1(new_n524), .C2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n532), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n518), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT79), .B(G90), .Z(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n524), .A2(new_n542), .B1(new_n535), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n541), .A2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n524), .A2(new_n547), .B1(new_n535), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n516), .A2(G56), .ZN(new_n551));
  INV_X1    g126(.A(G68), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(new_n512), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT80), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n553), .B2(new_n554), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n550), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(new_n521), .A2(G53), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n525), .A2(G91), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n567), .B(new_n568), .C1(new_n518), .C2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G168), .ZN(G286));
  NAND2_X1  g146(.A1(new_n525), .A2(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n521), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(new_n525), .A2(G86), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT82), .Z(new_n577));
  NAND2_X1  g152(.A1(new_n516), .A2(G61), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(KEYINPUT81), .B1(G73), .B2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n579), .B1(KEYINPUT81), .B2(new_n578), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G48), .B2(new_n521), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n525), .A2(G85), .B1(G47), .B2(new_n521), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n518), .B2(new_n584), .ZN(G290));
  INV_X1    g160(.A(G868), .ZN(new_n586));
  NOR2_X1   g161(.A1(G171), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  XNOR2_X1  g164(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n590));
  OR3_X1    g165(.A1(new_n524), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n524), .B2(new_n589), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G54), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n594), .A2(new_n518), .B1(new_n595), .B2(new_n535), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n588), .B1(G868), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT83), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(KEYINPUT83), .B2(new_n587), .ZN(G284));
  OAI21_X1  g175(.A(new_n599), .B1(KEYINPUT83), .B2(new_n587), .ZN(G321));
  NAND2_X1  g176(.A1(G299), .A2(new_n586), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n586), .B2(G168), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(new_n586), .B2(G168), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n558), .A2(new_n586), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n593), .A2(new_n596), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n609), .B2(new_n586), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g186(.A1(new_n473), .A2(new_n461), .A3(new_n485), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n492), .A2(G123), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n494), .A2(G135), .ZN(new_n617));
  OR2_X1    g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G111), .C2(new_n471), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n615), .A2(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(KEYINPUT14), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n628), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(G401));
  XNOR2_X1  g213(.A(G2072), .B(G2078), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT87), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2084), .B(G2090), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT86), .ZN(new_n642));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n645));
  OAI21_X1  g220(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2096), .B(G2100), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n642), .A2(new_n643), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n645), .B1(new_n650), .B2(new_n644), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n648), .B(new_n651), .Z(G227));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT89), .ZN(new_n654));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n655), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n658), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n654), .A2(KEYINPUT90), .A3(new_n655), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(new_n665), .A3(new_n658), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT91), .B(KEYINPUT20), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n661), .B(new_n662), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  OR3_X1    g244(.A1(new_n668), .A2(new_n669), .A3(G1991), .ZN(new_n670));
  OAI21_X1  g245(.A(G1991), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  AND3_X1   g246(.A1(new_n670), .A2(G1996), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(G1996), .B1(new_n670), .B2(new_n671), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n676), .B2(new_n677), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(G229));
  NAND2_X1  g257(.A1(G299), .A2(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(KEYINPUT23), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G20), .ZN(new_n686));
  MUX2_X1   g261(.A(KEYINPUT23), .B(new_n684), .S(new_n686), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1956), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n558), .A2(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n685), .A2(G19), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G1341), .ZN(new_n692));
  NOR2_X1   g267(.A1(G5), .A2(G16), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G171), .B2(G16), .ZN(new_n694));
  OAI22_X1  g269(.A1(new_n691), .A2(new_n692), .B1(new_n694), .B2(G1961), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n685), .A2(G4), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n597), .B2(new_n685), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1348), .ZN(new_n699));
  NOR4_X1   g274(.A1(new_n688), .A2(new_n695), .A3(new_n696), .A4(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(KEYINPUT92), .A2(G29), .ZN(new_n701));
  NOR2_X1   g276(.A1(KEYINPUT92), .A2(G29), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G35), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G162), .B2(new_n704), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT29), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G2090), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(G26), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT94), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n492), .A2(G128), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n494), .A2(G140), .ZN(new_n713));
  OR2_X1    g288(.A1(G104), .A2(G2105), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n714), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT93), .Z(new_n716));
  NAND3_X1  g291(.A1(new_n712), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n711), .B1(new_n717), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G2067), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n704), .A2(G27), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G164), .B2(new_n704), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n719), .B1(G2078), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G2078), .B2(new_n721), .ZN(new_n723));
  OAI22_X1  g298(.A1(KEYINPUT97), .A2(G2072), .B1(G29), .B2(G33), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n494), .A2(G139), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT95), .B(KEYINPUT25), .Z(new_n726));
  NAND3_X1  g301(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n461), .A2(new_n485), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n729), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n725), .B(new_n728), .C1(new_n471), .C2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT96), .Z(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n724), .B1(new_n733), .B2(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(KEYINPUT97), .A2(G2072), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n700), .A2(new_n708), .A3(new_n723), .A4(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT24), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(G34), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(G34), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n704), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n489), .B2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G2084), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n694), .A2(G1961), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT101), .Z(new_n747));
  NOR2_X1   g322(.A1(G168), .A2(new_n685), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n685), .B2(G21), .ZN(new_n749));
  INV_X1    g324(.A(G1966), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT31), .B(G11), .Z(new_n752));
  XOR2_X1   g327(.A(KEYINPUT100), .B(KEYINPUT30), .Z(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(G28), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n753), .B2(G28), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n620), .A2(new_n704), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n749), .B2(new_n750), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n747), .A2(new_n751), .A3(new_n756), .A4(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT102), .Z(new_n760));
  NOR3_X1   g335(.A1(new_n737), .A2(new_n745), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n742), .A2(G32), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n494), .A2(G141), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT98), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n492), .A2(G129), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT26), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n473), .A2(G105), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n764), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT99), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n762), .B1(new_n773), .B2(new_n742), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT27), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1996), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n761), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n685), .A2(G22), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n685), .ZN(new_n779));
  INV_X1    g354(.A(G1971), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G23), .ZN(new_n782));
  INV_X1    g357(.A(G288), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G16), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT33), .B(G1976), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G305), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(new_n685), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G6), .B2(new_n685), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT32), .B(G1981), .Z(new_n790));
  AOI21_X1  g365(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n781), .B(new_n791), .C1(new_n789), .C2(new_n790), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT34), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n492), .A2(G119), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n494), .A2(G131), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n471), .A2(G107), .ZN(new_n796));
  OAI21_X1  g371(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n794), .B(new_n795), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G25), .B(new_n798), .S(new_n703), .Z(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT35), .B(G1991), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G24), .B(G290), .S(G16), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1986), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n793), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(KEYINPUT36), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT36), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n793), .A2(new_n807), .A3(new_n804), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n777), .B1(new_n806), .B2(new_n808), .ZN(G311));
  INV_X1    g384(.A(G311), .ZN(G150));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  INV_X1    g386(.A(G55), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n524), .A2(new_n811), .B1(new_n535), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT104), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(new_n518), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n559), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n558), .A2(new_n816), .A3(new_n814), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n597), .A2(G559), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT39), .Z(new_n825));
  AOI21_X1  g400(.A(G860), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n825), .B2(new_n823), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n817), .A2(G860), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(G145));
  INV_X1    g405(.A(KEYINPUT106), .ZN(new_n831));
  INV_X1    g406(.A(new_n717), .ZN(new_n832));
  INV_X1    g407(.A(new_n510), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT105), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n835));
  INV_X1    g410(.A(new_n501), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g412(.A(KEYINPUT105), .B(new_n501), .C1(new_n502), .C2(KEYINPUT4), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n773), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n771), .B(KEYINPUT99), .ZN(new_n841));
  INV_X1    g416(.A(new_n839), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n832), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n840), .A2(new_n843), .A3(new_n832), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n731), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n846), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n733), .B1(new_n848), .B2(new_n844), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n494), .A2(G142), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n471), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G130), .B2(new_n492), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G162), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n489), .B(new_n620), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n798), .B(new_n613), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n847), .A2(new_n849), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n859), .B1(new_n847), .B2(new_n849), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n831), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n847), .A2(new_n849), .ZN(new_n865));
  INV_X1    g440(.A(new_n859), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n867), .A2(KEYINPUT106), .A3(new_n861), .A4(new_n860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT40), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT40), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n864), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(G395));
  NAND2_X1  g448(.A1(new_n817), .A2(new_n586), .ZN(new_n874));
  AND2_X1   g449(.A1(G303), .A2(new_n787), .ZN(new_n875));
  NOR2_X1   g450(.A1(G303), .A2(new_n787), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(G288), .B(KEYINPUT108), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G290), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n875), .B2(new_n876), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(KEYINPUT109), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(G299), .B(new_n597), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(KEYINPUT41), .ZN(new_n888));
  NAND2_X1  g463(.A1(G299), .A2(new_n597), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT107), .ZN(new_n890));
  XNOR2_X1  g465(.A(G299), .B(new_n608), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(KEYINPUT107), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n888), .B1(new_n892), .B2(KEYINPUT41), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n820), .B(new_n609), .ZN(new_n894));
  MUX2_X1   g469(.A(new_n893), .B(new_n892), .S(new_n894), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n886), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n874), .B1(new_n896), .B2(new_n586), .ZN(G295));
  OAI21_X1  g472(.A(new_n874), .B1(new_n896), .B2(new_n586), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT112), .ZN(new_n899));
  XNOR2_X1  g474(.A(G168), .B(G301), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n820), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n820), .A2(new_n900), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n892), .A2(new_n901), .A3(new_n902), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n893), .A2(new_n903), .B1(new_n904), .B2(KEYINPUT111), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n904), .A2(KEYINPUT111), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n899), .B(new_n861), .C1(new_n907), .C2(new_n883), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n883), .B1(new_n905), .B2(new_n906), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT112), .B1(new_n909), .B2(G37), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n905), .A2(new_n883), .A3(new_n906), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT113), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT43), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT113), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n912), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n903), .A2(KEYINPUT41), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n883), .B1(new_n918), .B2(new_n887), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n918), .A2(new_n892), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n861), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n916), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT44), .B1(new_n914), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n911), .B2(new_n913), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n916), .A2(new_n922), .A3(KEYINPUT43), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n925), .B1(new_n928), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g504(.A(G1384), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n839), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n488), .A2(G40), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n476), .A2(new_n934), .A3(new_n478), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT114), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n936), .B(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n717), .B(G2067), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT45), .B1(new_n839), .B2(new_n930), .ZN(new_n942));
  INV_X1    g517(.A(G1996), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n935), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n938), .A2(new_n841), .ZN(new_n945));
  OAI221_X1 g520(.A(new_n941), .B1(new_n841), .B2(new_n944), .C1(new_n945), .C2(new_n943), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT115), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n798), .A2(new_n800), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G2067), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n832), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n939), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n798), .A2(new_n800), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n938), .B1(new_n953), .B2(new_n948), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n936), .A2(G1986), .A3(G290), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT48), .Z(new_n956));
  NAND3_X1  g531(.A1(new_n947), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n944), .B(KEYINPUT46), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n945), .A2(new_n941), .A3(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT47), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n952), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT49), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT119), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n581), .A2(new_n576), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(G1981), .ZN(new_n966));
  INV_X1    g541(.A(G1981), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n577), .A2(new_n581), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n964), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n581), .B2(new_n576), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(KEYINPUT119), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n963), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n577), .A2(new_n581), .A3(new_n967), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT119), .B1(new_n973), .B2(new_n970), .ZN(new_n974));
  INV_X1    g549(.A(new_n971), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n975), .A3(KEYINPUT49), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n839), .A2(new_n930), .A3(new_n935), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n977), .A2(G8), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1976), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n977), .B(G8), .C1(new_n980), .C2(G288), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n783), .A2(G1976), .ZN(new_n982));
  OR3_X1    g557(.A1(new_n981), .A2(KEYINPUT52), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(KEYINPUT52), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n979), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n986));
  AND3_X1   g561(.A1(G303), .A2(G8), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(G303), .A2(G8), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(KEYINPUT118), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n987), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n930), .B1(new_n503), .B2(new_n510), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n935), .B1(new_n993), .B2(KEYINPUT45), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n839), .A2(KEYINPUT45), .A3(new_n930), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n839), .A2(KEYINPUT116), .A3(KEYINPUT45), .A4(new_n930), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G1971), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n476), .A2(new_n934), .A3(new_n478), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(KEYINPUT117), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n839), .A2(new_n1004), .A3(new_n930), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n992), .A2(new_n1006), .A3(KEYINPUT50), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1003), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G2090), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n991), .B(G8), .C1(new_n1000), .C2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n985), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n931), .A2(KEYINPUT50), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n993), .A2(new_n1004), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1012), .A2(new_n935), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI22_X1  g590(.A1(new_n1015), .A2(G2090), .B1(new_n999), .B2(G1971), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n991), .B1(new_n1016), .B2(G8), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n935), .B1(new_n932), .B2(new_n992), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n750), .B1(new_n942), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1003), .A2(new_n1005), .A3(new_n744), .A4(new_n1007), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(G8), .A3(G168), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1011), .A2(new_n1017), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(G8), .B1(new_n1000), .B2(new_n1009), .ZN(new_n1024));
  INV_X1    g599(.A(new_n991), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1023), .A2(KEYINPUT63), .B1(new_n1011), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1010), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n979), .A2(new_n980), .A3(new_n783), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n968), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1031), .A2(new_n985), .B1(new_n1033), .B2(new_n978), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1036), .B(G8), .C1(new_n1021), .C2(G286), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G168), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1021), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  AOI211_X1 g616(.A(new_n1036), .B(new_n1039), .C1(new_n1021), .C2(G8), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT124), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1039), .B1(new_n1021), .B2(G8), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT51), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT124), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n1040), .A4(new_n1037), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT62), .ZN(new_n1049));
  INV_X1    g624(.A(G2078), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n999), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  INV_X1    g627(.A(G1961), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1051), .A2(new_n1052), .B1(new_n1053), .B2(new_n1008), .ZN(new_n1054));
  OR4_X1    g629(.A1(new_n1052), .A2(new_n942), .A3(new_n1018), .A4(G2078), .ZN(new_n1055));
  AOI21_X1  g630(.A(G301), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT62), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1043), .A2(new_n1057), .A3(new_n1047), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1049), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT56), .B(G2072), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n999), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(G1956), .B2(new_n1014), .ZN(new_n1062));
  XNOR2_X1  g637(.A(G299), .B(KEYINPUT57), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  INV_X1    g640(.A(G1348), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1008), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n977), .A2(KEYINPUT120), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n839), .A2(new_n935), .A3(new_n1069), .A4(new_n930), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n950), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n597), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1064), .B1(new_n1065), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n1075));
  AOI211_X1 g650(.A(G1996), .B(new_n994), .C1(new_n997), .C2(new_n998), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT58), .B(G1341), .Z(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1075), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n997), .A2(new_n998), .ZN(new_n1081));
  INV_X1    g656(.A(new_n994), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n943), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1077), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(KEYINPUT121), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT59), .B1(new_n1087), .B2(new_n559), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n1089));
  AOI211_X1 g664(.A(new_n1089), .B(new_n558), .C1(new_n1080), .C2(new_n1086), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1072), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n597), .B1(new_n1072), .B2(new_n1092), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1067), .A2(new_n1071), .A3(KEYINPUT60), .A4(new_n608), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1096), .A2(new_n1095), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1093), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1074), .B1(new_n1091), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n933), .B1(new_n479), .B2(KEYINPUT125), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(KEYINPUT125), .B2(new_n479), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1103), .A2(KEYINPUT126), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n942), .A2(new_n1052), .A3(G2078), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(KEYINPUT126), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1104), .A2(new_n1081), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1008), .A2(new_n1053), .ZN(new_n1108));
  AOI211_X1 g683(.A(G2078), .B(new_n994), .C1(new_n997), .C2(new_n998), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1107), .B(new_n1108), .C1(KEYINPUT53), .C2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(G171), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1101), .B1(new_n1056), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1054), .A2(G301), .A3(new_n1055), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1110), .A2(G171), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1114), .A3(KEYINPUT54), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1014), .A2(G1956), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1063), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(KEYINPUT61), .A3(new_n1117), .A4(new_n1061), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1072), .A2(new_n597), .B1(KEYINPUT122), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1065), .B(new_n1118), .C1(new_n1064), .C2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1112), .A2(new_n1115), .A3(new_n1048), .A4(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1059), .B1(new_n1100), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1035), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(G290), .B(G1986), .Z(new_n1126));
  OAI211_X1 g701(.A(new_n947), .B(new_n954), .C1(new_n936), .C2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n962), .B1(new_n1125), .B2(new_n1127), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g703(.A1(new_n913), .A2(new_n923), .A3(new_n861), .A4(new_n921), .ZN(new_n1130));
  AOI21_X1  g704(.A(new_n916), .B1(new_n910), .B2(new_n908), .ZN(new_n1131));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1131), .B2(new_n923), .ZN(new_n1132));
  INV_X1    g706(.A(G319), .ZN(new_n1133));
  NOR3_X1   g707(.A1(G401), .A2(new_n1133), .A3(G227), .ZN(new_n1134));
  NAND3_X1  g708(.A1(new_n680), .A2(new_n681), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g709(.A(new_n1135), .B1(new_n864), .B2(new_n868), .ZN(new_n1136));
  AND2_X1   g710(.A1(new_n1132), .A2(new_n1136), .ZN(G308));
  NAND2_X1  g711(.A1(new_n1132), .A2(new_n1136), .ZN(G225));
endmodule


