//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT64), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT65), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(G137), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(new_n468), .ZN(G160));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  NOR3_X1   g050(.A1(new_n474), .A2(new_n475), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(KEYINPUT67), .B1(new_n462), .B2(new_n461), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n474), .A2(new_n461), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n471), .A2(new_n473), .A3(G126), .A4(G2105), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n462), .A2(KEYINPUT68), .A3(G126), .A4(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(new_n461), .B2(G114), .ZN(new_n491));
  NOR2_X1   g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT69), .B(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n462), .A2(new_n495), .A3(G138), .A4(new_n461), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n471), .A2(new_n473), .A3(G138), .A4(new_n461), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(KEYINPUT69), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n490), .A2(new_n494), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(G50), .A3(G543), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT70), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n505), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n504), .B1(new_n516), .B2(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n512), .B1(new_n507), .B2(new_n510), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n502), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT71), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n518), .A2(new_n521), .A3(new_n502), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT72), .B(G88), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(G166));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n502), .A2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n529), .A2(KEYINPUT73), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n528), .A2(G543), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT74), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n528), .A2(new_n534), .A3(G543), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n520), .A2(G89), .A3(new_n522), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT75), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n520), .A2(new_n522), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  INV_X1    g121(.A(G651), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT76), .B(G52), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n533), .B2(new_n535), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(G171));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n520), .A2(new_n522), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(G81), .B1(new_n536), .B2(G43), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n553), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n555), .A2(new_n558), .A3(new_n553), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  XOR2_X1   g140(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n566));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G188));
  AOI22_X1  g144(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(new_n547), .ZN(new_n571));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n532), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR3_X1   g151(.A1(new_n532), .A2(KEYINPUT9), .A3(new_n573), .ZN(new_n577));
  OAI221_X1 g152(.A(new_n571), .B1(new_n545), .B2(new_n572), .C1(new_n576), .C2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  AOI21_X1  g154(.A(KEYINPUT80), .B1(new_n517), .B2(new_n524), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n517), .A2(new_n524), .A3(KEYINPUT80), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G303));
  NAND2_X1  g158(.A1(new_n554), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n528), .A2(G49), .A3(G543), .A4(new_n531), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND3_X1  g162(.A1(new_n520), .A2(G86), .A3(new_n522), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n514), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n591), .A2(KEYINPUT81), .A3(G651), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n547), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n502), .A2(G48), .A3(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n588), .A2(new_n592), .A3(new_n595), .A4(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(new_n554), .A2(G85), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(new_n547), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n536), .A2(G47), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(G290));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(G171), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT83), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OR3_X1    g183(.A1(new_n545), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n514), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n536), .A2(G54), .B1(G651), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT10), .B1(new_n545), .B2(new_n608), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n609), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n607), .B1(G868), .B2(new_n616), .ZN(G284));
  OAI21_X1  g192(.A(new_n607), .B1(G868), .B2(new_n616), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT84), .Z(new_n620));
  NOR2_X1   g195(.A1(new_n576), .A2(new_n577), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n571), .B1(new_n545), .B2(new_n572), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n620), .B1(G868), .B2(new_n623), .ZN(G297));
  OAI21_X1  g199(.A(new_n620), .B1(G868), .B2(new_n623), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n616), .B1(new_n626), .B2(G860), .ZN(G148));
  NOR2_X1   g202(.A1(new_n615), .A2(G559), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g207(.A1(new_n478), .A2(G135), .B1(G123), .B2(new_n480), .ZN(new_n633));
  NOR2_X1   g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT85), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2435), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2438), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2443), .B(G2446), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(G14), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(KEYINPUT88), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT87), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(KEYINPUT88), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT89), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n658), .B(KEYINPUT17), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n662), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(new_n662), .A3(new_n665), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n659), .A2(new_n661), .A3(new_n665), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT86), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(new_n640), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT90), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  INV_X1    g261(.A(new_n683), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n686), .B1(new_n680), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n680), .A2(KEYINPUT91), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT22), .B(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  INV_X1    g273(.A(G34), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n699), .A2(KEYINPUT24), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(KEYINPUT24), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G160), .B2(new_n698), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G2084), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G5), .A2(G16), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G171), .B2(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n478), .A2(G141), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT26), .Z(new_n711));
  NAND3_X1  g286(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n480), .A2(G129), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n709), .A2(new_n711), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT98), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT99), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G29), .B2(G32), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G1996), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n706), .B1(G1961), .B2(new_n708), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT101), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G16), .A2(G19), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n562), .B2(G16), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G1341), .Z(new_n725));
  NOR2_X1   g300(.A1(G4), .A2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n616), .B2(G16), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n727), .A2(G1348), .B1(new_n708), .B2(G1961), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n698), .A2(G35), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n698), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT104), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT29), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n725), .B(new_n728), .C1(G2090), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n718), .A2(new_n719), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n727), .A2(G1348), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT96), .B1(G29), .B2(G33), .ZN(new_n736));
  OR3_X1    g311(.A1(KEYINPUT96), .A2(G29), .A3(G33), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n478), .A2(G139), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT97), .Z(new_n739));
  NAND3_X1  g314(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT25), .Z(new_n741));
  AOI22_X1  g316(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n739), .B(new_n741), .C1(new_n461), .C2(new_n742), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n736), .B(new_n737), .C1(new_n743), .C2(new_n698), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(G2072), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(G2072), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n735), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n703), .A2(G2084), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n698), .A2(G26), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n478), .A2(G140), .B1(G128), .B2(new_n480), .ZN(new_n752));
  NOR2_X1   g327(.A1(G104), .A2(G2105), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n751), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2067), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT30), .B(G28), .Z(new_n758));
  XOR2_X1   g333(.A(KEYINPUT103), .B(G2078), .Z(new_n759));
  NOR2_X1   g334(.A1(G164), .A2(new_n698), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n698), .A2(G27), .ZN(new_n761));
  OAI21_X1  g336(.A(KEYINPUT102), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(KEYINPUT102), .B2(new_n761), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n757), .B1(G29), .B2(new_n758), .C1(new_n759), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n759), .B2(new_n763), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n734), .A2(new_n747), .A3(new_n748), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n636), .A2(new_n698), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT100), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n733), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n732), .A2(G2090), .ZN(new_n770));
  INV_X1    g345(.A(G16), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n771), .A2(KEYINPUT23), .A3(G20), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT23), .ZN(new_n773));
  INV_X1    g348(.A(G20), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(G16), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n772), .B(new_n775), .C1(new_n623), .C2(new_n771), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT105), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1956), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n770), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT106), .ZN(new_n780));
  AND3_X1   g355(.A1(new_n722), .A2(new_n769), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT31), .B(G11), .ZN(new_n782));
  NOR2_X1   g357(.A1(G166), .A2(new_n771), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n771), .B2(G22), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G23), .ZN(new_n789));
  INV_X1    g364(.A(G288), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(G16), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT33), .B(G1976), .Z(new_n792));
  XOR2_X1   g367(.A(new_n791), .B(new_n792), .Z(new_n793));
  MUX2_X1   g368(.A(G6), .B(G305), .S(G16), .Z(new_n794));
  XOR2_X1   g369(.A(KEYINPUT32), .B(G1981), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n788), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(KEYINPUT34), .ZN(new_n798));
  INV_X1    g373(.A(G290), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G16), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G16), .B2(G24), .ZN(new_n801));
  INV_X1    g376(.A(G1986), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT34), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n788), .A2(new_n793), .A3(new_n804), .A4(new_n796), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT94), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n801), .B2(new_n802), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n798), .A2(new_n803), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n478), .A2(G131), .B1(G119), .B2(new_n480), .ZN(new_n809));
  OR2_X1    g384(.A1(G95), .A2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n810), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT92), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  MUX2_X1   g388(.A(G25), .B(new_n813), .S(G29), .Z(new_n814));
  XOR2_X1   g389(.A(KEYINPUT35), .B(G1991), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT93), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n808), .A2(KEYINPUT36), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT36), .B1(new_n808), .B2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n771), .A2(G21), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G168), .B2(new_n771), .ZN(new_n822));
  INV_X1    g397(.A(G1966), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n781), .A2(new_n782), .A3(new_n820), .A4(new_n824), .ZN(G150));
  INV_X1    g400(.A(G150), .ZN(G311));
  NAND2_X1  g401(.A1(new_n536), .A2(G55), .ZN(new_n827));
  INV_X1    g402(.A(G93), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(new_n545), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n547), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n561), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n559), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT107), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT107), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n562), .A2(new_n837), .A3(new_n833), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n555), .A2(new_n558), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n832), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n836), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n615), .A2(new_n626), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n842), .B(new_n843), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n841), .B(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT108), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n833), .A2(G860), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT37), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(G145));
  XNOR2_X1  g425(.A(new_n500), .B(KEYINPUT109), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n478), .A2(G142), .B1(G130), .B2(new_n480), .ZN(new_n852));
  NOR2_X1   g427(.A1(G106), .A2(G2105), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n851), .B(new_n855), .Z(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n755), .B(new_n813), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(new_n639), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n636), .B(G160), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n484), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n861), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n743), .A2(new_n715), .ZN(new_n864));
  INV_X1    g439(.A(new_n716), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n865), .B2(new_n743), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n866), .B1(new_n862), .B2(new_n863), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n857), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n862), .A2(new_n863), .ZN(new_n871));
  INV_X1    g446(.A(new_n866), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n856), .A3(new_n867), .ZN(new_n874));
  INV_X1    g449(.A(G37), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT110), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT110), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n870), .A2(new_n874), .A3(new_n878), .A4(new_n875), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n877), .A2(KEYINPUT40), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT40), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(G395));
  XNOR2_X1  g457(.A(new_n841), .B(new_n629), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n615), .B(G299), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT41), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n884), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT42), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(G305), .B(KEYINPUT111), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n525), .ZN(new_n892));
  XNOR2_X1  g467(.A(G290), .B(G288), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n892), .B(new_n893), .Z(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n895), .A2(KEYINPUT112), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n883), .A2(new_n886), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n897), .B(new_n898), .C1(new_n883), .C2(new_n888), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n890), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n896), .B1(new_n890), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(G868), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n833), .A2(new_n605), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(G295));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n903), .ZN(G331));
  XOR2_X1   g480(.A(G171), .B(G286), .Z(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n841), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n836), .A2(new_n838), .A3(new_n840), .A4(new_n906), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n884), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n895), .B(new_n910), .C1(new_n911), .C2(new_n885), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n908), .A2(new_n884), .A3(new_n909), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n885), .B1(new_n908), .B2(new_n909), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n894), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n915), .A3(new_n875), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n912), .A2(new_n915), .A3(new_n918), .A4(new_n875), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(KEYINPUT44), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(G397));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n925));
  XOR2_X1   g500(.A(KEYINPUT113), .B(G1384), .Z(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(G164), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G160), .A2(G40), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G1996), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n716), .A2(new_n930), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n813), .A2(new_n816), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n715), .A2(G1996), .ZN(new_n933));
  INV_X1    g508(.A(G2067), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n755), .B(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n813), .A2(new_n816), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n929), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n799), .A2(new_n802), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT114), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n799), .A2(new_n802), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n929), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT115), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n938), .A2(KEYINPUT115), .A3(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT125), .ZN(new_n948));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n500), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n925), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n499), .A2(new_n496), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n493), .B1(new_n488), .B2(new_n489), .ZN(new_n953));
  AOI21_X1  g528(.A(G1384), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT45), .ZN(new_n955));
  INV_X1    g530(.A(G40), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n465), .A2(new_n468), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(G2078), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n951), .A2(new_n955), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n950), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n500), .A2(KEYINPUT50), .A3(new_n949), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n928), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n960), .B1(new_n964), .B2(G1961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT123), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT123), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n967), .B(new_n960), .C1(new_n964), .C2(G1961), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n957), .B1(new_n954), .B2(KEYINPUT45), .ZN(new_n970));
  INV_X1    g545(.A(new_n926), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT116), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n928), .B1(new_n950), .B2(new_n925), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n976), .A3(new_n972), .ZN(new_n977));
  INV_X1    g552(.A(G2078), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n958), .ZN(new_n980));
  AOI21_X1  g555(.A(G301), .B1(new_n969), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n517), .A2(KEYINPUT80), .A3(new_n524), .ZN(new_n983));
  OAI21_X1  g558(.A(G8), .B1(new_n983), .B2(new_n580), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(G303), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(G8), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n985), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(G1971), .B1(new_n974), .B2(new_n977), .ZN(new_n990));
  INV_X1    g565(.A(G2090), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n964), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n989), .B(G8), .C1(new_n990), .C2(new_n993), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n990), .B2(new_n993), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT118), .B(G86), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n520), .A2(new_n522), .A3(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n1000), .A2(new_n592), .A3(new_n595), .A4(new_n598), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1001), .A2(G1981), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G305), .A2(G1981), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n998), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n950), .A2(new_n928), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1001), .A2(G1981), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1004), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1007), .ZN(new_n1011));
  INV_X1    g586(.A(G1976), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G288), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT52), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n1012), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1015), .B(new_n1007), .C1(new_n1012), .C2(G288), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1010), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n981), .A2(new_n994), .A3(new_n997), .A4(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n950), .A2(new_n925), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n823), .B1(new_n970), .B2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g595(.A(new_n961), .B(G1384), .C1(new_n952), .C2(new_n953), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT50), .B1(new_n500), .B2(new_n949), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n705), .B(new_n957), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G286), .A2(G8), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT51), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1006), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1026), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT62), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(G286), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1030), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n948), .B1(new_n1018), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1030), .A2(new_n1037), .A3(new_n1035), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT62), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n994), .A2(new_n997), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n966), .A2(new_n968), .B1(new_n958), .B2(new_n979), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1010), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1044), .A2(new_n1045), .A3(G301), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1043), .A2(new_n1046), .A3(KEYINPUT125), .A4(new_n1038), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1040), .A2(new_n1042), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1010), .A2(new_n1012), .A3(new_n790), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1003), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1011), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1025), .B2(G286), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1033), .A2(KEYINPUT119), .A3(G168), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n997), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1017), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1051), .B1(new_n1056), .B2(KEYINPUT63), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1048), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n994), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT63), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1041), .A2(new_n994), .A3(new_n997), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n927), .A2(new_n972), .A3(new_n957), .A4(new_n959), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n957), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1067));
  INV_X1    g642(.A(G1961), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1064), .A2(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AND4_X1   g644(.A1(G301), .A2(new_n980), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1063), .B1(new_n981), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1044), .A2(G301), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n980), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(new_n1074), .A3(KEYINPUT54), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1062), .A2(new_n1071), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n970), .A2(new_n973), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT56), .B(G2072), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1956), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1067), .A2(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n571), .B(KEYINPUT120), .C1(new_n572), .C2(new_n545), .ZN(new_n1084));
  NAND3_X1  g659(.A1(G299), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1083), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n623), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1348), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1067), .A2(new_n1089), .B1(new_n934), .B2(new_n1005), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1082), .A2(new_n1088), .B1(new_n615), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1081), .A3(new_n1079), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1090), .A2(KEYINPUT60), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1005), .A2(new_n934), .ZN(new_n1096));
  OAI211_X1 g671(.A(KEYINPUT60), .B(new_n1096), .C1(new_n964), .C2(G1348), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n616), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1090), .A2(KEYINPUT60), .A3(new_n615), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1092), .A2(KEYINPUT61), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n975), .A2(new_n972), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT121), .B1(new_n1105), .B2(G1996), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1077), .A2(new_n1107), .A3(new_n930), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n950), .B2(new_n928), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(KEYINPUT59), .A3(new_n562), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT59), .B1(new_n1111), .B2(new_n562), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1094), .B1(new_n1104), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1061), .B1(new_n1076), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1017), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n947), .B1(new_n1058), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n940), .A2(new_n929), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT48), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n938), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n1123));
  OAI22_X1  g698(.A1(new_n1123), .A2(new_n932), .B1(G2067), .B2(new_n755), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n929), .ZN(new_n1125));
  INV_X1    g700(.A(new_n715), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n935), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1127), .A2(new_n929), .B1(new_n1128), .B2(KEYINPUT46), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(KEYINPUT46), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n929), .B2(new_n930), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n929), .A2(new_n930), .A3(new_n1130), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT47), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1122), .A2(new_n1125), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT127), .B1(new_n1119), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n947), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1100), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1101), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1103), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1114), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1112), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1093), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1144), .A2(new_n1071), .A3(new_n1075), .A4(new_n1062), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1045), .B1(new_n1145), .B2(new_n1061), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1048), .A2(new_n1057), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1137), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT127), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1135), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1136), .A2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g727(.A1(new_n877), .A2(new_n879), .ZN(new_n1154));
  NOR2_X1   g728(.A1(G227), .A2(G401), .ZN(new_n1155));
  INV_X1    g729(.A(G319), .ZN(new_n1156));
  NOR2_X1   g730(.A1(G229), .A2(new_n1156), .ZN(new_n1157));
  AND4_X1   g731(.A1(new_n1154), .A2(new_n920), .A3(new_n1155), .A4(new_n1157), .ZN(G308));
  NAND4_X1  g732(.A1(new_n1154), .A2(new_n920), .A3(new_n1155), .A4(new_n1157), .ZN(G225));
endmodule


