//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n575, new_n578, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n451), .A2(new_n456), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(G2104), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR3_X1   g038(.A1(new_n463), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n464));
  OAI21_X1  g039(.A(G101), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n461), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n465), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  INV_X1    g049(.A(new_n469), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  INV_X1    g051(.A(G124), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n461), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI221_X1 g056(.A(new_n476), .B1(new_n477), .B2(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT68), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(KEYINPUT70), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G138), .B1(new_n484), .B2(new_n485), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n469), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(KEYINPUT71), .B2(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n478), .A2(new_n491), .A3(new_n461), .A4(new_n486), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(new_n498), .A3(G2104), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n495), .A2(new_n494), .A3(new_n499), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n493), .B1(new_n501), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT72), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT72), .A2(G543), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n505), .B(KEYINPUT5), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT72), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT72), .A2(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT73), .B1(new_n513), .B2(KEYINPUT5), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n508), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n504), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n515), .A2(G88), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n518), .A2(new_n524), .ZN(G166));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n526), .B1(new_n519), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n519), .A2(new_n526), .A3(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n515), .A2(G89), .A3(new_n519), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XOR2_X1   g108(.A(new_n533), .B(KEYINPUT7), .Z(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n534), .B1(new_n515), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n531), .A2(new_n532), .A3(new_n536), .ZN(G168));
  INV_X1    g112(.A(new_n529), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n527), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n515), .A2(new_n519), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n504), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n504), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n515), .A2(new_n519), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n549), .A2(G81), .B1(new_n530), .B2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OR3_X1    g133(.A1(new_n521), .A2(KEYINPUT9), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n521), .B2(new_n558), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n549), .A2(G91), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n515), .A2(KEYINPUT75), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT5), .B1(new_n506), .B2(new_n507), .ZN(new_n564));
  INV_X1    g139(.A(new_n514), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(new_n567), .A3(new_n508), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n563), .A2(G65), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n562), .B1(new_n571), .B2(G651), .ZN(new_n572));
  AOI211_X1 g147(.A(KEYINPUT76), .B(new_n504), .C1(new_n569), .C2(new_n570), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n561), .B1(new_n572), .B2(new_n573), .ZN(G299));
  NAND2_X1  g149(.A1(new_n530), .A2(G52), .ZN(new_n575));
  OAI221_X1 g150(.A(new_n575), .B1(new_n542), .B2(new_n541), .C1(new_n544), .C2(new_n504), .ZN(G301));
  NAND3_X1  g151(.A1(new_n531), .A2(new_n532), .A3(new_n536), .ZN(G286));
  AOI22_X1  g152(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n520), .B(new_n523), .C1(new_n578), .C2(new_n504), .ZN(G303));
  OAI21_X1  g154(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n522), .A2(G49), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n541), .ZN(G288));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n566), .B2(new_n508), .ZN(new_n585));
  AND2_X1   g160(.A1(G73), .A2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT77), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n589), .B(G651), .C1(new_n585), .C2(new_n586), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n522), .A2(G48), .ZN(new_n592));
  INV_X1    g167(.A(G86), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n541), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n504), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n549), .A2(G85), .B1(new_n530), .B2(G47), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G290));
  NAND3_X1  g176(.A1(G301), .A2(KEYINPUT78), .A3(G868), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(G171), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n549), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n541), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n530), .A2(G54), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n563), .A2(G66), .A3(new_n568), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n504), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n602), .B(new_n605), .C1(new_n616), .C2(G868), .ZN(G284));
  XNOR2_X1  g192(.A(G284), .B(KEYINPUT79), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  XOR2_X1   g196(.A(G297), .B(KEYINPUT80), .Z(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n551), .A2(new_n604), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n613), .A2(new_n614), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n611), .B(new_n610), .C1(new_n626), .C2(new_n504), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n625), .B1(new_n628), .B2(new_n604), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g205(.A1(new_n462), .A2(new_n464), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n478), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT81), .B(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT82), .Z(new_n637));
  INV_X1    g212(.A(new_n479), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n461), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n475), .A2(new_n642), .A3(G135), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n475), .B2(G135), .ZN(new_n644));
  OAI221_X1 g219(.A(new_n639), .B1(new_n640), .B2(new_n641), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  OAI211_X1 g221(.A(new_n637), .B(new_n646), .C1(new_n635), .C2(new_n634), .ZN(G156));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n660), .A2(G14), .A3(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT84), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT17), .ZN(new_n665));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2084), .B(G2090), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n664), .B2(new_n667), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n665), .B2(new_n667), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n666), .A2(new_n668), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  OR3_X1    g249(.A1(new_n669), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(KEYINPUT85), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(KEYINPUT85), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT86), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  NAND3_X1  g265(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n692), .B(new_n695), .C1(new_n686), .C2(new_n694), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(G229));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G6), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n594), .B1(new_n588), .B2(new_n590), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT32), .B(G1981), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G23), .B(G288), .S(G16), .Z(new_n710));
  XOR2_X1   g285(.A(KEYINPUT33), .B(G1976), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT87), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n707), .A2(new_n708), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n704), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n704), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  AND4_X1   g293(.A1(new_n709), .A2(new_n713), .A3(new_n714), .A4(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G25), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n638), .A2(G119), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n475), .A2(G131), .ZN(new_n726));
  OR2_X1    g301(.A1(G95), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(new_n723), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n704), .A2(G24), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G290), .B2(G16), .ZN(new_n735));
  INV_X1    g310(.A(G1986), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n736), .B2(new_n735), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n721), .A2(new_n722), .A3(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT36), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n704), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT23), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n620), .B2(new_n704), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1956), .ZN(new_n744));
  NOR2_X1   g319(.A1(G29), .A2(G35), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G162), .B2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT100), .B(KEYINPUT29), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2090), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n638), .A2(G129), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n631), .A2(G105), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n475), .A2(G141), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT26), .Z(new_n754));
  NAND4_X1  g329(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(new_n723), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n723), .B2(G32), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT93), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  XOR2_X1   g337(.A(KEYINPUT95), .B(G28), .Z(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n766), .B1(new_n723), .B2(new_n645), .C1(new_n758), .C2(new_n759), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n723), .A2(G33), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT25), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n478), .A2(G127), .ZN(new_n771));
  NAND2_X1  g346(.A1(G115), .A2(G2104), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n461), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n770), .B(new_n773), .C1(G139), .C2(new_n475), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n768), .B1(new_n774), .B2(new_n723), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT91), .B(G2072), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n767), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n723), .A2(G26), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT28), .ZN(new_n780));
  OR2_X1    g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT90), .Z(new_n783));
  AOI22_X1  g358(.A1(new_n638), .A2(G128), .B1(G140), .B2(new_n475), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n780), .B1(new_n785), .B2(new_n723), .ZN(new_n786));
  INV_X1    g361(.A(G2067), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT24), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(G34), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(G34), .ZN(new_n791));
  AOI21_X1  g366(.A(G29), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(G160), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(G29), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT92), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G2084), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n761), .A2(new_n778), .A3(new_n788), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n704), .A2(G5), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G171), .B2(new_n704), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G1961), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT96), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n552), .A2(G16), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G16), .B2(G19), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT89), .B(G1341), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n704), .A2(G21), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G168), .B2(new_n704), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT94), .B(G1966), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n803), .A2(new_n804), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n801), .B(new_n809), .C1(new_n806), .C2(new_n808), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n803), .A2(new_n804), .B1(G1961), .B2(new_n799), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n749), .A2(new_n797), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G4), .A2(G16), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT88), .Z(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n616), .B2(G16), .ZN(new_n815));
  INV_X1    g390(.A(G1348), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n795), .A2(G2084), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n723), .A2(G27), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT98), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G164), .B2(new_n723), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G2078), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT99), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n812), .A2(new_n817), .A3(new_n819), .A4(new_n824), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n740), .A2(new_n744), .A3(new_n825), .ZN(G311));
  OR3_X1    g401(.A1(new_n740), .A2(new_n744), .A3(new_n825), .ZN(G150));
  NAND2_X1  g402(.A1(new_n515), .A2(G67), .ZN(new_n828));
  INV_X1    g403(.A(G80), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n513), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G651), .ZN(new_n831));
  OAI21_X1  g406(.A(G55), .B1(new_n538), .B2(new_n527), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n515), .A2(G93), .A3(new_n519), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n834), .B1(new_n832), .B2(new_n833), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G860), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT37), .Z(new_n840));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n552), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n832), .A2(new_n833), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT101), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n844), .A2(new_n835), .B1(G651), .B2(new_n830), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(KEYINPUT102), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n552), .A2(new_n845), .A3(KEYINPUT102), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT38), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n623), .B2(new_n627), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n849), .B(KEYINPUT38), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n627), .A2(new_n623), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n852), .A2(KEYINPUT39), .A3(new_n855), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n858), .A2(KEYINPUT103), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT103), .B1(new_n858), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n840), .B1(new_n860), .B2(new_n861), .ZN(G145));
  XNOR2_X1  g437(.A(new_n785), .B(new_n774), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n489), .A2(new_n492), .A3(new_n495), .A4(new_n499), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n863), .B(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(new_n755), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n755), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n475), .A2(G142), .ZN(new_n870));
  INV_X1    g445(.A(G130), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n461), .A2(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  OAI221_X1 g448(.A(new_n870), .B1(new_n871), .B2(new_n479), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n633), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n729), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(KEYINPUT104), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n869), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n867), .B(new_n868), .C1(KEYINPUT104), .C2(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(KEYINPUT104), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G162), .B(G160), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n645), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n876), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n885), .A2(KEYINPUT105), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n883), .B1(new_n869), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n867), .A2(new_n886), .A3(new_n868), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g467(.A(KEYINPUT108), .ZN(new_n893));
  XNOR2_X1  g468(.A(G288), .B(KEYINPUT107), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(G305), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n896));
  XNOR2_X1  g471(.A(G288), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n706), .ZN(new_n898));
  INV_X1    g473(.A(G47), .ZN(new_n899));
  INV_X1    g474(.A(G85), .ZN(new_n900));
  OAI22_X1  g475(.A1(new_n539), .A2(new_n899), .B1(new_n541), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(G166), .B1(new_n598), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n599), .A2(G303), .A3(new_n600), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n895), .A2(new_n898), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n895), .B2(new_n898), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n893), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n895), .A2(new_n898), .ZN(new_n908));
  INV_X1    g483(.A(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n895), .A2(new_n898), .A3(new_n904), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(KEYINPUT108), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT42), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n913), .A2(KEYINPUT42), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n905), .A2(new_n906), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT109), .B1(new_n917), .B2(KEYINPUT42), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n915), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n849), .B(new_n628), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n620), .A2(new_n627), .ZN(new_n921));
  NAND2_X1  g496(.A1(G299), .A2(new_n616), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n572), .A2(new_n573), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n925), .A2(KEYINPUT106), .A3(new_n561), .A4(new_n627), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(G299), .B2(new_n616), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n928), .A3(new_n922), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(G299), .B2(new_n616), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n929), .A2(new_n930), .B1(new_n921), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n924), .B1(new_n932), .B2(new_n920), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n919), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n919), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(G868), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(G868), .B2(new_n845), .ZN(G295));
  OAI21_X1  g512(.A(new_n936), .B1(G868), .B2(new_n845), .ZN(G331));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(G301), .B2(G168), .ZN(new_n941));
  NAND3_X1  g516(.A1(G171), .A2(KEYINPUT111), .A3(G286), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(G171), .B2(G286), .ZN(new_n945));
  NAND3_X1  g520(.A1(G301), .A2(KEYINPUT110), .A3(G168), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n847), .B2(new_n848), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n842), .A2(new_n846), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n845), .A2(KEYINPUT102), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n838), .A2(new_n841), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n552), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n950), .A2(new_n953), .A3(new_n947), .A4(new_n943), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n932), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n923), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n913), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n957), .B(new_n913), .C1(new_n932), .C2(new_n955), .ZN(new_n959));
  INV_X1    g534(.A(G37), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n939), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n923), .A2(new_n930), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n926), .A2(new_n928), .A3(new_n931), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n949), .A2(new_n954), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n913), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n957), .A2(KEYINPUT112), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n955), .B1(new_n963), .B2(new_n964), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n968), .B(new_n969), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n972), .A2(KEYINPUT43), .A3(new_n960), .A4(new_n959), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n962), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT44), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT43), .B1(new_n958), .B2(new_n961), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n972), .A2(new_n939), .A3(new_n960), .A4(new_n959), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(new_n980), .ZN(G397));
  OAI21_X1  g556(.A(G8), .B1(KEYINPUT121), .B2(KEYINPUT51), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G1384), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT116), .B1(G164), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n473), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n475), .A2(G137), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n988), .A3(G40), .A4(new_n465), .ZN(new_n989));
  INV_X1    g564(.A(G1384), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n864), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n989), .B1(new_n991), .B2(new_n983), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n495), .A2(new_n494), .A3(new_n499), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n489), .B(new_n492), .C1(new_n993), .C2(new_n500), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(new_n995), .A3(new_n984), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n986), .A2(new_n992), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n994), .B2(new_n990), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n864), .A2(new_n998), .A3(new_n990), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n470), .A2(new_n1001), .A3(new_n473), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G2084), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n997), .A2(new_n807), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n982), .B1(new_n1006), .B2(G168), .ZN(new_n1007));
  NAND2_X1  g582(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n991), .A2(new_n983), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n996), .A2(new_n1010), .A3(new_n1002), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n995), .B1(new_n994), .B2(new_n984), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n807), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1007), .A2(new_n1008), .B1(G286), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(G168), .A3(new_n1014), .ZN(new_n1017));
  INV_X1    g592(.A(new_n982), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1008), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT122), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(new_n1018), .A3(new_n1008), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(G8), .A3(G286), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT122), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n1019), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT62), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1016), .A2(new_n1020), .A3(KEYINPUT122), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1026), .B1(new_n1025), .B2(new_n1019), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT62), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n983), .B1(G164), .B2(G1384), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n864), .A2(new_n984), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n1002), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1033), .B1(new_n1036), .B2(G2078), .ZN(new_n1037));
  INV_X1    g612(.A(G1961), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n999), .B2(new_n1003), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1033), .A2(G2078), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n986), .A2(new_n992), .A3(new_n996), .A4(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G171), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT123), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n991), .A2(new_n989), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(new_n1009), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G288), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT52), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1049), .B(new_n1054), .C1(new_n1051), .C2(G288), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT49), .ZN(new_n1057));
  AOI211_X1 g632(.A(G1981), .B(new_n594), .C1(new_n588), .C2(new_n590), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n595), .B2(new_n587), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1057), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n595), .A2(new_n587), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(G1981), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1064), .A3(new_n1049), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1066));
  INV_X1    g641(.A(G2090), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n1002), .A4(new_n1000), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT45), .B1(new_n994), .B2(new_n990), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1002), .A2(new_n1035), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n717), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1009), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT55), .B(G8), .C1(new_n518), .C2(new_n524), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT114), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(G166), .B2(new_n1009), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n1077));
  NAND4_X1  g652(.A1(G303), .A2(new_n1077), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1074), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1072), .A2(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1056), .A2(new_n1065), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n989), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n994), .A2(new_n998), .A3(new_n990), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1067), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1009), .B1(new_n1071), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n1086));
  OR3_X1    g661(.A1(new_n1085), .A2(new_n1079), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1085), .B2(new_n1079), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1047), .A2(new_n1081), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1028), .A2(new_n1032), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1028), .A2(new_n1090), .A3(KEYINPUT125), .A4(new_n1032), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1048), .A2(new_n787), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n816), .B1(new_n999), .B2(new_n1003), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n627), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(new_n561), .C1(new_n572), .C2(new_n573), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT56), .B(G2072), .Z(new_n1101));
  NOR3_X1   g676(.A1(new_n1069), .A2(new_n1070), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1956), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1098), .A2(new_n1100), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1096), .A2(new_n1095), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n616), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1097), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(KEYINPUT120), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1105), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1069), .A2(new_n1070), .A3(G1996), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT58), .B(G1341), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1048), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n552), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(KEYINPUT59), .B(new_n552), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n616), .A2(new_n1122), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(KEYINPUT61), .B2(new_n1105), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1112), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1109), .B(new_n1114), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1103), .B2(new_n1102), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT53), .B1(KEYINPUT124), .B2(G2078), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(KEYINPUT124), .B2(G2078), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n992), .A2(new_n1035), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1037), .A2(new_n1039), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(G171), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1037), .A2(G301), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(KEYINPUT54), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1081), .A2(new_n1138), .A3(new_n1089), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1045), .B(new_n1046), .C1(G171), .C2(new_n1135), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1130), .A2(new_n1131), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(G288), .A2(G1976), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1058), .B1(new_n1065), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1056), .A2(new_n1065), .ZN(new_n1146));
  OAI22_X1  g721(.A1(new_n1145), .A2(new_n1050), .B1(new_n1146), .B2(new_n1080), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1072), .A2(new_n1148), .ZN(new_n1149));
  AOI211_X1 g724(.A(KEYINPUT118), .B(new_n1009), .C1(new_n1068), .C2(new_n1071), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1074), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1015), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1081), .A2(new_n1153), .A3(KEYINPUT119), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1006), .A2(new_n1009), .A3(G286), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1152), .B1(new_n1072), .B2(new_n1148), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1157), .B(KEYINPUT63), .C1(new_n1158), .C2(new_n1150), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1056), .A2(new_n1065), .A3(new_n1080), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1156), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1155), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1081), .A2(new_n1089), .A3(new_n1157), .ZN(new_n1163));
  XOR2_X1   g738(.A(KEYINPUT117), .B(KEYINPUT63), .Z(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1147), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1093), .A2(new_n1094), .A3(new_n1143), .A4(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(G290), .A2(G1986), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(G290), .A2(G1986), .ZN(new_n1170));
  OR3_X1    g745(.A1(new_n1169), .A2(KEYINPUT113), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1010), .A2(new_n989), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1169), .B2(KEYINPUT113), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n785), .B(G2067), .ZN(new_n1175));
  INV_X1    g750(.A(G1996), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n755), .B(new_n1176), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n730), .A2(new_n732), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n730), .A2(new_n732), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1171), .A2(new_n1174), .B1(new_n1172), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1167), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT48), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1170), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT48), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1184), .A2(new_n1185), .A3(new_n1173), .ZN(new_n1186));
  AOI211_X1 g761(.A(new_n1183), .B(new_n1186), .C1(new_n1172), .C2(new_n1180), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT46), .Z(new_n1189));
  AOI21_X1  g764(.A(new_n1173), .B1(new_n1175), .B2(new_n756), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT47), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n785), .A2(new_n787), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1193), .B1(new_n1194), .B2(new_n1179), .ZN(new_n1195));
  AOI211_X1 g770(.A(new_n1187), .B(new_n1192), .C1(new_n1172), .C2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1182), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g772(.A1(new_n681), .A2(G319), .A3(new_n682), .ZN(new_n1199));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g775(.A1(new_n681), .A2(KEYINPUT126), .A3(G319), .A4(new_n682), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g777(.A(G401), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1205), .A2(KEYINPUT127), .ZN(new_n1206));
  AOI21_X1  g780(.A(G229), .B1(new_n884), .B2(new_n890), .ZN(new_n1207));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n1208));
  NAND3_X1  g782(.A1(new_n1203), .A2(new_n1208), .A3(new_n1204), .ZN(new_n1209));
  AND4_X1   g783(.A1(new_n978), .A2(new_n1206), .A3(new_n1207), .A4(new_n1209), .ZN(G308));
  NAND4_X1  g784(.A1(new_n978), .A2(new_n1206), .A3(new_n1207), .A4(new_n1209), .ZN(G225));
endmodule


