

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727;

  XNOR2_X1 U363 ( .A(n557), .B(KEYINPUT85), .ZN(n573) );
  AND2_X1 U364 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X2 U365 ( .A(n353), .B(n348), .ZN(n506) );
  NOR2_X2 U366 ( .A1(n625), .A2(n563), .ZN(n537) );
  XNOR2_X2 U367 ( .A(n531), .B(n530), .ZN(n625) );
  XNOR2_X2 U368 ( .A(G478), .B(n342), .ZN(n511) );
  INV_X1 U369 ( .A(n528), .ZN(n603) );
  XNOR2_X1 U370 ( .A(G143), .B(KEYINPUT65), .ZN(n404) );
  NOR2_X1 U371 ( .A1(n548), .A2(n505), .ZN(n673) );
  XNOR2_X1 U372 ( .A(n553), .B(n552), .ZN(n639) );
  AND2_X1 U373 ( .A1(n570), .A2(n393), .ZN(n553) );
  XNOR2_X1 U374 ( .A(n495), .B(n363), .ZN(n727) );
  NAND2_X1 U375 ( .A1(n396), .A2(n346), .ZN(n395) );
  XNOR2_X1 U376 ( .A(n716), .B(n427), .ZN(n475) );
  XNOR2_X1 U377 ( .A(n404), .B(G128), .ZN(n476) );
  XNOR2_X1 U378 ( .A(n426), .B(G146), .ZN(n716) );
  XNOR2_X1 U379 ( .A(n439), .B(G110), .ZN(n483) );
  INV_X1 U380 ( .A(G119), .ZN(n439) );
  XNOR2_X1 U381 ( .A(G113), .B(G104), .ZN(n418) );
  XNOR2_X1 U382 ( .A(n365), .B(n364), .ZN(n614) );
  INV_X1 U383 ( .A(KEYINPUT41), .ZN(n364) );
  NOR2_X1 U384 ( .A1(n619), .A2(n618), .ZN(n365) );
  INV_X1 U385 ( .A(n725), .ZN(n356) );
  INV_X1 U386 ( .A(n727), .ZN(n355) );
  XNOR2_X1 U387 ( .A(n425), .B(n397), .ZN(n712) );
  XOR2_X1 U388 ( .A(G137), .B(G131), .Z(n397) );
  INV_X1 U389 ( .A(KEYINPUT4), .ZN(n426) );
  XNOR2_X1 U390 ( .A(n386), .B(KEYINPUT70), .ZN(n602) );
  OR2_X1 U391 ( .A1(n554), .A2(n598), .ZN(n386) );
  OR2_X1 U392 ( .A1(n676), .A2(G902), .ZN(n377) );
  XNOR2_X1 U393 ( .A(n712), .B(n475), .ZN(n467) );
  XOR2_X1 U394 ( .A(G119), .B(G116), .Z(n463) );
  XNOR2_X1 U395 ( .A(KEYINPUT3), .B(G113), .ZN(n462) );
  NAND2_X1 U396 ( .A1(n391), .A2(n580), .ZN(n388) );
  XNOR2_X1 U397 ( .A(KEYINPUT18), .B(G125), .ZN(n477) );
  XNOR2_X1 U398 ( .A(n384), .B(n383), .ZN(n523) );
  INV_X1 U399 ( .A(KEYINPUT39), .ZN(n383) );
  AND2_X1 U400 ( .A1(n474), .A2(n345), .ZN(n382) );
  XNOR2_X1 U401 ( .A(n603), .B(n394), .ZN(n548) );
  INV_X1 U402 ( .A(KEYINPUT87), .ZN(n394) );
  NAND2_X1 U403 ( .A1(n585), .A2(n580), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n488), .B(n487), .ZN(n705) );
  NOR2_X1 U405 ( .A1(n633), .A2(n344), .ZN(n369) );
  INV_X1 U406 ( .A(n597), .ZN(n367) );
  XNOR2_X1 U407 ( .A(n381), .B(n380), .ZN(n714) );
  INV_X1 U408 ( .A(KEYINPUT10), .ZN(n380) );
  XNOR2_X1 U409 ( .A(G140), .B(G125), .ZN(n381) );
  NOR2_X1 U410 ( .A1(n583), .A2(n350), .ZN(n390) );
  XOR2_X1 U411 ( .A(G140), .B(G110), .Z(n429) );
  NAND2_X1 U412 ( .A1(n345), .A2(n616), .ZN(n619) );
  XNOR2_X1 U413 ( .A(n423), .B(n422), .ZN(n510) );
  XNOR2_X1 U414 ( .A(n421), .B(G475), .ZN(n422) );
  XNOR2_X1 U415 ( .A(n520), .B(KEYINPUT72), .ZN(n521) );
  XOR2_X1 U416 ( .A(KEYINPUT92), .B(KEYINPUT75), .Z(n442) );
  XNOR2_X1 U417 ( .A(G137), .B(G128), .ZN(n441) );
  XNOR2_X1 U418 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n438) );
  XOR2_X1 U419 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n407) );
  XNOR2_X1 U420 ( .A(n476), .B(n405), .ZN(n425) );
  XNOR2_X1 U421 ( .A(n714), .B(G146), .ZN(n436) );
  XNOR2_X1 U422 ( .A(n467), .B(n378), .ZN(n676) );
  XNOR2_X1 U423 ( .A(n431), .B(G104), .ZN(n378) );
  XNOR2_X1 U424 ( .A(n430), .B(n398), .ZN(n431) );
  XNOR2_X1 U425 ( .A(KEYINPUT78), .B(G107), .ZN(n398) );
  NOR2_X1 U426 ( .A1(n548), .A2(n547), .ZN(n393) );
  NAND2_X1 U427 ( .A1(n528), .A2(n347), .ZN(n611) );
  XNOR2_X1 U428 ( .A(n448), .B(n387), .ZN(n554) );
  XNOR2_X1 U429 ( .A(n340), .B(n451), .ZN(n387) );
  NOR2_X1 U430 ( .A1(n691), .A2(G902), .ZN(n448) );
  XNOR2_X1 U431 ( .A(n452), .B(n385), .ZN(n562) );
  NOR2_X1 U432 ( .A1(n498), .A2(n602), .ZN(n452) );
  XNOR2_X1 U433 ( .A(n467), .B(n466), .ZN(n641) );
  INV_X1 U434 ( .A(G475), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n705), .B(n354), .ZN(n585) );
  XNOR2_X1 U436 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n363) );
  NAND2_X1 U437 ( .A1(n360), .A2(n357), .ZN(n725) );
  NAND2_X1 U438 ( .A1(n359), .A2(n358), .ZN(n357) );
  XNOR2_X1 U439 ( .A(KEYINPUT35), .B(KEYINPUT83), .ZN(n541) );
  XNOR2_X1 U440 ( .A(n379), .B(KEYINPUT31), .ZN(n670) );
  NOR2_X1 U441 ( .A1(n611), .A2(n563), .ZN(n379) );
  NAND2_X1 U442 ( .A1(n506), .A2(n616), .ZN(n507) );
  XNOR2_X1 U443 ( .A(n691), .B(n692), .ZN(n693) );
  AND2_X1 U444 ( .A1(n369), .A2(n366), .ZN(n636) );
  OR2_X1 U445 ( .A1(n595), .A2(KEYINPUT2), .ZN(n339) );
  INV_X1 U446 ( .A(n583), .ZN(n391) );
  AND2_X1 U447 ( .A1(G217), .A2(n447), .ZN(n340) );
  XOR2_X1 U448 ( .A(KEYINPUT74), .B(G469), .Z(n341) );
  OR2_X1 U449 ( .A1(G902), .A2(n687), .ZN(n342) );
  XOR2_X1 U450 ( .A(KEYINPUT23), .B(KEYINPUT91), .Z(n343) );
  OR2_X1 U451 ( .A1(G953), .A2(n593), .ZN(n344) );
  XNOR2_X1 U452 ( .A(KEYINPUT38), .B(n526), .ZN(n345) );
  NOR2_X1 U453 ( .A1(n618), .A2(n598), .ZN(n346) );
  BUF_X1 U454 ( .A(n549), .Z(n563) );
  AND2_X1 U455 ( .A1(n560), .A2(n607), .ZN(n347) );
  AND2_X1 U456 ( .A1(n489), .A2(G210), .ZN(n348) );
  XOR2_X1 U457 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n349) );
  NOR2_X1 U458 ( .A1(n596), .A2(KEYINPUT67), .ZN(n350) );
  OR2_X1 U459 ( .A1(n596), .A2(KEYINPUT81), .ZN(n351) );
  XNOR2_X2 U460 ( .A(n352), .B(KEYINPUT45), .ZN(n697) );
  NAND2_X2 U461 ( .A1(n578), .A2(n577), .ZN(n352) );
  XNOR2_X2 U462 ( .A(n468), .B(n469), .ZN(n607) );
  NOR2_X1 U463 ( .A1(n589), .A2(n696), .ZN(n590) );
  NOR2_X1 U464 ( .A1(n685), .A2(n696), .ZN(n686) );
  XNOR2_X1 U465 ( .A(n481), .B(n480), .ZN(n354) );
  NAND2_X1 U466 ( .A1(n523), .A2(n349), .ZN(n362) );
  NAND2_X1 U467 ( .A1(n356), .A2(n355), .ZN(n496) );
  NOR2_X1 U468 ( .A1(n667), .A2(n349), .ZN(n358) );
  INV_X1 U469 ( .A(n523), .ZN(n359) );
  AND2_X1 U470 ( .A1(n362), .A2(n361), .ZN(n360) );
  NAND2_X1 U471 ( .A1(n667), .A2(n349), .ZN(n361) );
  NAND2_X1 U472 ( .A1(n368), .A2(n367), .ZN(n366) );
  NAND2_X1 U473 ( .A1(n339), .A2(n351), .ZN(n368) );
  NOR2_X1 U474 ( .A1(n584), .A2(n597), .ZN(n690) );
  NAND2_X1 U475 ( .A1(n370), .A2(n373), .ZN(n643) );
  NOR2_X1 U476 ( .A1(n597), .A2(n371), .ZN(n370) );
  INV_X1 U477 ( .A(G472), .ZN(n371) );
  NAND2_X1 U478 ( .A1(n372), .A2(n373), .ZN(n684) );
  NOR2_X1 U479 ( .A1(n597), .A2(n375), .ZN(n372) );
  NAND2_X1 U480 ( .A1(n374), .A2(n373), .ZN(n588) );
  INV_X1 U481 ( .A(n584), .ZN(n373) );
  NOR2_X1 U482 ( .A1(n597), .A2(n376), .ZN(n374) );
  INV_X1 U483 ( .A(G210), .ZN(n376) );
  XNOR2_X2 U484 ( .A(n377), .B(n341), .ZN(n498) );
  NAND2_X1 U485 ( .A1(n392), .A2(n390), .ZN(n389) );
  NAND2_X1 U486 ( .A1(n389), .A2(n388), .ZN(n584) );
  XNOR2_X2 U487 ( .A(n498), .B(n497), .ZN(n528) );
  INV_X1 U488 ( .A(n392), .ZN(n594) );
  NOR2_X2 U489 ( .A1(n392), .A2(n596), .ZN(n597) );
  NAND2_X1 U490 ( .A1(n562), .A2(n474), .ZN(n513) );
  NAND2_X1 U491 ( .A1(n562), .A2(n382), .ZN(n384) );
  INV_X1 U492 ( .A(KEYINPUT95), .ZN(n385) );
  NAND2_X1 U493 ( .A1(n579), .A2(n697), .ZN(n392) );
  XNOR2_X2 U494 ( .A(n395), .B(n550), .ZN(n570) );
  INV_X1 U495 ( .A(n549), .ZN(n396) );
  INV_X1 U496 ( .A(n506), .ZN(n526) );
  XNOR2_X2 U497 ( .A(n507), .B(KEYINPUT19), .ZN(n659) );
  XNOR2_X1 U498 ( .A(n496), .B(KEYINPUT46), .ZN(n519) );
  NAND2_X1 U499 ( .A1(n529), .A2(n528), .ZN(n531) );
  INV_X1 U500 ( .A(G134), .ZN(n405) );
  INV_X1 U501 ( .A(KEYINPUT125), .ZN(n692) );
  OR2_X1 U502 ( .A1(n718), .A2(G952), .ZN(n644) );
  XNOR2_X1 U503 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U504 ( .A(n636), .B(n635), .ZN(G75) );
  XNOR2_X1 U505 ( .A(G116), .B(G107), .ZN(n482) );
  INV_X1 U506 ( .A(KEYINPUT64), .ZN(n399) );
  XNOR2_X2 U507 ( .A(n399), .B(G953), .ZN(n718) );
  NAND2_X1 U508 ( .A1(n718), .A2(G234), .ZN(n402) );
  XNOR2_X1 U509 ( .A(KEYINPUT8), .B(KEYINPUT71), .ZN(n400) );
  XNOR2_X1 U510 ( .A(n400), .B(KEYINPUT82), .ZN(n401) );
  XNOR2_X1 U511 ( .A(n402), .B(n401), .ZN(n435) );
  NAND2_X1 U512 ( .A1(G217), .A2(n435), .ZN(n403) );
  XOR2_X1 U513 ( .A(n482), .B(n403), .Z(n411) );
  XNOR2_X1 U514 ( .A(G122), .B(KEYINPUT9), .ZN(n406) );
  XNOR2_X1 U515 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U516 ( .A(n408), .B(KEYINPUT104), .Z(n409) );
  XNOR2_X1 U517 ( .A(n425), .B(n409), .ZN(n410) );
  XNOR2_X1 U518 ( .A(n411), .B(n410), .ZN(n687) );
  XOR2_X1 U519 ( .A(G131), .B(KEYINPUT99), .Z(n413) );
  NOR2_X1 U520 ( .A1(G953), .A2(G237), .ZN(n459) );
  NAND2_X1 U521 ( .A1(G214), .A2(n459), .ZN(n412) );
  XNOR2_X1 U522 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U523 ( .A(KEYINPUT100), .B(KEYINPUT11), .Z(n415) );
  XNOR2_X1 U524 ( .A(G143), .B(KEYINPUT12), .ZN(n414) );
  XNOR2_X1 U525 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U526 ( .A(n417), .B(n416), .Z(n420) );
  XNOR2_X1 U527 ( .A(n418), .B(G122), .ZN(n487) );
  XNOR2_X1 U528 ( .A(n436), .B(n487), .ZN(n419) );
  XNOR2_X1 U529 ( .A(n420), .B(n419), .ZN(n682) );
  NOR2_X1 U530 ( .A1(G902), .A2(n682), .ZN(n423) );
  XNOR2_X1 U531 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n421) );
  XNOR2_X1 U532 ( .A(KEYINPUT102), .B(n510), .ZN(n508) );
  NOR2_X1 U533 ( .A1(n511), .A2(n508), .ZN(n424) );
  XNOR2_X2 U534 ( .A(KEYINPUT105), .B(n424), .ZN(n667) );
  XNOR2_X1 U535 ( .A(KEYINPUT68), .B(G101), .ZN(n427) );
  NAND2_X1 U536 ( .A1(G227), .A2(n718), .ZN(n428) );
  XNOR2_X1 U537 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U538 ( .A(G902), .B(KEYINPUT15), .ZN(n580) );
  NAND2_X1 U539 ( .A1(n580), .A2(G234), .ZN(n432) );
  XNOR2_X1 U540 ( .A(n432), .B(KEYINPUT20), .ZN(n447) );
  AND2_X1 U541 ( .A1(n447), .A2(G221), .ZN(n434) );
  INV_X1 U542 ( .A(KEYINPUT21), .ZN(n433) );
  XNOR2_X1 U543 ( .A(n434), .B(n433), .ZN(n598) );
  NAND2_X1 U544 ( .A1(G221), .A2(n435), .ZN(n437) );
  XNOR2_X1 U545 ( .A(n437), .B(n436), .ZN(n446) );
  XNOR2_X1 U546 ( .A(n343), .B(n438), .ZN(n440) );
  XNOR2_X1 U547 ( .A(n440), .B(n483), .ZN(n444) );
  XNOR2_X1 U548 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U549 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U550 ( .A(n446), .B(n445), .ZN(n691) );
  XOR2_X1 U551 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n450) );
  XNOR2_X1 U552 ( .A(KEYINPUT93), .B(KEYINPUT77), .ZN(n449) );
  XOR2_X1 U553 ( .A(n450), .B(n449), .Z(n451) );
  NAND2_X1 U554 ( .A1(G234), .A2(G237), .ZN(n453) );
  XNOR2_X1 U555 ( .A(n453), .B(KEYINPUT88), .ZN(n454) );
  XNOR2_X1 U556 ( .A(KEYINPUT14), .B(n454), .ZN(n455) );
  NAND2_X1 U557 ( .A1(G952), .A2(n455), .ZN(n631) );
  NOR2_X1 U558 ( .A1(n631), .A2(G953), .ZN(n534) );
  NAND2_X1 U559 ( .A1(G902), .A2(n455), .ZN(n532) );
  NOR2_X1 U560 ( .A1(n718), .A2(n532), .ZN(n456) );
  XNOR2_X1 U561 ( .A(n456), .B(KEYINPUT107), .ZN(n457) );
  NOR2_X1 U562 ( .A1(G900), .A2(n457), .ZN(n458) );
  NOR2_X1 U563 ( .A1(n534), .A2(n458), .ZN(n490) );
  XNOR2_X1 U564 ( .A(G472), .B(KEYINPUT97), .ZN(n469) );
  XOR2_X1 U565 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n461) );
  NAND2_X1 U566 ( .A1(n459), .A2(G210), .ZN(n460) );
  XNOR2_X1 U567 ( .A(n461), .B(n460), .ZN(n465) );
  XNOR2_X1 U568 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U569 ( .A(n465), .B(n464), .ZN(n466) );
  NOR2_X1 U570 ( .A1(n641), .A2(G902), .ZN(n468) );
  INV_X1 U571 ( .A(G902), .ZN(n471) );
  INV_X1 U572 ( .A(G237), .ZN(n470) );
  NAND2_X1 U573 ( .A1(n471), .A2(n470), .ZN(n489) );
  NAND2_X1 U574 ( .A1(n489), .A2(G214), .ZN(n616) );
  NAND2_X1 U575 ( .A1(n607), .A2(n616), .ZN(n472) );
  XNOR2_X1 U576 ( .A(KEYINPUT30), .B(n472), .ZN(n473) );
  NOR2_X1 U577 ( .A1(n490), .A2(n473), .ZN(n474) );
  XNOR2_X1 U578 ( .A(n476), .B(n475), .ZN(n481) );
  NAND2_X1 U579 ( .A1(n718), .A2(G224), .ZN(n479) );
  XNOR2_X1 U580 ( .A(n477), .B(KEYINPUT17), .ZN(n478) );
  XNOR2_X1 U581 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U582 ( .A(n483), .B(n482), .ZN(n486) );
  XNOR2_X1 U583 ( .A(KEYINPUT76), .B(KEYINPUT3), .ZN(n484) );
  XNOR2_X1 U584 ( .A(n484), .B(KEYINPUT16), .ZN(n485) );
  XNOR2_X1 U585 ( .A(n486), .B(n485), .ZN(n488) );
  INV_X1 U586 ( .A(n607), .ZN(n561) );
  NOR2_X1 U587 ( .A1(n490), .A2(n598), .ZN(n491) );
  NAND2_X1 U588 ( .A1(n491), .A2(n554), .ZN(n502) );
  NOR2_X1 U589 ( .A1(n561), .A2(n502), .ZN(n492) );
  XOR2_X1 U590 ( .A(KEYINPUT28), .B(n492), .Z(n493) );
  NOR2_X1 U591 ( .A1(n498), .A2(n493), .ZN(n658) );
  INV_X1 U592 ( .A(n511), .ZN(n494) );
  NAND2_X1 U593 ( .A1(n510), .A2(n494), .ZN(n618) );
  NAND2_X1 U594 ( .A1(n658), .A2(n614), .ZN(n495) );
  INV_X1 U595 ( .A(KEYINPUT1), .ZN(n497) );
  INV_X1 U596 ( .A(n667), .ZN(n500) );
  INV_X1 U597 ( .A(KEYINPUT6), .ZN(n499) );
  XNOR2_X1 U598 ( .A(n607), .B(n499), .ZN(n568) );
  NAND2_X1 U599 ( .A1(n500), .A2(n568), .ZN(n501) );
  NOR2_X1 U600 ( .A1(n502), .A2(n501), .ZN(n503) );
  NAND2_X1 U601 ( .A1(n503), .A2(n616), .ZN(n524) );
  NOR2_X1 U602 ( .A1(n524), .A2(n526), .ZN(n504) );
  XOR2_X1 U603 ( .A(KEYINPUT36), .B(n504), .Z(n505) );
  NAND2_X1 U604 ( .A1(n658), .A2(n659), .ZN(n664) );
  NAND2_X1 U605 ( .A1(n508), .A2(n511), .ZN(n671) );
  AND2_X1 U606 ( .A1(n667), .A2(n671), .ZN(n620) );
  NOR2_X1 U607 ( .A1(n664), .A2(n620), .ZN(n509) );
  XNOR2_X1 U608 ( .A(n509), .B(KEYINPUT47), .ZN(n515) );
  INV_X1 U609 ( .A(n510), .ZN(n512) );
  NAND2_X1 U610 ( .A1(n512), .A2(n511), .ZN(n538) );
  NOR2_X1 U611 ( .A1(n513), .A2(n538), .ZN(n514) );
  NAND2_X1 U612 ( .A1(n514), .A2(n506), .ZN(n637) );
  NAND2_X1 U613 ( .A1(n515), .A2(n637), .ZN(n516) );
  NOR2_X1 U614 ( .A1(n673), .A2(n516), .ZN(n517) );
  XNOR2_X1 U615 ( .A(KEYINPUT73), .B(n517), .ZN(n518) );
  NOR2_X1 U616 ( .A1(n519), .A2(n518), .ZN(n522) );
  INV_X1 U617 ( .A(KEYINPUT48), .ZN(n520) );
  XNOR2_X1 U618 ( .A(n522), .B(n521), .ZN(n711) );
  NOR2_X1 U619 ( .A1(n523), .A2(n671), .ZN(n675) );
  OR2_X1 U620 ( .A1(n524), .A2(n528), .ZN(n525) );
  XNOR2_X1 U621 ( .A(n525), .B(KEYINPUT43), .ZN(n527) );
  AND2_X1 U622 ( .A1(n527), .A2(n526), .ZN(n638) );
  OR2_X1 U623 ( .A1(n675), .A2(n638), .ZN(n710) );
  NOR2_X1 U624 ( .A1(n711), .A2(n710), .ZN(n579) );
  INV_X1 U625 ( .A(n602), .ZN(n560) );
  AND2_X1 U626 ( .A1(n560), .A2(n568), .ZN(n529) );
  XOR2_X1 U627 ( .A(KEYINPUT86), .B(KEYINPUT33), .Z(n530) );
  XNOR2_X1 U628 ( .A(G898), .B(KEYINPUT89), .ZN(n701) );
  NAND2_X1 U629 ( .A1(G953), .A2(n701), .ZN(n706) );
  NOR2_X1 U630 ( .A1(n532), .A2(n706), .ZN(n533) );
  OR2_X1 U631 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U632 ( .A1(n659), .A2(n535), .ZN(n536) );
  XNOR2_X1 U633 ( .A(n536), .B(KEYINPUT0), .ZN(n549) );
  XNOR2_X1 U634 ( .A(n537), .B(KEYINPUT34), .ZN(n540) );
  INV_X1 U635 ( .A(n538), .ZN(n539) );
  NAND2_X1 U636 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X2 U637 ( .A(n542), .B(n541), .ZN(n726) );
  INV_X1 U638 ( .A(KEYINPUT44), .ZN(n543) );
  NAND2_X1 U639 ( .A1(n726), .A2(n543), .ZN(n544) );
  XNOR2_X1 U640 ( .A(n544), .B(KEYINPUT69), .ZN(n559) );
  INV_X1 U641 ( .A(KEYINPUT80), .ZN(n545) );
  XNOR2_X1 U642 ( .A(n568), .B(n545), .ZN(n546) );
  XNOR2_X1 U643 ( .A(n554), .B(KEYINPUT106), .ZN(n599) );
  NAND2_X1 U644 ( .A1(n546), .A2(n599), .ZN(n547) );
  INV_X1 U645 ( .A(KEYINPUT22), .ZN(n550) );
  XNOR2_X1 U646 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n551) );
  XNOR2_X1 U647 ( .A(n551), .B(KEYINPUT66), .ZN(n552) );
  NAND2_X1 U648 ( .A1(n561), .A2(n554), .ZN(n555) );
  NOR2_X1 U649 ( .A1(n528), .A2(n555), .ZN(n556) );
  NAND2_X1 U650 ( .A1(n556), .A2(n570), .ZN(n656) );
  NAND2_X1 U651 ( .A1(n639), .A2(n656), .ZN(n557) );
  XNOR2_X1 U652 ( .A(n573), .B(KEYINPUT84), .ZN(n558) );
  NAND2_X1 U653 ( .A1(n559), .A2(n558), .ZN(n578) );
  AND2_X1 U654 ( .A1(n562), .A2(n561), .ZN(n564) );
  NAND2_X1 U655 ( .A1(n564), .A2(n396), .ZN(n651) );
  NAND2_X1 U656 ( .A1(n670), .A2(n651), .ZN(n565) );
  XNOR2_X1 U657 ( .A(n565), .B(KEYINPUT98), .ZN(n567) );
  INV_X1 U658 ( .A(n620), .ZN(n566) );
  NAND2_X1 U659 ( .A1(n567), .A2(n566), .ZN(n572) );
  OR2_X1 U660 ( .A1(n568), .A2(n599), .ZN(n569) );
  NOR2_X1 U661 ( .A1(n528), .A2(n569), .ZN(n571) );
  NAND2_X1 U662 ( .A1(n571), .A2(n570), .ZN(n647) );
  AND2_X1 U663 ( .A1(n572), .A2(n647), .ZN(n576) );
  NAND2_X1 U664 ( .A1(n726), .A2(n573), .ZN(n574) );
  NAND2_X1 U665 ( .A1(n574), .A2(KEYINPUT44), .ZN(n575) );
  INV_X1 U666 ( .A(KEYINPUT2), .ZN(n596) );
  INV_X1 U667 ( .A(n580), .ZN(n581) );
  NAND2_X1 U668 ( .A1(n581), .A2(KEYINPUT2), .ZN(n582) );
  AND2_X1 U669 ( .A1(n582), .A2(KEYINPUT67), .ZN(n583) );
  XOR2_X1 U670 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n586) );
  XOR2_X1 U671 ( .A(n586), .B(n585), .Z(n587) );
  XNOR2_X1 U672 ( .A(n588), .B(n587), .ZN(n589) );
  INV_X1 U673 ( .A(n644), .ZN(n696) );
  XNOR2_X1 U674 ( .A(n590), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U675 ( .A(n625), .ZN(n591) );
  NAND2_X1 U676 ( .A1(n614), .A2(n591), .ZN(n592) );
  XOR2_X1 U677 ( .A(KEYINPUT122), .B(n592), .Z(n593) );
  NOR2_X1 U678 ( .A1(n594), .A2(KEYINPUT81), .ZN(n595) );
  XOR2_X1 U679 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n601) );
  NAND2_X1 U680 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U681 ( .A(n601), .B(n600), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U683 ( .A(n604), .B(KEYINPUT50), .ZN(n605) );
  XNOR2_X1 U684 ( .A(KEYINPUT117), .B(n605), .ZN(n606) );
  NOR2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U688 ( .A(KEYINPUT51), .B(n612), .Z(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U690 ( .A(KEYINPUT118), .B(n615), .Z(n627) );
  NOR2_X1 U691 ( .A1(n345), .A2(n616), .ZN(n617) );
  NOR2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n623) );
  NOR2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U694 ( .A(KEYINPUT119), .B(n621), .Z(n622) );
  NOR2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n628), .B(KEYINPUT52), .ZN(n629) );
  XNOR2_X1 U699 ( .A(KEYINPUT120), .B(n629), .ZN(n630) );
  NOR2_X1 U700 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U701 ( .A(n632), .B(KEYINPUT121), .Z(n633) );
  INV_X1 U702 ( .A(KEYINPUT123), .ZN(n634) );
  XNOR2_X1 U703 ( .A(n634), .B(KEYINPUT53), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n637), .B(G143), .ZN(G45) );
  XOR2_X1 U705 ( .A(n638), .B(G140), .Z(G42) );
  XNOR2_X1 U706 ( .A(n639), .B(G119), .ZN(G21) );
  XOR2_X1 U707 ( .A(KEYINPUT110), .B(KEYINPUT62), .Z(n640) );
  XNOR2_X1 U708 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U709 ( .A(n643), .B(n642), .ZN(n645) );
  NAND2_X1 U710 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U711 ( .A(n646), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U712 ( .A(G101), .B(n647), .ZN(G3) );
  NOR2_X1 U713 ( .A1(n667), .A2(n651), .ZN(n648) );
  XOR2_X1 U714 ( .A(G104), .B(n648), .Z(G6) );
  XOR2_X1 U715 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n650) );
  XNOR2_X1 U716 ( .A(KEYINPUT111), .B(KEYINPUT27), .ZN(n649) );
  XNOR2_X1 U717 ( .A(n650), .B(n649), .ZN(n655) );
  NOR2_X1 U718 ( .A1(n671), .A2(n651), .ZN(n653) );
  XNOR2_X1 U719 ( .A(G107), .B(KEYINPUT26), .ZN(n652) );
  XNOR2_X1 U720 ( .A(n653), .B(n652), .ZN(n654) );
  XOR2_X1 U721 ( .A(n655), .B(n654), .Z(G9) );
  XNOR2_X1 U722 ( .A(G110), .B(n656), .ZN(G12) );
  INV_X1 U723 ( .A(n671), .ZN(n657) );
  NAND2_X1 U724 ( .A1(n658), .A2(n657), .ZN(n661) );
  INV_X1 U725 ( .A(n659), .ZN(n660) );
  NOR2_X1 U726 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U727 ( .A(G128), .B(KEYINPUT29), .ZN(n662) );
  XNOR2_X1 U728 ( .A(n663), .B(n662), .ZN(G30) );
  NOR2_X1 U729 ( .A1(n664), .A2(n667), .ZN(n665) );
  XOR2_X1 U730 ( .A(KEYINPUT114), .B(n665), .Z(n666) );
  XNOR2_X1 U731 ( .A(G146), .B(n666), .ZN(G48) );
  NOR2_X1 U732 ( .A1(n667), .A2(n670), .ZN(n669) );
  XNOR2_X1 U733 ( .A(G113), .B(KEYINPUT115), .ZN(n668) );
  XNOR2_X1 U734 ( .A(n669), .B(n668), .ZN(G15) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U736 ( .A(G116), .B(n672), .Z(G18) );
  XNOR2_X1 U737 ( .A(G125), .B(n673), .ZN(n674) );
  XNOR2_X1 U738 ( .A(n674), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U739 ( .A(G134), .B(n675), .Z(G36) );
  NAND2_X1 U740 ( .A1(n690), .A2(G469), .ZN(n680) );
  XOR2_X1 U741 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n678) );
  XNOR2_X1 U742 ( .A(n676), .B(KEYINPUT124), .ZN(n677) );
  XNOR2_X1 U743 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U744 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U745 ( .A1(n696), .A2(n681), .ZN(G54) );
  XOR2_X1 U746 ( .A(n682), .B(KEYINPUT59), .Z(n683) );
  XNOR2_X1 U747 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U748 ( .A(n686), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U749 ( .A1(n690), .A2(G478), .ZN(n688) );
  XNOR2_X1 U750 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X1 U751 ( .A1(n696), .A2(n689), .ZN(G63) );
  NAND2_X1 U752 ( .A1(n690), .A2(G217), .ZN(n694) );
  NOR2_X1 U753 ( .A1(n696), .A2(n695), .ZN(G66) );
  INV_X1 U754 ( .A(n697), .ZN(n698) );
  NOR2_X1 U755 ( .A1(n698), .A2(G953), .ZN(n703) );
  NAND2_X1 U756 ( .A1(G953), .A2(G224), .ZN(n699) );
  XOR2_X1 U757 ( .A(KEYINPUT61), .B(n699), .Z(n700) );
  NOR2_X1 U758 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U759 ( .A1(n703), .A2(n702), .ZN(n709) );
  XNOR2_X1 U760 ( .A(G101), .B(KEYINPUT126), .ZN(n704) );
  XNOR2_X1 U761 ( .A(n705), .B(n704), .ZN(n707) );
  NAND2_X1 U762 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n709), .B(n708), .ZN(G69) );
  OR2_X1 U764 ( .A1(n711), .A2(n710), .ZN(n717) );
  XOR2_X1 U765 ( .A(KEYINPUT127), .B(n712), .Z(n713) );
  XNOR2_X1 U766 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U767 ( .A(n716), .B(n715), .ZN(n720) );
  XNOR2_X1 U768 ( .A(n717), .B(n720), .ZN(n719) );
  NAND2_X1 U769 ( .A1(n719), .A2(n718), .ZN(n724) );
  XNOR2_X1 U770 ( .A(G227), .B(n720), .ZN(n721) );
  NAND2_X1 U771 ( .A1(n721), .A2(G900), .ZN(n722) );
  NAND2_X1 U772 ( .A1(n722), .A2(G953), .ZN(n723) );
  NAND2_X1 U773 ( .A1(n724), .A2(n723), .ZN(G72) );
  XOR2_X1 U774 ( .A(n725), .B(G131), .Z(G33) );
  XNOR2_X1 U775 ( .A(n726), .B(G122), .ZN(G24) );
  XOR2_X1 U776 ( .A(G137), .B(n727), .Z(G39) );
endmodule

