//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968;
  OAI21_X1  g000(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT92), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT93), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NOR3_X1   g005(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n204), .B(KEYINPUT93), .ZN(new_n209));
  INV_X1    g008(.A(new_n207), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n214), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  OR3_X1    g014(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT15), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n208), .A2(new_n211), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n210), .A2(KEYINPUT90), .A3(new_n202), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  OAI22_X1  g019(.A1(new_n202), .A2(KEYINPUT90), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(KEYINPUT15), .B(new_n212), .C1(new_n218), .C2(new_n221), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n217), .A2(KEYINPUT94), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT94), .B1(new_n217), .B2(new_n222), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT7), .ZN(new_n227));
  INV_X1    g026(.A(G99gat), .ZN(new_n228));
  INV_X1    g027(.A(G106gat), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT8), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n227), .B(new_n230), .C1(G85gat), .C2(G92gat), .ZN(new_n231));
  XOR2_X1   g030(.A(G99gat), .B(G106gat), .Z(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n225), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n223), .B2(new_n224), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT95), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n217), .A2(KEYINPUT17), .A3(new_n222), .ZN(new_n239));
  OAI211_X1 g038(.A(KEYINPUT95), .B(new_n235), .C1(new_n223), .C2(new_n224), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT101), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n234), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n238), .A2(new_n242), .A3(new_n239), .A4(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n233), .ZN(new_n245));
  INV_X1    g044(.A(G232gat), .ZN(new_n246));
  INV_X1    g045(.A(G233gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n243), .A2(new_n245), .B1(KEYINPUT41), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n248), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT41), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n243), .A2(new_n245), .A3(new_n251), .A4(new_n250), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G134gat), .B(G162gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(G190gat), .B(G218gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n253), .A2(new_n254), .A3(new_n258), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G127gat), .B(G155gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(G231gat), .A2(G233gat), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G15gat), .B(G22gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT96), .ZN(new_n268));
  INV_X1    g067(.A(G1gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n267), .ZN(new_n270));
  OAI22_X1  g069(.A1(new_n268), .A2(new_n269), .B1(new_n270), .B2(KEYINPUT16), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(new_n269), .B2(new_n268), .ZN(new_n272));
  INV_X1    g071(.A(G8gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G57gat), .B(G64gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT9), .ZN(new_n276));
  NAND2_X1  g075(.A1(G71gat), .A2(G78gat), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(G71gat), .B(G78gat), .Z(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n278), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT21), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OR3_X1    g082(.A1(new_n274), .A2(KEYINPUT100), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT100), .B1(new_n274), .B2(new_n283), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT99), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT99), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n284), .A2(new_n288), .A3(new_n285), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n281), .A2(new_n282), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n291), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n287), .A2(new_n293), .A3(new_n289), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n266), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n297));
  XNOR2_X1  g096(.A(G183gat), .B(G211gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n292), .A2(new_n294), .A3(new_n266), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n299), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n292), .A2(new_n294), .A3(new_n266), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(new_n295), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n262), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT4), .ZN(new_n307));
  INV_X1    g106(.A(G134gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G127gat), .ZN(new_n309));
  INV_X1    g108(.A(G127gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G134gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT68), .ZN(new_n312));
  OR3_X1    g111(.A1(new_n310), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(G113gat), .B(G120gat), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n312), .B(new_n313), .C1(KEYINPUT1), .C2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G120gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G113gat), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G120gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT1), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n323), .A2(KEYINPUT69), .A3(new_n313), .A4(new_n312), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n309), .A2(new_n311), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n322), .A2(new_n326), .A3(KEYINPUT70), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT70), .B1(new_n322), .B2(new_n326), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G141gat), .B(G148gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  OR2_X1    g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(KEYINPUT2), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n332), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n334), .B(new_n333), .C1(new_n331), .C2(KEYINPUT2), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n307), .B1(new_n330), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(KEYINPUT3), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n330), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n339), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n325), .A2(new_n346), .A3(new_n329), .A4(KEYINPUT4), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n340), .A2(new_n344), .A3(new_n345), .A4(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n345), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n325), .A2(new_n346), .A3(new_n329), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n346), .B1(new_n325), .B2(new_n329), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n354), .A2(KEYINPUT5), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(KEYINPUT5), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n349), .A3(new_n348), .ZN(new_n358));
  XOR2_X1   g157(.A(G1gat), .B(G29gat), .Z(new_n359));
  XNOR2_X1  g158(.A(G57gat), .B(G85gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(new_n358), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n364), .B1(new_n356), .B2(new_n358), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(KEYINPUT6), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n367), .B1(new_n369), .B2(new_n365), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT86), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n374));
  AND2_X1   g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(G197gat), .A2(G204gat), .ZN(new_n376));
  OAI22_X1  g175(.A1(new_n374), .A2(KEYINPUT77), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n374), .A2(KEYINPUT77), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(G211gat), .B(G218gat), .Z(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n374), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n374), .A2(KEYINPUT77), .ZN(new_n385));
  INV_X1    g184(.A(new_n376), .ZN(new_n386));
  NAND2_X1  g185(.A1(G197gat), .A2(G204gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n380), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n373), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n381), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G226gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n247), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(KEYINPUT29), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT26), .ZN(new_n398));
  NOR2_X1   g197(.A1(G169gat), .A2(G176gat), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n400), .A2(new_n401), .B1(G183gat), .B2(G190gat), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT28), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT27), .ZN(new_n404));
  INV_X1    g203(.A(G183gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n407));
  AOI21_X1  g206(.A(G190gat), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT67), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n403), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G190gat), .ZN(new_n411));
  AND2_X1   g210(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n402), .A2(new_n410), .A3(new_n415), .ZN(new_n416));
  AND3_X1   g215(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT25), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n397), .ZN(new_n423));
  INV_X1    g222(.A(G169gat), .ZN(new_n424));
  INV_X1    g223(.A(G176gat), .ZN(new_n425));
  AND4_X1   g224(.A1(KEYINPUT64), .A2(new_n424), .A3(new_n425), .A4(KEYINPUT23), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT64), .B1(new_n399), .B2(KEYINPUT23), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n399), .A2(KEYINPUT23), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n422), .A2(new_n423), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n416), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT25), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n397), .A2(KEYINPUT65), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT24), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(new_n405), .B2(new_n411), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT66), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n420), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT66), .B1(new_n417), .B2(new_n418), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n399), .A2(KEYINPUT23), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n397), .A2(KEYINPUT65), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n429), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n432), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT79), .B1(new_n431), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n436), .B1(new_n435), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n421), .B1(new_n418), .B2(KEYINPUT66), .ZN(new_n448));
  OAI22_X1  g247(.A1(new_n447), .A2(new_n448), .B1(KEYINPUT65), .B2(new_n397), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT25), .B1(new_n449), .B2(new_n442), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT79), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n430), .A4(new_n416), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n396), .B1(new_n445), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n430), .A3(new_n416), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n454), .A2(new_n393), .A3(new_n247), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n392), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT30), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n445), .A2(new_n394), .A3(new_n452), .ZN(new_n458));
  INV_X1    g257(.A(new_n392), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n454), .A2(new_n395), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n456), .A2(new_n457), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G64gat), .B(G92gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(G36gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT80), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(new_n273), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n457), .B1(new_n456), .B2(new_n461), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI211_X1 g268(.A(new_n457), .B(new_n466), .C1(new_n456), .C2(new_n461), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n372), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n461), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT30), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n466), .A3(new_n462), .ZN(new_n474));
  INV_X1    g273(.A(new_n470), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT86), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT31), .B(G50gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(G78gat), .B(G106gat), .Z(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G228gat), .A2(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT29), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n381), .A2(new_n391), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n346), .B1(new_n484), .B2(new_n341), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n381), .A2(new_n391), .B1(new_n342), .B2(new_n483), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G22gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n483), .B1(new_n389), .B2(new_n390), .ZN(new_n489));
  INV_X1    g288(.A(new_n377), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n380), .B1(new_n490), .B2(new_n385), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n341), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n339), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n342), .A2(new_n483), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n392), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n481), .A3(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n487), .A2(new_n488), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n488), .B1(new_n487), .B2(new_n496), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n480), .B1(new_n499), .B2(KEYINPUT84), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n487), .A2(new_n496), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(G22gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n488), .A3(new_n496), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n502), .A2(KEYINPUT84), .A3(new_n503), .A4(new_n480), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n478), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(KEYINPUT84), .A3(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n479), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(new_n477), .A3(new_n504), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n471), .A2(new_n476), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT71), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n431), .B2(new_n444), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n450), .A2(KEYINPUT71), .A3(new_n430), .A4(new_n416), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n330), .A3(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n454), .A2(new_n511), .A3(new_n325), .A4(new_n329), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G227gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(new_n247), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n516), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n516), .B2(new_n519), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n514), .A2(new_n518), .A3(new_n515), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G43gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(G71gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(new_n228), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT33), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(KEYINPUT32), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT73), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n524), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n527), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n524), .B2(KEYINPUT32), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT33), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n524), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n535), .A2(KEYINPUT72), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT72), .B1(new_n535), .B2(new_n537), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n523), .B(new_n533), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT76), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n524), .A2(KEYINPUT32), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n542), .A3(new_n527), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT72), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n535), .A2(KEYINPUT72), .A3(new_n537), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n523), .B1(new_n547), .B2(new_n533), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT76), .ZN(new_n551));
  INV_X1    g350(.A(new_n523), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n371), .B(new_n510), .C1(new_n549), .C2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT35), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n506), .A2(new_n509), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n550), .A2(new_n552), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT75), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n560), .A3(new_n540), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n550), .A2(KEYINPUT75), .A3(new_n552), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n469), .A2(new_n470), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n356), .A2(new_n358), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n363), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT83), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n567), .A3(new_n366), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT83), .B1(new_n368), .B2(KEYINPUT6), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(new_n365), .ZN(new_n570));
  INV_X1    g369(.A(new_n367), .ZN(new_n571));
  AOI211_X1 g370(.A(new_n556), .B(new_n564), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n555), .A2(new_n556), .B1(new_n563), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n365), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n574), .B1(new_n369), .B2(new_n567), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n367), .B1(new_n575), .B2(new_n569), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n506), .A2(KEYINPUT85), .A3(new_n509), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT85), .B1(new_n506), .B2(new_n509), .ZN(new_n578));
  OAI22_X1  g377(.A1(new_n576), .A2(new_n564), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT37), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n472), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n472), .A2(new_n580), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT38), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n466), .B1(new_n472), .B2(KEYINPUT38), .ZN(new_n585));
  OR3_X1    g384(.A1(new_n453), .A2(new_n455), .A3(new_n392), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n458), .A2(new_n460), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n586), .B(KEYINPUT37), .C1(new_n587), .C2(new_n459), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT38), .ZN(new_n589));
  INV_X1    g388(.A(new_n466), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n588), .A2(new_n581), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n370), .A2(new_n584), .A3(new_n585), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n340), .A2(new_n344), .A3(new_n347), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n351), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT87), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n595), .A2(new_n596), .A3(new_n363), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n595), .B2(new_n363), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n352), .A2(new_n353), .A3(new_n351), .ZN(new_n599));
  AOI211_X1 g398(.A(new_n594), .B(new_n599), .C1(new_n351), .C2(new_n593), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT88), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT40), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n603), .A2(new_n471), .A3(new_n365), .A4(new_n476), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT40), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n592), .B(new_n557), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n559), .A2(KEYINPUT76), .A3(new_n540), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n607), .A2(new_n608), .A3(new_n553), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(new_n561), .B2(new_n562), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n579), .B(new_n606), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n573), .A2(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n233), .A2(new_n281), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n233), .A2(new_n281), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n613), .A2(new_n616), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(G230gat), .A3(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(new_n425), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G204gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n620), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n619), .B(KEYINPUT102), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(new_n615), .B2(new_n617), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n625), .B1(new_n631), .B2(new_n622), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G113gat), .B(G141gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G169gat), .B(G197gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n274), .B1(new_n223), .B2(new_n224), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT97), .ZN(new_n642));
  INV_X1    g441(.A(new_n274), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n238), .A2(new_n643), .A3(new_n239), .A4(new_n240), .ZN(new_n644));
  NAND2_X1  g443(.A1(G229gat), .A2(G233gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT18), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n640), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n642), .B1(new_n274), .B2(new_n225), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n645), .B(KEYINPUT13), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n642), .A2(new_n644), .A3(KEYINPUT18), .A4(new_n645), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n648), .A3(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n650), .A2(new_n655), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND4_X1   g457(.A1(new_n306), .A2(new_n612), .A3(new_n633), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n576), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g460(.A1(new_n471), .A2(new_n476), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n659), .B(new_n663), .C1(KEYINPUT16), .C2(G8gat), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT103), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n273), .B1(new_n659), .B2(new_n663), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n665), .B2(KEYINPUT42), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(KEYINPUT103), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(G1325gat));
  NAND2_X1  g470(.A1(new_n607), .A2(new_n553), .ZN(new_n672));
  AOI21_X1  g471(.A(G15gat), .B1(new_n659), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n609), .A2(new_n610), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n659), .A2(G15gat), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n577), .A2(new_n578), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n659), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(new_n262), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n573), .B2(new_n611), .ZN(new_n683));
  INV_X1    g482(.A(new_n305), .ZN(new_n684));
  INV_X1    g483(.A(new_n633), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n650), .A2(new_n655), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n650), .A2(new_n655), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n219), .A3(new_n576), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT45), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n260), .A2(KEYINPUT104), .A3(new_n261), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT104), .B1(new_n260), .B2(new_n261), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n612), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n683), .B2(new_n697), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n699), .A2(new_n689), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n576), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT105), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n692), .B1(new_n702), .B2(new_n219), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g504(.A(KEYINPUT106), .B(new_n692), .C1(new_n702), .C2(new_n219), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1328gat));
  NAND3_X1  g506(.A1(new_n690), .A2(new_n220), .A3(new_n663), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT46), .Z(new_n709));
  NAND2_X1  g508(.A1(new_n700), .A2(new_n663), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n220), .B2(new_n711), .ZN(G1329gat));
  NAND2_X1  g511(.A1(new_n700), .A2(new_n674), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G43gat), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715));
  INV_X1    g514(.A(G43gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n690), .A2(new_n716), .A3(new_n672), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n715), .B1(new_n714), .B2(new_n717), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT47), .B1(new_n717), .B2(KEYINPUT107), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1330gat));
  INV_X1    g521(.A(G50gat), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n700), .B2(new_n678), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n690), .A2(new_n723), .A3(new_n678), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(KEYINPUT109), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n728), .B(new_n723), .C1(new_n700), .C2(new_n558), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n725), .B1(new_n730), .B2(KEYINPUT48), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n727), .A2(KEYINPUT48), .B1(new_n729), .B2(new_n731), .ZN(G1331gat));
  NOR3_X1   g531(.A1(new_n262), .A2(new_n658), .A3(new_n305), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n612), .A2(new_n685), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n576), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n663), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  AOI21_X1  g539(.A(G71gat), .B1(new_n734), .B2(new_n672), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n734), .A2(G71gat), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n674), .B2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n678), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n684), .A2(new_n658), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n683), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n683), .A2(KEYINPUT51), .A3(new_n747), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n633), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n576), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n684), .A2(new_n658), .A3(new_n633), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n699), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G85gat), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n753), .B1(new_n758), .B2(new_n576), .ZN(G1336gat));
  NAND2_X1  g558(.A1(new_n750), .A2(new_n751), .ZN(new_n760));
  INV_X1    g559(.A(G92gat), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n760), .A2(new_n761), .A3(new_n685), .A4(new_n663), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n697), .B1(new_n612), .B2(new_n262), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n764));
  INV_X1    g563(.A(new_n261), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n258), .B1(new_n253), .B2(new_n254), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n767), .A2(new_n693), .A3(new_n697), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n573), .B2(new_n611), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n663), .B(new_n754), .C1(new_n763), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G92gat), .ZN(new_n771));
  XOR2_X1   g570(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n772));
  NAND3_X1  g571(.A1(new_n762), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(KEYINPUT110), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n770), .A2(new_n775), .A3(G92gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n762), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT52), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n777), .B2(KEYINPUT52), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n773), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(KEYINPUT113), .B(new_n773), .C1(new_n779), .C2(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1337gat));
  NAND3_X1  g584(.A1(new_n752), .A2(new_n228), .A3(new_n672), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n756), .A2(new_n674), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n788), .B2(new_n228), .ZN(G1338gat));
  NAND3_X1  g588(.A1(new_n752), .A2(new_n229), .A3(new_n558), .ZN(new_n790));
  XOR2_X1   g589(.A(KEYINPUT114), .B(G106gat), .Z(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n755), .B2(new_n557), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n791), .B1(new_n755), .B2(new_n677), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n790), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT53), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n794), .A2(new_n795), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n796), .A2(new_n799), .A3(new_n800), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n651), .A2(new_n652), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n645), .B1(new_n642), .B2(new_n644), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n638), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n653), .A2(new_n648), .A3(new_n640), .A4(new_n654), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n805), .A3(new_n685), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n620), .B(KEYINPUT54), .C1(new_n618), .C2(new_n628), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n625), .B1(new_n630), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n807), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n810), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(KEYINPUT55), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n626), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n806), .B1(new_n688), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(new_n694), .B2(new_n695), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n804), .A2(new_n805), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n767), .A2(new_n693), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n684), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n733), .A2(new_n633), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n563), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n576), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n663), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n320), .A3(new_n658), .ZN(new_n829));
  INV_X1    g628(.A(new_n826), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n677), .A2(new_n672), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n822), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G113gat), .B1(new_n833), .B2(new_n688), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n829), .A2(new_n834), .ZN(G1340gat));
  NAND3_X1  g634(.A1(new_n828), .A2(new_n318), .A3(new_n685), .ZN(new_n836));
  OAI21_X1  g635(.A(G120gat), .B1(new_n833), .B2(new_n633), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1341gat));
  AOI21_X1  g637(.A(G127gat), .B1(new_n828), .B2(new_n684), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n305), .A2(new_n310), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n832), .B2(new_n840), .ZN(G1342gat));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n576), .A3(new_n262), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(G134gat), .A3(new_n663), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT56), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n833), .B2(new_n682), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1343gat));
  INV_X1    g645(.A(G141gat), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n848), .B(new_n558), .C1(new_n820), .C2(new_n821), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n674), .A2(new_n830), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT117), .B1(new_n808), .B2(new_n810), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT55), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n626), .B(new_n852), .C1(new_n686), .C2(new_n687), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n262), .B1(new_n853), .B2(new_n806), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n819), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT118), .B(new_n262), .C1(new_n806), .C2(new_n853), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n305), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n733), .A2(new_n633), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n677), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n849), .B(new_n850), .C1(new_n860), .C2(new_n848), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT119), .ZN(new_n862));
  INV_X1    g661(.A(new_n806), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n851), .B(new_n807), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(new_n656), .B2(new_n657), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n865), .B2(new_n626), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT118), .B1(new_n866), .B2(new_n262), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n854), .A2(new_n855), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n819), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n821), .B1(new_n869), .B2(new_n305), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT57), .B1(new_n870), .B2(new_n677), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n871), .A2(new_n872), .A3(new_n849), .A4(new_n850), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n862), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n847), .B1(new_n874), .B2(new_n658), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n822), .A2(new_n557), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n876), .A2(new_n847), .A3(new_n658), .A4(new_n850), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT58), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n877), .B(KEYINPUT120), .Z(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  OAI21_X1  g680(.A(G141gat), .B1(new_n861), .B2(new_n688), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n879), .A2(new_n883), .ZN(G1344gat));
  AOI21_X1  g683(.A(new_n633), .B1(new_n862), .B2(new_n873), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n262), .A2(new_n818), .ZN(new_n886));
  OAI211_X1 g685(.A(KEYINPUT122), .B(new_n886), .C1(new_n866), .C2(new_n262), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n262), .A2(new_n818), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n854), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n305), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n859), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n821), .A2(KEYINPUT121), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n848), .A3(new_n678), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT57), .B1(new_n822), .B2(new_n557), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n850), .A2(KEYINPUT59), .A3(new_n685), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n885), .A2(KEYINPUT59), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n876), .A2(new_n850), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(G148gat), .B1(new_n902), .B2(new_n685), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n900), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n903), .ZN(G1345gat));
  AOI21_X1  g703(.A(G155gat), .B1(new_n902), .B2(new_n684), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n305), .B1(new_n862), .B2(new_n873), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(G155gat), .ZN(G1346gat));
  INV_X1    g706(.A(G162gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n902), .A2(new_n908), .A3(new_n262), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n874), .A2(new_n696), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n908), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n576), .A2(new_n662), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n824), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n424), .A3(new_n658), .ZN(new_n915));
  INV_X1    g714(.A(new_n912), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n822), .A2(new_n831), .A3(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n658), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n915), .B1(new_n922), .B2(new_n424), .ZN(G1348gat));
  NAND3_X1  g722(.A1(new_n921), .A2(G176gat), .A3(new_n685), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n425), .B1(new_n913), .B2(new_n633), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n920), .A3(new_n684), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G183gat), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n914), .B(new_n684), .C1(new_n413), .C2(new_n412), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n932), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n914), .A2(new_n411), .A3(new_n696), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT124), .Z(new_n936));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n920), .A3(new_n262), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G190gat), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n936), .A2(new_n940), .A3(new_n941), .ZN(G1351gat));
  NOR2_X1   g741(.A1(new_n674), .A2(new_n916), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n898), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n946), .B1(new_n945), .B2(new_n898), .ZN(new_n947));
  OAI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n688), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n876), .A2(new_n943), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n949), .A2(G197gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n948), .B1(new_n688), .B2(new_n950), .ZN(G1352gat));
  XOR2_X1   g750(.A(KEYINPUT126), .B(G204gat), .Z(new_n952));
  OAI21_X1  g751(.A(new_n952), .B1(new_n947), .B2(new_n633), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n949), .A2(new_n633), .A3(new_n952), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1353gat));
  OR3_X1    g755(.A1(new_n949), .A2(G211gat), .A3(new_n305), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n896), .A2(new_n897), .A3(new_n684), .A4(new_n943), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT127), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n963), .B(new_n957), .C1(new_n959), .C2(new_n960), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1354gat));
  OAI21_X1  g764(.A(G218gat), .B1(new_n947), .B2(new_n682), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n949), .A2(G218gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(new_n696), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1355gat));
endmodule


