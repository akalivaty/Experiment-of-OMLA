

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744;

  XNOR2_X1 U377 ( .A(n400), .B(n440), .ZN(n465) );
  NAND2_X1 U378 ( .A1(n384), .A2(n381), .ZN(n531) );
  XNOR2_X1 U379 ( .A(KEYINPUT41), .B(n503), .ZN(n541) );
  XNOR2_X2 U380 ( .A(n536), .B(KEYINPUT40), .ZN(n744) );
  XNOR2_X2 U381 ( .A(G104), .B(KEYINPUT77), .ZN(n380) );
  XNOR2_X2 U382 ( .A(n470), .B(n469), .ZN(n553) );
  OR2_X2 U383 ( .A1(n655), .A2(n640), .ZN(n470) );
  XNOR2_X2 U384 ( .A(n456), .B(n455), .ZN(n715) );
  XNOR2_X2 U385 ( .A(n364), .B(n435), .ZN(n456) );
  NOR2_X2 U386 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X2 U387 ( .A(n531), .B(n408), .ZN(n451) );
  AND2_X2 U388 ( .A1(n667), .A2(n664), .ZN(n362) );
  XNOR2_X2 U389 ( .A(n605), .B(KEYINPUT32), .ZN(n667) );
  INV_X2 U390 ( .A(G953), .ZN(n733) );
  XNOR2_X1 U391 ( .A(G119), .B(G116), .ZN(n366) );
  XNOR2_X1 U392 ( .A(G113), .B(KEYINPUT73), .ZN(n365) );
  AND2_X1 U393 ( .A1(n573), .A2(n572), .ZN(n575) );
  NOR2_X1 U394 ( .A1(n552), .A2(n391), .ZN(n573) );
  AND2_X1 U395 ( .A1(n620), .A2(n388), .ZN(n360) );
  AND2_X1 U396 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U397 ( .A1(n710), .A2(n359), .ZN(n617) );
  XNOR2_X1 U398 ( .A(n611), .B(KEYINPUT31), .ZN(n710) );
  NOR2_X1 U399 ( .A1(n615), .A2(n599), .ZN(n600) );
  XNOR2_X1 U400 ( .A(n590), .B(n393), .ZN(n615) );
  NOR2_X1 U401 ( .A1(n588), .A2(n587), .ZN(n590) );
  AND2_X1 U402 ( .A1(n386), .A2(n385), .ZN(n384) );
  XNOR2_X1 U403 ( .A(n465), .B(n405), .ZN(n683) );
  XNOR2_X1 U404 ( .A(n366), .B(n365), .ZN(n364) );
  XNOR2_X1 U405 ( .A(G143), .B(G128), .ZN(n480) );
  INV_X1 U406 ( .A(KEYINPUT67), .ZN(n397) );
  INV_X1 U407 ( .A(n409), .ZN(n355) );
  NAND2_X2 U408 ( .A1(n608), .A2(n362), .ZN(n621) );
  XNOR2_X2 U409 ( .A(n377), .B(n376), .ZN(n608) );
  AND2_X2 U410 ( .A1(n645), .A2(n644), .ZN(n356) );
  AND2_X2 U411 ( .A1(n645), .A2(n644), .ZN(n682) );
  NAND2_X1 U412 ( .A1(n384), .A2(n381), .ZN(n357) );
  NAND2_X1 U413 ( .A1(n369), .A2(n368), .ZN(n367) );
  AND2_X2 U414 ( .A1(n450), .A2(n451), .ZN(n510) );
  INV_X1 U415 ( .A(KEYINPUT86), .ZN(n388) );
  NAND2_X1 U416 ( .A1(n371), .A2(n370), .ZN(n369) );
  NAND2_X1 U417 ( .A1(n387), .A2(KEYINPUT86), .ZN(n373) );
  NAND2_X1 U418 ( .A1(n360), .A2(n375), .ZN(n374) );
  NOR2_X1 U419 ( .A1(n537), .A2(n529), .ZN(n545) );
  NAND2_X1 U420 ( .A1(n383), .A2(n486), .ZN(n382) );
  XNOR2_X1 U421 ( .A(n380), .B(G107), .ZN(n379) );
  XNOR2_X1 U422 ( .A(n594), .B(n593), .ZN(n378) );
  XNOR2_X1 U423 ( .A(n544), .B(n543), .ZN(n552) );
  NAND2_X1 U424 ( .A1(n407), .A2(G902), .ZN(n385) );
  XNOR2_X1 U425 ( .A(G134), .B(G107), .ZN(n475) );
  XNOR2_X1 U426 ( .A(n713), .B(KEYINPUT74), .ZN(n400) );
  NOR2_X1 U427 ( .A1(KEYINPUT2), .A2(n638), .ZN(n625) );
  AND2_X1 U428 ( .A1(n389), .A2(n613), .ZN(n535) );
  INV_X1 U429 ( .A(KEYINPUT1), .ZN(n408) );
  XNOR2_X1 U430 ( .A(n555), .B(n554), .ZN(n588) );
  NAND2_X1 U431 ( .A1(n642), .A2(n641), .ZN(n645) );
  XNOR2_X1 U432 ( .A(n648), .B(n647), .ZN(n649) );
  INV_X1 U433 ( .A(KEYINPUT35), .ZN(n376) );
  NAND2_X1 U434 ( .A1(n361), .A2(n358), .ZN(n619) );
  XNOR2_X1 U435 ( .A(n619), .B(G101), .ZN(G3) );
  AND2_X1 U436 ( .A1(n560), .A2(n609), .ZN(n358) );
  NOR2_X1 U437 ( .A1(n615), .A2(n614), .ZN(n359) );
  AND2_X1 U438 ( .A1(n606), .A2(n409), .ZN(n361) );
  XNOR2_X1 U439 ( .A(n379), .B(n396), .ZN(n713) );
  AND2_X1 U440 ( .A1(KEYINPUT44), .A2(KEYINPUT86), .ZN(n363) );
  NOR2_X1 U441 ( .A1(n372), .A2(n367), .ZN(n623) );
  NAND2_X1 U442 ( .A1(n621), .A2(n363), .ZN(n368) );
  INV_X1 U443 ( .A(KEYINPUT44), .ZN(n370) );
  INV_X1 U444 ( .A(n621), .ZN(n371) );
  NAND2_X1 U445 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U446 ( .A1(n621), .A2(KEYINPUT44), .ZN(n375) );
  INV_X1 U447 ( .A(n608), .ZN(n668) );
  NAND2_X1 U448 ( .A1(n378), .A2(n596), .ZN(n377) );
  OR2_X1 U449 ( .A1(n683), .A2(n382), .ZN(n381) );
  INV_X1 U450 ( .A(n407), .ZN(n383) );
  NAND2_X1 U451 ( .A1(n683), .A2(n407), .ZN(n386) );
  INV_X1 U452 ( .A(n620), .ZN(n387) );
  AND2_X1 U453 ( .A1(n545), .A2(n530), .ZN(n389) );
  OR2_X1 U454 ( .A1(G902), .A2(n648), .ZN(n390) );
  XNOR2_X1 U455 ( .A(KEYINPUT82), .B(n701), .ZN(n391) );
  XOR2_X1 U456 ( .A(KEYINPUT87), .B(KEYINPUT36), .Z(n392) );
  XOR2_X1 U457 ( .A(n589), .B(KEYINPUT0), .Z(n393) );
  AND2_X1 U458 ( .A1(G221), .A2(n483), .ZN(n394) );
  XNOR2_X1 U459 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n543) );
  XNOR2_X1 U460 ( .A(G137), .B(KEYINPUT5), .ZN(n441) );
  XNOR2_X1 U461 ( .A(KEYINPUT106), .B(KEYINPUT30), .ZN(n527) );
  XNOR2_X1 U462 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U463 ( .A(n528), .B(n527), .ZN(n529) );
  BUF_X1 U464 ( .A(n636), .Z(n718) );
  NOR2_X2 U465 ( .A1(n624), .A2(n718), .ZN(n643) );
  INV_X1 U466 ( .A(KEYINPUT60), .ZN(n653) );
  XNOR2_X1 U467 ( .A(n634), .B(n633), .ZN(G75) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n395) );
  XNOR2_X1 U469 ( .A(n395), .B(KEYINPUT14), .ZN(n523) );
  NAND2_X1 U470 ( .A1(G952), .A2(n523), .ZN(n522) );
  XOR2_X1 U471 ( .A(KEYINPUT90), .B(G110), .Z(n396) );
  XNOR2_X1 U472 ( .A(n397), .B(KEYINPUT4), .ZN(n398) );
  XNOR2_X1 U473 ( .A(n480), .B(n398), .ZN(n731) );
  XNOR2_X1 U474 ( .A(KEYINPUT66), .B(G101), .ZN(n399) );
  XNOR2_X1 U475 ( .A(n731), .B(n399), .ZN(n440) );
  XNOR2_X1 U476 ( .A(G131), .B(KEYINPUT69), .ZN(n489) );
  XNOR2_X1 U477 ( .A(n489), .B(G134), .ZN(n442) );
  INV_X1 U478 ( .A(G140), .ZN(n665) );
  XNOR2_X1 U479 ( .A(n665), .B(G137), .ZN(n410) );
  INV_X1 U480 ( .A(n410), .ZN(n401) );
  XNOR2_X1 U481 ( .A(n442), .B(n401), .ZN(n729) );
  XNOR2_X1 U482 ( .A(G146), .B(KEYINPUT80), .ZN(n403) );
  NAND2_X1 U483 ( .A1(n733), .A2(G227), .ZN(n402) );
  XNOR2_X1 U484 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U485 ( .A(n729), .B(n404), .ZN(n405) );
  XNOR2_X1 U486 ( .A(KEYINPUT72), .B(G469), .ZN(n406) );
  XNOR2_X1 U487 ( .A(n406), .B(KEYINPUT71), .ZN(n407) );
  INV_X1 U488 ( .A(n451), .ZN(n409) );
  XNOR2_X1 U489 ( .A(G119), .B(G128), .ZN(n411) );
  XNOR2_X1 U490 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U491 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n413) );
  XNOR2_X1 U492 ( .A(G110), .B(KEYINPUT79), .ZN(n412) );
  XNOR2_X1 U493 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U494 ( .A(n415), .B(n414), .Z(n419) );
  XNOR2_X1 U495 ( .A(G146), .B(G125), .ZN(n461) );
  XNOR2_X1 U496 ( .A(n461), .B(KEYINPUT10), .ZN(n728) );
  XOR2_X1 U497 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n417) );
  NAND2_X1 U498 ( .A1(G234), .A2(n733), .ZN(n416) );
  XNOR2_X1 U499 ( .A(n417), .B(n416), .ZN(n483) );
  XNOR2_X1 U500 ( .A(n728), .B(n394), .ZN(n418) );
  XNOR2_X1 U501 ( .A(n419), .B(n418), .ZN(n674) );
  INV_X1 U502 ( .A(G902), .ZN(n486) );
  NAND2_X1 U503 ( .A1(n674), .A2(n486), .ZN(n427) );
  XNOR2_X1 U504 ( .A(KEYINPUT78), .B(KEYINPUT25), .ZN(n423) );
  XOR2_X1 U505 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n421) );
  XNOR2_X1 U506 ( .A(KEYINPUT15), .B(G902), .ZN(n635) );
  NAND2_X1 U507 ( .A1(G234), .A2(n635), .ZN(n420) );
  XNOR2_X1 U508 ( .A(n421), .B(n420), .ZN(n428) );
  NAND2_X1 U509 ( .A1(G217), .A2(n428), .ZN(n422) );
  XNOR2_X1 U510 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U511 ( .A(KEYINPUT96), .B(KEYINPUT98), .Z(n424) );
  XNOR2_X1 U512 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U513 ( .A(n427), .B(n426), .ZN(n609) );
  AND2_X1 U514 ( .A1(n428), .A2(G221), .ZN(n429) );
  XNOR2_X1 U515 ( .A(n429), .B(KEYINPUT21), .ZN(n597) );
  NAND2_X1 U516 ( .A1(n609), .A2(n597), .ZN(n532) );
  NAND2_X1 U517 ( .A1(n409), .A2(n532), .ZN(n430) );
  XOR2_X1 U518 ( .A(KEYINPUT50), .B(n430), .Z(n449) );
  INV_X1 U519 ( .A(n609), .ZN(n602) );
  INV_X1 U520 ( .A(n597), .ZN(n431) );
  NAND2_X1 U521 ( .A1(n602), .A2(n431), .ZN(n434) );
  XNOR2_X1 U522 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n432) );
  XNOR2_X1 U523 ( .A(n432), .B(KEYINPUT49), .ZN(n433) );
  XNOR2_X1 U524 ( .A(n434), .B(n433), .ZN(n447) );
  XNOR2_X1 U525 ( .A(KEYINPUT91), .B(KEYINPUT3), .ZN(n435) );
  XOR2_X1 U526 ( .A(KEYINPUT100), .B(KEYINPUT76), .Z(n437) );
  NOR2_X1 U527 ( .A1(G953), .A2(G237), .ZN(n495) );
  NAND2_X1 U528 ( .A1(n495), .A2(G210), .ZN(n436) );
  XNOR2_X1 U529 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U530 ( .A(n456), .B(n438), .ZN(n439) );
  XNOR2_X1 U531 ( .A(n440), .B(n439), .ZN(n445) );
  XOR2_X1 U532 ( .A(n443), .B(G146), .Z(n444) );
  XNOR2_X1 U533 ( .A(n445), .B(n444), .ZN(n669) );
  NAND2_X1 U534 ( .A1(n669), .A2(n486), .ZN(n446) );
  XNOR2_X2 U535 ( .A(n446), .B(G472), .ZN(n526) );
  INV_X1 U536 ( .A(n526), .ZN(n612) );
  NAND2_X1 U537 ( .A1(n447), .A2(n612), .ZN(n448) );
  NOR2_X1 U538 ( .A1(n449), .A2(n448), .ZN(n453) );
  INV_X1 U539 ( .A(n532), .ZN(n450) );
  NAND2_X1 U540 ( .A1(n510), .A2(n526), .ZN(n610) );
  INV_X1 U541 ( .A(n610), .ZN(n452) );
  NOR2_X1 U542 ( .A1(n453), .A2(n452), .ZN(n454) );
  XNOR2_X1 U543 ( .A(KEYINPUT51), .B(n454), .ZN(n504) );
  XNOR2_X1 U544 ( .A(KEYINPUT16), .B(G122), .ZN(n455) );
  XOR2_X1 U545 ( .A(KEYINPUT18), .B(KEYINPUT88), .Z(n459) );
  NAND2_X1 U546 ( .A1(G224), .A2(n733), .ZN(n457) );
  XNOR2_X1 U547 ( .A(n457), .B(KEYINPUT81), .ZN(n458) );
  XNOR2_X1 U548 ( .A(n459), .B(n458), .ZN(n463) );
  XNOR2_X1 U549 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n460) );
  XNOR2_X1 U550 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U551 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U552 ( .A(n715), .B(n464), .ZN(n466) );
  XNOR2_X1 U553 ( .A(n466), .B(n465), .ZN(n655) );
  INV_X1 U554 ( .A(n635), .ZN(n640) );
  INV_X1 U555 ( .A(G237), .ZN(n467) );
  NAND2_X1 U556 ( .A1(n486), .A2(n467), .ZN(n473) );
  NAND2_X1 U557 ( .A1(n473), .A2(G210), .ZN(n468) );
  XNOR2_X1 U558 ( .A(n468), .B(KEYINPUT93), .ZN(n469) );
  BUF_X1 U559 ( .A(n553), .Z(n471) );
  XNOR2_X1 U560 ( .A(KEYINPUT75), .B(KEYINPUT38), .ZN(n472) );
  XNOR2_X1 U561 ( .A(n471), .B(n472), .ZN(n530) );
  NAND2_X1 U562 ( .A1(n473), .A2(G214), .ZN(n474) );
  XNOR2_X1 U563 ( .A(n474), .B(KEYINPUT94), .ZN(n564) );
  AND2_X1 U564 ( .A1(n530), .A2(n564), .ZN(n507) );
  XOR2_X1 U565 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n476) );
  XNOR2_X1 U566 ( .A(n476), .B(n475), .ZN(n478) );
  XNOR2_X1 U567 ( .A(KEYINPUT103), .B(KEYINPUT7), .ZN(n477) );
  XNOR2_X1 U568 ( .A(n478), .B(n477), .ZN(n482) );
  XNOR2_X1 U569 ( .A(G116), .B(G122), .ZN(n479) );
  XNOR2_X1 U570 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U571 ( .A(n482), .B(n481), .ZN(n485) );
  AND2_X1 U572 ( .A1(n483), .A2(G217), .ZN(n484) );
  XNOR2_X1 U573 ( .A(n485), .B(n484), .ZN(n679) );
  NAND2_X1 U574 ( .A1(n679), .A2(n486), .ZN(n488) );
  INV_X1 U575 ( .A(G478), .ZN(n487) );
  XNOR2_X1 U576 ( .A(n488), .B(n487), .ZN(n547) );
  XNOR2_X1 U577 ( .A(KEYINPUT13), .B(G475), .ZN(n502) );
  XOR2_X1 U578 ( .A(n728), .B(G122), .Z(n492) );
  INV_X1 U579 ( .A(n489), .ZN(n490) );
  XNOR2_X1 U580 ( .A(G113), .B(n490), .ZN(n491) );
  XNOR2_X1 U581 ( .A(n492), .B(n491), .ZN(n501) );
  XOR2_X1 U582 ( .A(KEYINPUT101), .B(G140), .Z(n494) );
  XNOR2_X1 U583 ( .A(G143), .B(G104), .ZN(n493) );
  XNOR2_X1 U584 ( .A(n494), .B(n493), .ZN(n499) );
  XOR2_X1 U585 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n497) );
  NAND2_X1 U586 ( .A1(G214), .A2(n495), .ZN(n496) );
  XNOR2_X1 U587 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U588 ( .A(n499), .B(n498), .Z(n500) );
  XNOR2_X1 U589 ( .A(n501), .B(n500), .ZN(n648) );
  XNOR2_X1 U590 ( .A(n502), .B(n390), .ZN(n546) );
  AND2_X1 U591 ( .A1(n547), .A2(n546), .ZN(n598) );
  NAND2_X1 U592 ( .A1(n507), .A2(n598), .ZN(n503) );
  NAND2_X1 U593 ( .A1(n504), .A2(n541), .ZN(n515) );
  OR2_X1 U594 ( .A1(n530), .A2(n564), .ZN(n505) );
  NAND2_X1 U595 ( .A1(n505), .A2(n598), .ZN(n509) );
  INV_X1 U596 ( .A(n546), .ZN(n506) );
  AND2_X1 U597 ( .A1(n547), .A2(n506), .ZN(n706) );
  OR2_X1 U598 ( .A1(n547), .A2(n506), .ZN(n697) );
  INV_X1 U599 ( .A(n697), .ZN(n709) );
  NOR2_X1 U600 ( .A1(n706), .A2(n709), .ZN(n558) );
  INV_X1 U601 ( .A(n558), .ZN(n616) );
  NAND2_X1 U602 ( .A1(n507), .A2(n616), .ZN(n508) );
  NAND2_X1 U603 ( .A1(n509), .A2(n508), .ZN(n513) );
  XNOR2_X1 U604 ( .A(n510), .B(KEYINPUT104), .ZN(n511) );
  XNOR2_X1 U605 ( .A(n526), .B(KEYINPUT6), .ZN(n560) );
  INV_X1 U606 ( .A(n560), .ZN(n601) );
  NAND2_X1 U607 ( .A1(n511), .A2(n601), .ZN(n512) );
  XNOR2_X2 U608 ( .A(n512), .B(KEYINPUT33), .ZN(n592) );
  NAND2_X1 U609 ( .A1(n513), .A2(n592), .ZN(n514) );
  NAND2_X1 U610 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U611 ( .A(n516), .B(KEYINPUT52), .ZN(n517) );
  XNOR2_X1 U612 ( .A(n517), .B(KEYINPUT115), .ZN(n518) );
  NOR2_X1 U613 ( .A1(n522), .A2(n518), .ZN(n520) );
  AND2_X1 U614 ( .A1(n592), .A2(n541), .ZN(n519) );
  NOR2_X1 U615 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U616 ( .A(KEYINPUT116), .B(n521), .ZN(n632) );
  NOR2_X1 U617 ( .A1(G953), .A2(n522), .ZN(n585) );
  NAND2_X1 U618 ( .A1(G902), .A2(n523), .ZN(n583) );
  OR2_X1 U619 ( .A1(n733), .A2(n583), .ZN(n524) );
  NOR2_X1 U620 ( .A1(G900), .A2(n524), .ZN(n525) );
  NOR2_X1 U621 ( .A1(n585), .A2(n525), .ZN(n537) );
  NAND2_X1 U622 ( .A1(n526), .A2(n564), .ZN(n528) );
  OR2_X1 U623 ( .A1(n357), .A2(n532), .ZN(n533) );
  XNOR2_X1 U624 ( .A(n533), .B(KEYINPUT99), .ZN(n613) );
  INV_X1 U625 ( .A(KEYINPUT39), .ZN(n534) );
  XNOR2_X1 U626 ( .A(n535), .B(n534), .ZN(n579) );
  NAND2_X1 U627 ( .A1(n579), .A2(n706), .ZN(n536) );
  NOR2_X1 U628 ( .A1(n609), .A2(n537), .ZN(n538) );
  NAND2_X1 U629 ( .A1(n538), .A2(n597), .ZN(n561) );
  NOR2_X1 U630 ( .A1(n561), .A2(n612), .ZN(n539) );
  XOR2_X1 U631 ( .A(KEYINPUT28), .B(n539), .Z(n540) );
  NOR2_X1 U632 ( .A1(n540), .A2(n357), .ZN(n557) );
  NAND2_X1 U633 ( .A1(n541), .A2(n557), .ZN(n542) );
  XNOR2_X1 U634 ( .A(n542), .B(KEYINPUT42), .ZN(n742) );
  NAND2_X1 U635 ( .A1(n744), .A2(n742), .ZN(n544) );
  INV_X1 U636 ( .A(n545), .ZN(n548) );
  OR2_X1 U637 ( .A1(n547), .A2(n546), .ZN(n595) );
  NOR2_X1 U638 ( .A1(n548), .A2(n595), .ZN(n549) );
  NAND2_X1 U639 ( .A1(n549), .A2(n471), .ZN(n551) );
  INV_X1 U640 ( .A(n613), .ZN(n550) );
  NOR2_X1 U641 ( .A1(n551), .A2(n550), .ZN(n701) );
  NAND2_X1 U642 ( .A1(n553), .A2(n564), .ZN(n555) );
  INV_X1 U643 ( .A(KEYINPUT19), .ZN(n554) );
  INV_X1 U644 ( .A(n588), .ZN(n556) );
  NAND2_X1 U645 ( .A1(n557), .A2(n556), .ZN(n703) );
  NOR2_X1 U646 ( .A1(n703), .A2(n558), .ZN(n559) );
  XNOR2_X1 U647 ( .A(n559), .B(KEYINPUT47), .ZN(n571) );
  INV_X1 U648 ( .A(n706), .ZN(n702) );
  NOR2_X1 U649 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U650 ( .A(n562), .B(KEYINPUT105), .ZN(n563) );
  NOR2_X1 U651 ( .A1(n702), .A2(n563), .ZN(n565) );
  NAND2_X1 U652 ( .A1(n565), .A2(n564), .ZN(n576) );
  INV_X1 U653 ( .A(n471), .ZN(n566) );
  NOR2_X1 U654 ( .A1(n576), .A2(n566), .ZN(n567) );
  XNOR2_X1 U655 ( .A(n567), .B(n392), .ZN(n568) );
  NAND2_X1 U656 ( .A1(n568), .A2(n451), .ZN(n569) );
  XNOR2_X1 U657 ( .A(n569), .B(KEYINPUT107), .ZN(n740) );
  INV_X1 U658 ( .A(n740), .ZN(n570) );
  AND2_X1 U659 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U660 ( .A(KEYINPUT48), .B(KEYINPUT70), .ZN(n574) );
  XNOR2_X1 U661 ( .A(n575), .B(n574), .ZN(n582) );
  NOR2_X1 U662 ( .A1(n576), .A2(n355), .ZN(n577) );
  XNOR2_X1 U663 ( .A(n577), .B(KEYINPUT43), .ZN(n578) );
  NOR2_X1 U664 ( .A1(n578), .A2(n471), .ZN(n666) );
  NAND2_X1 U665 ( .A1(n579), .A2(n709), .ZN(n712) );
  INV_X1 U666 ( .A(n712), .ZN(n580) );
  NOR2_X1 U667 ( .A1(n666), .A2(n580), .ZN(n581) );
  AND2_X2 U668 ( .A1(n582), .A2(n581), .ZN(n638) );
  NAND2_X1 U669 ( .A1(n638), .A2(KEYINPUT2), .ZN(n624) );
  OR2_X1 U670 ( .A1(n733), .A2(G898), .ZN(n716) );
  NOR2_X1 U671 ( .A1(n583), .A2(n716), .ZN(n584) );
  OR2_X1 U672 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U673 ( .A(n586), .B(KEYINPUT95), .ZN(n587) );
  INV_X1 U674 ( .A(KEYINPUT65), .ZN(n589) );
  INV_X1 U675 ( .A(n615), .ZN(n591) );
  NAND2_X1 U676 ( .A1(n592), .A2(n591), .ZN(n594) );
  INV_X1 U677 ( .A(KEYINPUT34), .ZN(n593) );
  INV_X1 U678 ( .A(n595), .ZN(n596) );
  NAND2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U680 ( .A(n600), .B(KEYINPUT22), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n560), .A2(n602), .ZN(n603) );
  NOR2_X1 U682 ( .A1(n603), .A2(n409), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n606), .A2(n604), .ZN(n605) );
  NOR2_X1 U684 ( .A1(n526), .A2(n609), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n361), .A2(n607), .ZN(n664) );
  OR2_X1 U686 ( .A1(n615), .A2(n610), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U689 ( .A(KEYINPUT85), .B(KEYINPUT45), .Z(n622) );
  XNOR2_X1 U690 ( .A(n623), .B(n622), .ZN(n636) );
  XNOR2_X1 U691 ( .A(n625), .B(KEYINPUT83), .ZN(n628) );
  INV_X1 U692 ( .A(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U693 ( .A1(n718), .A2(n626), .ZN(n627) );
  NAND2_X1 U694 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U695 ( .A1(n643), .A2(n629), .ZN(n630) );
  NOR2_X1 U696 ( .A1(G953), .A2(n630), .ZN(n631) );
  NAND2_X1 U697 ( .A1(n632), .A2(n631), .ZN(n634) );
  XNOR2_X1 U698 ( .A(KEYINPUT117), .B(KEYINPUT53), .ZN(n633) );
  XNOR2_X1 U699 ( .A(n637), .B(KEYINPUT84), .ZN(n639) );
  NAND2_X1 U700 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U701 ( .A1(n640), .A2(KEYINPUT2), .ZN(n641) );
  INV_X1 U702 ( .A(n643), .ZN(n644) );
  NAND2_X1 U703 ( .A1(n682), .A2(G475), .ZN(n650) );
  XNOR2_X1 U704 ( .A(KEYINPUT89), .B(KEYINPUT122), .ZN(n646) );
  XOR2_X1 U705 ( .A(n646), .B(KEYINPUT59), .Z(n647) );
  XNOR2_X1 U706 ( .A(n650), .B(n649), .ZN(n652) );
  INV_X1 U707 ( .A(G952), .ZN(n651) );
  NAND2_X1 U708 ( .A1(n651), .A2(G953), .ZN(n689) );
  NAND2_X1 U709 ( .A1(n652), .A2(n689), .ZN(n654) );
  XNOR2_X1 U710 ( .A(n654), .B(n653), .ZN(G60) );
  NAND2_X1 U711 ( .A1(n356), .A2(G210), .ZN(n659) );
  XNOR2_X1 U712 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n656) );
  XNOR2_X1 U713 ( .A(n656), .B(KEYINPUT55), .ZN(n657) );
  XNOR2_X1 U714 ( .A(n655), .B(n657), .ZN(n658) );
  XNOR2_X1 U715 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U716 ( .A1(n660), .A2(n689), .ZN(n662) );
  INV_X1 U717 ( .A(KEYINPUT56), .ZN(n661) );
  XNOR2_X1 U718 ( .A(n662), .B(n661), .ZN(G51) );
  XOR2_X1 U719 ( .A(G110), .B(KEYINPUT109), .Z(n663) );
  XNOR2_X1 U720 ( .A(n664), .B(n663), .ZN(G12) );
  XNOR2_X1 U721 ( .A(n666), .B(n665), .ZN(G42) );
  XNOR2_X1 U722 ( .A(n667), .B(G119), .ZN(G21) );
  XOR2_X1 U723 ( .A(n668), .B(G122), .Z(G24) );
  NAND2_X1 U724 ( .A1(n682), .A2(G472), .ZN(n671) );
  XNOR2_X1 U725 ( .A(n669), .B(KEYINPUT62), .ZN(n670) );
  XNOR2_X1 U726 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U727 ( .A1(n672), .A2(n689), .ZN(n673) );
  XNOR2_X1 U728 ( .A(n673), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U729 ( .A1(n356), .A2(G217), .ZN(n676) );
  XNOR2_X1 U730 ( .A(n674), .B(KEYINPUT123), .ZN(n675) );
  XNOR2_X1 U731 ( .A(n676), .B(n675), .ZN(n677) );
  INV_X1 U732 ( .A(n689), .ZN(n680) );
  NOR2_X1 U733 ( .A1(n677), .A2(n680), .ZN(G66) );
  NAND2_X1 U734 ( .A1(n356), .A2(G478), .ZN(n678) );
  XOR2_X1 U735 ( .A(n679), .B(n678), .Z(n681) );
  NOR2_X1 U736 ( .A1(n681), .A2(n680), .ZN(G63) );
  NAND2_X1 U737 ( .A1(n682), .A2(G469), .ZN(n688) );
  XOR2_X1 U738 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n685) );
  XNOR2_X1 U739 ( .A(KEYINPUT120), .B(KEYINPUT119), .ZN(n684) );
  XNOR2_X1 U740 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U741 ( .A(n683), .B(n686), .ZN(n687) );
  XNOR2_X1 U742 ( .A(n688), .B(n687), .ZN(n690) );
  NAND2_X1 U743 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U744 ( .A(n691), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U745 ( .A1(n359), .A2(n706), .ZN(n692) );
  XNOR2_X1 U746 ( .A(n692), .B(G104), .ZN(G6) );
  XNOR2_X1 U747 ( .A(G107), .B(KEYINPUT108), .ZN(n696) );
  XOR2_X1 U748 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n694) );
  NAND2_X1 U749 ( .A1(n359), .A2(n709), .ZN(n693) );
  XNOR2_X1 U750 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U751 ( .A(n696), .B(n695), .ZN(G9) );
  NOR2_X1 U752 ( .A1(n703), .A2(n697), .ZN(n699) );
  XNOR2_X1 U753 ( .A(KEYINPUT110), .B(KEYINPUT29), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U755 ( .A(G128), .B(n700), .ZN(G30) );
  XOR2_X1 U756 ( .A(G143), .B(n701), .Z(G45) );
  NOR2_X1 U757 ( .A1(n703), .A2(n702), .ZN(n705) );
  XNOR2_X1 U758 ( .A(G146), .B(KEYINPUT111), .ZN(n704) );
  XNOR2_X1 U759 ( .A(n705), .B(n704), .ZN(G48) );
  NAND2_X1 U760 ( .A1(n710), .A2(n706), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n707), .B(KEYINPUT112), .ZN(n708) );
  XNOR2_X1 U762 ( .A(G113), .B(n708), .ZN(G15) );
  NAND2_X1 U763 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U764 ( .A(n711), .B(G116), .ZN(G18) );
  XNOR2_X1 U765 ( .A(G134), .B(n712), .ZN(G36) );
  XOR2_X1 U766 ( .A(n713), .B(G101), .Z(n714) );
  XNOR2_X1 U767 ( .A(n715), .B(n714), .ZN(n717) );
  NAND2_X1 U768 ( .A1(n717), .A2(n716), .ZN(n726) );
  INV_X1 U769 ( .A(n718), .ZN(n719) );
  NAND2_X1 U770 ( .A1(n719), .A2(n733), .ZN(n724) );
  NAND2_X1 U771 ( .A1(G224), .A2(G953), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n720), .B(KEYINPUT61), .ZN(n721) );
  XNOR2_X1 U773 ( .A(KEYINPUT124), .B(n721), .ZN(n722) );
  NAND2_X1 U774 ( .A1(G898), .A2(n722), .ZN(n723) );
  NAND2_X1 U775 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U776 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U777 ( .A(KEYINPUT125), .B(n727), .ZN(G69) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U779 ( .A(n730), .B(KEYINPUT126), .ZN(n732) );
  XOR2_X1 U780 ( .A(n732), .B(n731), .Z(n735) );
  XNOR2_X1 U781 ( .A(n638), .B(n735), .ZN(n734) );
  NAND2_X1 U782 ( .A1(n734), .A2(n733), .ZN(n739) );
  XOR2_X1 U783 ( .A(G227), .B(n735), .Z(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U785 ( .A1(n737), .A2(G953), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n739), .A2(n738), .ZN(G72) );
  XNOR2_X1 U787 ( .A(G125), .B(n740), .ZN(n741) );
  XNOR2_X1 U788 ( .A(n741), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U789 ( .A(G137), .B(n742), .Z(n743) );
  XNOR2_X1 U790 ( .A(KEYINPUT127), .B(n743), .ZN(G39) );
  XNOR2_X1 U791 ( .A(G131), .B(n744), .ZN(G33) );
endmodule

