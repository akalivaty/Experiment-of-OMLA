//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G227), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT4), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G101), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n197), .A2(KEYINPUT83), .A3(new_n198), .A4(G101), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n192), .A2(new_n195), .A3(new_n203), .A4(new_n196), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n198), .B1(new_n197), .B2(G101), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n201), .A2(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n207), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(KEYINPUT0), .A3(G128), .A4(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n208), .A2(new_n210), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n207), .A2(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT0), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT65), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT65), .B1(new_n220), .B2(new_n221), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n219), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n206), .A2(new_n215), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n216), .B1(new_n208), .B2(new_n210), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n230));
  OAI21_X1  g044(.A(G128), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n219), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT67), .B(G146), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n214), .B(new_n233), .C1(new_n234), .C2(new_n216), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n196), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n191), .A2(G107), .ZN(new_n238));
  OAI21_X1  g052(.A(G101), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n204), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(KEYINPUT10), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n235), .A2(KEYINPUT84), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT84), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n212), .A2(new_n245), .A3(new_n214), .A4(new_n233), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n230), .B1(G143), .B2(new_n207), .ZN(new_n247));
  OAI22_X1  g061(.A1(new_n229), .A2(new_n213), .B1(new_n221), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n241), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT10), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n243), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AOI211_X1 g066(.A(KEYINPUT85), .B(KEYINPUT10), .C1(new_n249), .C2(new_n241), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n228), .B(new_n242), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT11), .A3(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n259), .A3(new_n263), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n190), .B1(new_n254), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT89), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n229), .A2(new_n213), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n231), .A2(new_n219), .B1(new_n269), .B2(new_n233), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n240), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n250), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT12), .A3(new_n265), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT86), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(new_n265), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT12), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n272), .A2(KEYINPUT86), .A3(KEYINPUT12), .A4(new_n265), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT89), .B(new_n190), .C1(new_n254), .C2(new_n265), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n268), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n190), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n250), .A2(new_n251), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT85), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n250), .A2(new_n243), .A3(new_n251), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n265), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n228), .A4(new_n242), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n254), .A2(new_n265), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n283), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n282), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  INV_X1    g108(.A(G469), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n295), .A2(KEYINPUT88), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(KEYINPUT88), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n293), .A2(new_n294), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n280), .A2(new_n289), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT87), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n280), .A2(new_n289), .A3(KEYINPUT87), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n283), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n291), .A2(new_n266), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n298), .B1(new_n306), .B2(new_n295), .ZN(new_n307));
  INV_X1    g121(.A(G221), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT9), .B(G234), .Z(new_n309));
  AOI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(new_n294), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G113), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n313), .A2(KEYINPUT2), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(KEYINPUT2), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT68), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT2), .B(G113), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(G116), .B(G119), .Z(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT69), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n320), .A2(new_n317), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT69), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n316), .A2(new_n319), .A3(new_n324), .A4(new_n320), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n206), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT5), .ZN(new_n328));
  INV_X1    g142(.A(G119), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(G116), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n320), .B2(new_n328), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n323), .B1(new_n331), .B2(new_n313), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n332), .A2(new_n240), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G122), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n332), .A2(new_n240), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n206), .B2(new_n326), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n335), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n340), .A3(KEYINPUT6), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n227), .A2(new_n215), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT79), .B(G125), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT90), .ZN(new_n345));
  INV_X1    g159(.A(new_n343), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n344), .A2(new_n345), .B1(new_n270), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G224), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(G953), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n347), .B(new_n350), .C1(new_n345), .C2(new_n344), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n346), .B1(new_n227), .B2(new_n215), .ZN(new_n352));
  OAI22_X1  g166(.A1(new_n352), .A2(KEYINPUT90), .B1(new_n236), .B2(new_n343), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n344), .A2(new_n345), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n349), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n334), .A2(new_n357), .A3(new_n336), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n341), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n335), .B(KEYINPUT8), .Z(new_n360));
  NAND2_X1  g174(.A1(new_n332), .A2(new_n240), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n333), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n339), .B2(new_n335), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT7), .ZN(new_n364));
  OAI22_X1  g178(.A1(new_n353), .A2(new_n354), .B1(new_n364), .B2(new_n349), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n363), .B(new_n365), .C1(new_n364), .C2(new_n351), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n359), .A2(new_n366), .A3(new_n294), .ZN(new_n367));
  OAI21_X1  g181(.A(G210), .B1(G237), .B2(G902), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(KEYINPUT91), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n369), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n359), .A2(new_n366), .A3(new_n294), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(G214), .B1(G237), .B2(G902), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G475), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT16), .ZN(new_n377));
  INV_X1    g191(.A(G140), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n343), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G125), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n378), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n343), .B2(G140), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n379), .B1(new_n383), .B2(new_n377), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n207), .ZN(new_n385));
  NOR2_X1   g199(.A1(G237), .A2(G953), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G214), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n216), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(G143), .A3(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G131), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT17), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(new_n263), .A3(new_n389), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(G146), .B(new_n379), .C1(new_n383), .C2(new_n377), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n390), .A2(KEYINPUT17), .A3(G131), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n385), .A2(new_n394), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n343), .A2(G140), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(G146), .A3(new_n381), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(G125), .A2(G140), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n381), .A2(KEYINPUT80), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT80), .B1(new_n381), .B2(new_n402), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n211), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n383), .A2(KEYINPUT92), .A3(G146), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT18), .A2(G131), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n390), .B(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n397), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G113), .B(G122), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(new_n191), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n397), .A2(new_n410), .A3(new_n413), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n376), .B1(new_n417), .B2(new_n294), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT19), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n403), .B2(new_n404), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n398), .A2(KEYINPUT19), .A3(new_n381), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n421), .A3(new_n211), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT93), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n391), .A2(new_n393), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT93), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n420), .A2(new_n421), .A3(new_n425), .A4(new_n211), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n423), .A2(new_n395), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n410), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n414), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n416), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n430), .A2(new_n431), .A3(new_n376), .A4(new_n294), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n413), .B1(new_n427), .B2(new_n410), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n397), .A2(new_n410), .A3(new_n413), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n376), .B(new_n294), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT20), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n418), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G952), .ZN(new_n438));
  AOI211_X1 g252(.A(G953), .B(new_n438), .C1(G234), .C2(G237), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT21), .B(G898), .Z(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n294), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n309), .A2(G217), .A3(new_n188), .ZN(new_n445));
  INV_X1    g259(.A(G122), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G116), .ZN(new_n447));
  INV_X1    g261(.A(G116), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G122), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G107), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n449), .A3(new_n194), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n216), .A2(G128), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n221), .A2(G143), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT13), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n456), .B(G134), .C1(KEYINPUT13), .C2(new_n454), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n455), .A3(new_n256), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n453), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n454), .A2(new_n455), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G134), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n458), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n448), .A2(KEYINPUT14), .A3(G122), .ZN(new_n463));
  OAI211_X1 g277(.A(G107), .B(new_n463), .C1(new_n450), .C2(KEYINPUT14), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n452), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT94), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n459), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n466), .B1(new_n459), .B2(new_n465), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n445), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n459), .A2(new_n465), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT94), .ZN(new_n472));
  INV_X1    g286(.A(new_n445), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n467), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n474), .A3(new_n294), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n477), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n437), .A2(new_n444), .A3(new_n481), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n312), .A2(new_n375), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT29), .ZN(new_n484));
  XOR2_X1   g298(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n326), .ZN(new_n487));
  INV_X1    g301(.A(new_n260), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n256), .A2(G137), .ZN(new_n489));
  OAI21_X1  g303(.A(G131), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n264), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n232), .B2(new_n235), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n265), .A2(new_n227), .A3(new_n215), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n487), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n494), .B1(new_n270), .B2(new_n491), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n326), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n486), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n496), .A2(new_n326), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(KEYINPUT28), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n386), .A2(G210), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(new_n203), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n498), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n505), .A2(KEYINPUT73), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT64), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n265), .A2(new_n227), .A3(new_n215), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n507), .B1(new_n492), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT70), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT30), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n496), .B2(KEYINPUT70), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT70), .B1(new_n496), .B2(new_n507), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n511), .B(new_n326), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n495), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n505), .B1(new_n516), .B2(new_n504), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT73), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n484), .B(new_n506), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n495), .A2(new_n497), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT28), .ZN(new_n522));
  INV_X1    g336(.A(new_n500), .ZN(new_n523));
  INV_X1    g337(.A(new_n504), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT29), .A4(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n525), .A2(KEYINPUT75), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(KEYINPUT75), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n526), .A2(new_n527), .A3(G902), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n524), .B1(new_n515), .B2(new_n495), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT73), .B1(new_n529), .B2(new_n505), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT74), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n484), .A4(new_n506), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n520), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G472), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT32), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n504), .B1(new_n498), .B2(new_n500), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n515), .A2(new_n524), .A3(new_n495), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT31), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n515), .A2(KEYINPUT31), .A3(new_n524), .A4(new_n495), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(G472), .A2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n535), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT72), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT72), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n540), .A2(new_n541), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n536), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT32), .B1(new_n549), .B2(new_n543), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n542), .A2(new_n535), .A3(new_n544), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n534), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT22), .B(G137), .ZN(new_n554));
  INV_X1    g368(.A(G234), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n308), .A2(new_n555), .A3(G953), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n554), .B(new_n556), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n385), .A2(new_n395), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n329), .A2(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT78), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n221), .A2(G119), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT78), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT23), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n221), .A2(G119), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n561), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT77), .B1(new_n562), .B2(new_n565), .ZN(new_n568));
  OR3_X1    g382(.A1(new_n562), .A2(KEYINPUT77), .A3(new_n565), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n566), .A2(new_n560), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT24), .B(G110), .Z(new_n572));
  AOI22_X1  g386(.A1(new_n570), .A2(G110), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n559), .A2(new_n573), .ZN(new_n574));
  OAI22_X1  g388(.A1(new_n570), .A2(G110), .B1(new_n571), .B2(new_n572), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n395), .A3(new_n405), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n574), .A2(new_n576), .A3(KEYINPUT81), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT81), .B1(new_n574), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n558), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(new_n576), .A3(new_n557), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n294), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT25), .ZN(new_n582));
  OAI21_X1  g396(.A(G217), .B1(new_n555), .B2(G902), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT76), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT25), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n579), .A2(new_n586), .A3(new_n294), .A4(new_n580), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n582), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n579), .A2(new_n580), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n585), .A2(G902), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n588), .A2(new_n591), .A3(KEYINPUT82), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT82), .B1(new_n588), .B2(new_n591), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n483), .A2(new_n553), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  OR2_X1    g410(.A1(new_n367), .A2(new_n368), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n367), .A2(new_n368), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n374), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n190), .B1(new_n299), .B2(new_n300), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n304), .B1(new_n600), .B2(new_n302), .ZN(new_n601));
  OAI21_X1  g415(.A(G469), .B1(new_n601), .B2(G902), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n310), .B(new_n599), .C1(new_n602), .C2(new_n298), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n549), .A2(new_n543), .ZN(new_n604));
  OAI21_X1  g418(.A(G472), .B1(new_n542), .B2(G902), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n604), .B(new_n605), .C1(new_n592), .C2(new_n593), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n475), .A2(new_n476), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n468), .A2(new_n469), .A3(new_n445), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n473), .B1(new_n472), .B2(new_n467), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n470), .A2(new_n474), .A3(KEYINPUT33), .ZN(new_n614));
  AOI21_X1  g428(.A(G902), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n609), .B1(new_n615), .B2(G478), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n437), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n443), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n603), .A2(new_n607), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  NOR2_X1   g436(.A1(new_n312), .A2(new_n606), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n432), .A2(KEYINPUT95), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n432), .A2(KEYINPUT95), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n436), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n481), .A2(new_n418), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n599), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n623), .A2(new_n444), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G107), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT96), .B(KEYINPUT35), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n604), .A2(new_n605), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n577), .A2(new_n578), .ZN(new_n636));
  OR2_X1    g450(.A1(new_n558), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n590), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n588), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n634), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT97), .A4(new_n640), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n483), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n442), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n439), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n310), .B(new_n651), .C1(new_n602), .C2(new_n298), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n553), .A2(new_n629), .A3(new_n640), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  AOI21_X1  g468(.A(new_n310), .B1(new_n602), .B2(new_n298), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n650), .B(KEYINPUT39), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT40), .ZN(new_n658));
  INV_X1    g472(.A(new_n521), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n538), .B1(new_n524), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G472), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n552), .A2(new_n546), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n437), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n665), .A2(new_n374), .A3(new_n480), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT99), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n373), .B(new_n669), .Z(new_n670));
  NOR4_X1   g484(.A1(new_n658), .A2(new_n640), .A3(new_n667), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n216), .ZN(G45));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n617), .B2(new_n650), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n437), .A2(new_n616), .A3(KEYINPUT101), .A4(new_n651), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n553), .A2(new_n603), .A3(new_n640), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  NAND2_X1  g492(.A1(new_n293), .A2(new_n294), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n298), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n681), .A2(new_n310), .A3(new_n599), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n553), .A2(new_n682), .A3(new_n594), .A4(new_n619), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NOR3_X1   g499(.A1(new_n681), .A2(new_n310), .A3(new_n443), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n553), .A2(new_n686), .A3(new_n594), .A4(new_n629), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  INV_X1    g502(.A(new_n482), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n553), .A2(new_n682), .A3(new_n689), .A4(new_n640), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  AND2_X1   g505(.A1(new_n588), .A2(new_n591), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n599), .A2(new_n481), .A3(new_n437), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n522), .A2(new_n523), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n504), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n544), .B1(new_n548), .B2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n605), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g512(.A(KEYINPUT102), .B(G472), .C1(new_n542), .C2(G902), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n686), .A2(new_n692), .A3(new_n693), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  NAND4_X1  g516(.A1(new_n682), .A2(new_n640), .A3(new_n676), .A4(new_n700), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G125), .ZN(G27));
  NAND3_X1  g518(.A1(new_n370), .A2(new_n374), .A3(new_n372), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n674), .A2(new_n675), .A3(new_n705), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n655), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n553), .A3(new_n594), .ZN(new_n708));
  NAND2_X1  g522(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n709));
  OR2_X1    g523(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  OR3_X1    g525(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT104), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT104), .B1(new_n550), .B2(new_n551), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n534), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n707), .A3(KEYINPUT42), .A4(new_n692), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G131), .ZN(G33));
  INV_X1    g531(.A(new_n628), .ZN(new_n718));
  AND4_X1   g532(.A1(new_n311), .A2(new_n307), .A3(new_n718), .A4(new_n650), .ZN(new_n719));
  INV_X1    g533(.A(new_n705), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n553), .A3(new_n594), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  OAI21_X1  g536(.A(G469), .B1(new_n601), .B2(KEYINPUT45), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n601), .A2(KEYINPUT45), .ZN(new_n726));
  OAI211_X1 g540(.A(KEYINPUT105), .B(G469), .C1(new_n601), .C2(KEYINPUT45), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(G469), .A2(G902), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n728), .A2(KEYINPUT46), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT46), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  INV_X1    g545(.A(new_n298), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n310), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n635), .A2(new_n640), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n735), .A2(KEYINPUT106), .ZN(new_n736));
  INV_X1    g550(.A(new_n616), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n437), .ZN(new_n738));
  XOR2_X1   g552(.A(new_n738), .B(KEYINPUT43), .Z(new_n739));
  NAND2_X1  g553(.A1(new_n735), .A2(KEYINPUT106), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n736), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AND4_X1   g558(.A1(new_n656), .A2(new_n734), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n705), .B(KEYINPUT107), .Z(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G137), .ZN(G39));
  XNOR2_X1  g563(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n733), .B2(new_n310), .ZN(new_n752));
  INV_X1    g566(.A(new_n553), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n728), .A2(new_n729), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n728), .A2(KEYINPUT46), .A3(new_n729), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n298), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n311), .A3(new_n750), .ZN(new_n759));
  INV_X1    g573(.A(new_n706), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n594), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n752), .A2(new_n753), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  INV_X1    g579(.A(new_n670), .ZN(new_n766));
  INV_X1    g580(.A(new_n738), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n692), .A2(new_n767), .A3(new_n374), .A4(new_n311), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT110), .Z(new_n769));
  INV_X1    g583(.A(new_n665), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n769), .B(new_n770), .C1(KEYINPUT49), .C2(new_n681), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n766), .B(new_n771), .C1(KEYINPUT49), .C2(new_n681), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(KEYINPUT111), .Z(new_n773));
  NAND4_X1  g587(.A1(new_n665), .A2(new_n652), .A3(new_n641), .A4(new_n693), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT115), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n653), .A2(new_n677), .A3(new_n703), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT52), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n549), .A2(KEYINPUT32), .A3(new_n543), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT72), .B1(new_n778), .B2(new_n545), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n547), .B1(new_n604), .B2(new_n535), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n640), .B1(new_n781), .B2(new_n664), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(KEYINPUT115), .A3(new_n652), .A4(new_n693), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n774), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n653), .A2(new_n677), .A3(new_n703), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n721), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n711), .B2(new_n715), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n480), .A2(new_n418), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n720), .A2(new_n626), .A3(new_n650), .A4(new_n793), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(KEYINPUT113), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(KEYINPUT113), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n553), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n700), .A2(new_n706), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n655), .B(new_n640), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n618), .B(KEYINPUT112), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n432), .A2(new_n436), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n627), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n375), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n623), .A2(new_n803), .A3(new_n804), .A4(new_n444), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n595), .A2(new_n644), .A3(new_n805), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n683), .A2(new_n687), .A3(new_n690), .A4(new_n701), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n792), .A2(new_n799), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n790), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n788), .B1(new_n786), .B2(new_n787), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n595), .A2(new_n644), .A3(new_n805), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n683), .A2(new_n687), .A3(new_n690), .A4(new_n701), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n799), .A4(new_n792), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n810), .A2(new_n813), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n809), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n739), .A2(new_n439), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n681), .A2(new_n310), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n824), .A2(new_n825), .A3(new_n720), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n714), .A2(new_n692), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT48), .Z(new_n829));
  NOR3_X1   g643(.A1(new_n829), .A2(new_n438), .A3(G953), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n810), .A2(new_n818), .ZN(new_n831));
  INV_X1    g645(.A(new_n790), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n831), .A2(new_n832), .B1(new_n819), .B2(new_n820), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n823), .B(new_n830), .C1(new_n822), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n752), .A2(new_n759), .ZN(new_n835));
  INV_X1    g649(.A(new_n681), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n310), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n700), .A2(new_n692), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n824), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n747), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n825), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n840), .A2(new_n374), .A3(new_n766), .A4(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT50), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n665), .A2(new_n649), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n594), .A3(new_n825), .A4(new_n720), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n847), .A2(new_n666), .A3(new_n737), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n826), .A2(new_n640), .A3(new_n700), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n842), .A2(new_n845), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n842), .A2(KEYINPUT116), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n842), .A2(new_n845), .A3(new_n848), .A4(new_n849), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n852), .A3(new_n851), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n847), .A2(new_n618), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n840), .A2(new_n599), .A3(new_n843), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n834), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(G952), .A2(G953), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n773), .B1(new_n860), .B2(new_n861), .ZN(G75));
  NAND2_X1  g676(.A1(new_n341), .A2(new_n358), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(new_n356), .Z(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT55), .ZN(new_n865));
  INV_X1    g679(.A(G210), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n821), .A2(new_n866), .A3(new_n294), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n865), .B1(new_n867), .B2(KEYINPUT56), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n188), .A2(G952), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n819), .A2(new_n820), .ZN(new_n871));
  INV_X1    g685(.A(new_n809), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(G210), .A3(G902), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT56), .ZN(new_n875));
  INV_X1    g689(.A(new_n865), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n868), .A2(new_n870), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT117), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n868), .A2(new_n877), .A3(new_n880), .A4(new_n870), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(G51));
  NAND2_X1  g696(.A1(new_n729), .A2(KEYINPUT57), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n729), .A2(KEYINPUT57), .ZN(new_n884));
  INV_X1    g698(.A(new_n823), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n821), .A2(new_n822), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n883), .B(new_n884), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n293), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n821), .A2(new_n294), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n728), .B(KEYINPUT118), .Z(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n869), .B1(new_n888), .B2(new_n891), .ZN(G54));
  NAND3_X1  g706(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .ZN(new_n893));
  INV_X1    g707(.A(new_n430), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n895), .A2(new_n896), .A3(new_n869), .ZN(G60));
  XNOR2_X1  g711(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n476), .A2(new_n294), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n898), .B(new_n899), .Z(new_n900));
  NAND2_X1  g714(.A1(new_n613), .A2(new_n614), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT119), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n900), .B(new_n902), .C1(new_n885), .C2(new_n886), .ZN(new_n903));
  INV_X1    g717(.A(new_n900), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n831), .A2(new_n832), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n871), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n904), .B1(new_n907), .B2(new_n823), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n903), .B(new_n870), .C1(new_n908), .C2(new_n902), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(G63));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT60), .Z(new_n912));
  XNOR2_X1  g726(.A(new_n638), .B(KEYINPUT121), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n873), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n873), .A2(new_n912), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n870), .B(new_n914), .C1(new_n915), .C2(new_n589), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT61), .B1(new_n914), .B2(KEYINPUT122), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(G66));
  OAI21_X1  g732(.A(G953), .B1(new_n441), .B2(new_n348), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n816), .B2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n863), .B1(G898), .B2(new_n188), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(G69));
  AOI21_X1  g736(.A(new_n776), .B1(new_n745), .B2(new_n747), .ZN(new_n923));
  INV_X1    g737(.A(new_n792), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n734), .A2(new_n656), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n827), .A2(new_n693), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n764), .A2(new_n923), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n513), .A2(new_n514), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(KEYINPUT30), .B2(new_n514), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n420), .A2(new_n421), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n930), .B(new_n931), .Z(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(G953), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n671), .A2(new_n776), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT62), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n553), .A2(new_n594), .A3(new_n720), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n657), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n745), .A2(new_n747), .B1(new_n803), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n764), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n934), .B1(new_n933), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(G900), .B1(KEYINPUT123), .B2(G227), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n933), .B(new_n942), .C1(KEYINPUT123), .C2(G900), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n932), .A2(G227), .A3(G900), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(G953), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n941), .A2(new_n945), .ZN(G72));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n764), .A2(new_n816), .A3(new_n923), .A4(new_n927), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n949));
  NAND2_X1  g763(.A1(G472), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n948), .A2(KEYINPUT125), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT125), .B1(new_n948), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n516), .A2(new_n524), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT126), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n952), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n764), .A2(new_n816), .A3(new_n936), .A4(new_n939), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n951), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n504), .B1(new_n515), .B2(new_n495), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n954), .A2(new_n960), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n906), .A2(new_n951), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n961), .A2(new_n870), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n947), .B1(new_n957), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n948), .A2(new_n951), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n948), .A2(KEYINPUT125), .A3(new_n951), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n969), .A3(new_n955), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n869), .B1(new_n959), .B2(new_n960), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n970), .A2(KEYINPUT127), .A3(new_n963), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n965), .A2(new_n972), .ZN(G57));
endmodule


