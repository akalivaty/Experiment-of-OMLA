//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946;
  NAND2_X1  g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT14), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT87), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n203), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NOR3_X1   g008(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(KEYINPUT87), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n202), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(KEYINPUT15), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n207), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n210), .A2(KEYINPUT88), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(new_n203), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n213), .A2(KEYINPUT15), .B1(KEYINPUT89), .B2(new_n202), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n202), .A2(KEYINPUT89), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n214), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT90), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G15gat), .B(G22gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT16), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(G1gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n230), .B(new_n231), .C1(G1gat), .C2(new_n228), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n227), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n234), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n223), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n235), .A2(KEYINPUT18), .A3(new_n236), .A4(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n234), .B(new_n223), .Z(new_n240));
  XOR2_X1   g039(.A(new_n236), .B(KEYINPUT13), .Z(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT18), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT92), .ZN(new_n248));
  XNOR2_X1  g047(.A(G169gat), .B(G197gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G113gat), .B(G141gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT12), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n244), .B(new_n247), .C1(new_n248), .C2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n254), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n248), .A3(new_n242), .ZN(new_n257));
  INV_X1    g056(.A(new_n247), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n256), .B(new_n257), .C1(new_n258), .C2(new_n243), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT100), .ZN(new_n261));
  INV_X1    g060(.A(G57gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(KEYINPUT93), .ZN(new_n263));
  INV_X1    g062(.A(G64gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G71gat), .A2(G78gat), .ZN(new_n266));
  OR2_X1    g065(.A1(G71gat), .A2(G78gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT9), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT9), .B1(new_n262), .B2(new_n264), .ZN(new_n271));
  NOR2_X1   g070(.A1(G57gat), .A2(G64gat), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n266), .B(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(KEYINPUT21), .ZN(new_n275));
  XNOR2_X1  g074(.A(G127gat), .B(G155gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G211gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n275), .B(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G183gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(KEYINPUT21), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n234), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n281), .B1(new_n234), .B2(new_n282), .ZN(new_n285));
  INV_X1    g084(.A(G231gat), .ZN(new_n286));
  INV_X1    g085(.A(G233gat), .ZN(new_n287));
  OAI22_X1  g086(.A1(new_n284), .A2(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n234), .A2(new_n282), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G183gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n286), .A2(new_n287), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n283), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n288), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n288), .B2(new_n292), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n280), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n288), .A2(new_n292), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n293), .ZN(new_n300));
  INV_X1    g099(.A(new_n279), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n278), .B(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n302), .A3(new_n295), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(G85gat), .A2(G92gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT7), .ZN(new_n308));
  NOR2_X1   g107(.A1(G85gat), .A2(G92gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(G99gat), .A2(G106gat), .ZN(new_n310));
  AOI211_X1 g109(.A(KEYINPUT97), .B(new_n309), .C1(KEYINPUT8), .C2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G85gat), .ZN(new_n312));
  INV_X1    g111(.A(G92gat), .ZN(new_n313));
  AOI22_X1  g112(.A1(KEYINPUT8), .A2(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT97), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n308), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G99gat), .B(G106gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n318), .B(new_n308), .C1(new_n311), .C2(new_n316), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT98), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(KEYINPUT98), .A3(new_n319), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n223), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n225), .B(KEYINPUT17), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n306), .B(new_n326), .C1(new_n327), .C2(new_n325), .ZN(new_n328));
  XNOR2_X1  g127(.A(G134gat), .B(G162gat), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n329), .B(new_n330), .Z(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n227), .A2(new_n324), .A3(new_n323), .ZN(new_n333));
  INV_X1    g132(.A(new_n331), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n306), .A4(new_n326), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT96), .B(KEYINPUT99), .ZN(new_n336));
  XNOR2_X1  g135(.A(G190gat), .B(G218gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n332), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(new_n332), .B2(new_n335), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n261), .B1(new_n305), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n304), .B(KEYINPUT100), .C1(new_n339), .C2(new_n340), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G211gat), .B(G218gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G197gat), .ZN(new_n350));
  INV_X1    g149(.A(G204gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G197gat), .A2(G204gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT22), .ZN(new_n354));
  NAND2_X1  g153(.A1(G211gat), .A2(G218gat), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n352), .A2(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT70), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n349), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n354), .ZN(new_n359));
  NOR2_X1   g158(.A1(G197gat), .A2(G204gat), .ZN(new_n360));
  AND2_X1   g159(.A1(G197gat), .A2(G204gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(KEYINPUT70), .A3(new_n348), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT27), .B1(new_n281), .B2(KEYINPUT65), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT65), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT27), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(G183gat), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT28), .ZN(new_n374));
  INV_X1    g173(.A(G190gat), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n370), .A2(new_n373), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT26), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384));
  AND2_X1   g183(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n375), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n384), .B1(new_n387), .B2(KEYINPUT28), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n380), .A2(KEYINPUT23), .ZN(new_n389));
  INV_X1    g188(.A(G169gat), .ZN(new_n390));
  INV_X1    g189(.A(G176gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n377), .A2(KEYINPUT23), .ZN(new_n394));
  NAND3_X1  g193(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(G183gat), .B2(G190gat), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n393), .B(new_n394), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n383), .A2(new_n388), .B1(KEYINPUT25), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT23), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n400), .A2(G169gat), .A3(G176gat), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n392), .B2(new_n389), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT25), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT64), .B1(new_n384), .B2(KEYINPUT24), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT64), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n402), .B(new_n403), .C1(new_n407), .C2(new_n396), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n369), .B1(new_n399), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n387), .A2(KEYINPUT28), .ZN(new_n410));
  INV_X1    g209(.A(new_n384), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n376), .A4(new_n382), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n398), .A2(KEYINPUT25), .ZN(new_n413));
  AND4_X1   g212(.A1(new_n412), .A2(new_n408), .A3(new_n413), .A4(new_n366), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n365), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT71), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n408), .A3(new_n366), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n408), .A2(new_n413), .A3(new_n412), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n368), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n419), .A3(new_n364), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(KEYINPUT71), .B(new_n365), .C1(new_n409), .C2(new_n414), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n347), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n423), .A2(KEYINPUT30), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n423), .A2(KEYINPUT74), .A3(KEYINPUT30), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT74), .B1(new_n423), .B2(KEYINPUT30), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n421), .A2(KEYINPUT72), .A3(new_n422), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT72), .B1(new_n421), .B2(new_n422), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT73), .B1(new_n430), .B2(new_n347), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT73), .ZN(new_n432));
  INV_X1    g231(.A(new_n347), .ZN(new_n433));
  NOR4_X1   g232(.A1(new_n428), .A2(new_n429), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n427), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n424), .B1(new_n435), .B2(KEYINPUT75), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT79), .ZN(new_n437));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(KEYINPUT5), .ZN(new_n440));
  XNOR2_X1  g239(.A(G155gat), .B(G162gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT2), .ZN(new_n442));
  INV_X1    g241(.A(G148gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(G141gat), .ZN(new_n444));
  INV_X1    g243(.A(G141gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G148gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n441), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G141gat), .B(G148gat), .ZN(new_n449));
  INV_X1    g248(.A(G155gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT76), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT76), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(G155gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n453), .A3(G162gat), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n449), .B1(new_n454), .B2(KEYINPUT2), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n448), .B1(new_n441), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT3), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(KEYINPUT2), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(new_n447), .A3(new_n441), .ZN(new_n460));
  INV_X1    g259(.A(new_n441), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(KEYINPUT2), .B2(new_n449), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT1), .ZN(new_n465));
  INV_X1    g264(.A(G113gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(G120gat), .ZN(new_n467));
  INV_X1    g266(.A(G120gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(G113gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n465), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G127gat), .B(G134gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(G113gat), .B(G120gat), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n470), .B(new_n471), .C1(KEYINPUT66), .C2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(KEYINPUT66), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n472), .A2(KEYINPUT1), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n458), .A2(new_n464), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT4), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n474), .B(new_n470), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n460), .A2(new_n462), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT77), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT77), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n477), .A2(new_n456), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n480), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n477), .A2(new_n456), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n480), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n486), .A2(KEYINPUT78), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT78), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n477), .A2(new_n456), .A3(new_n484), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n484), .B1(new_n477), .B2(new_n456), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT4), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(new_n494), .B2(new_n488), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n440), .B(new_n479), .C1(new_n490), .C2(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n483), .B(new_n485), .C1(new_n480), .C2(new_n439), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n479), .B(new_n497), .C1(new_n480), .C2(new_n487), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n492), .A2(new_n493), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n482), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n439), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(KEYINPUT5), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G1gat), .B(G29gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(G85gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT0), .B(G57gat), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n506), .B(new_n507), .Z(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n437), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n504), .A2(new_n509), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n496), .A2(new_n503), .A3(KEYINPUT79), .A4(new_n508), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n504), .A2(KEYINPUT6), .A3(new_n509), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G78gat), .B(G106gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT31), .B(G50gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G228gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(new_n287), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT80), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n362), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n359), .B(KEYINPUT80), .C1(new_n360), .C2(new_n361), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n349), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n362), .A2(new_n522), .A3(new_n348), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n367), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n457), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n482), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n463), .A2(new_n367), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n365), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n521), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n364), .B1(new_n367), .B2(new_n463), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n358), .A2(new_n367), .A3(new_n363), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n456), .B1(new_n457), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n521), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n519), .B1(new_n538), .B2(G22gat), .ZN(new_n539));
  INV_X1    g338(.A(G22gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n532), .B2(new_n537), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT81), .B1(new_n532), .B2(new_n537), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n534), .A2(new_n457), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n531), .B(new_n521), .C1(new_n456), .C2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n456), .B1(new_n527), .B2(new_n457), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n536), .B1(new_n546), .B2(new_n533), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT81), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n545), .A2(new_n547), .A3(new_n548), .A4(G22gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n541), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n550), .A2(KEYINPUT82), .A3(new_n519), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT82), .B1(new_n550), .B2(new_n519), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n542), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n399), .A2(new_n481), .A3(new_n408), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n418), .A2(new_n477), .ZN(new_n555));
  NAND2_X1  g354(.A1(G227gat), .A2(G233gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT33), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT67), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G15gat), .B(G43gat), .Z(new_n563));
  XNOR2_X1  g362(.A(G71gat), .B(G99gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n558), .A2(KEYINPUT32), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n558), .A2(KEYINPUT67), .A3(new_n559), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n562), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n554), .A2(new_n555), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n556), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT34), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n571), .B1(new_n556), .B2(KEYINPUT68), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n570), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n565), .A2(KEYINPUT33), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n558), .A2(KEYINPUT32), .A3(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n568), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n574), .B1(new_n568), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT69), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT69), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n553), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT75), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n583), .B(new_n427), .C1(new_n431), .C2(new_n434), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n436), .A2(new_n516), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT35), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT85), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n496), .A2(new_n503), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n496), .B2(new_n503), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n509), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n590), .A2(new_n511), .A3(new_n513), .A4(new_n510), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n515), .ZN(new_n592));
  INV_X1    g391(.A(new_n424), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n427), .B(new_n593), .C1(new_n431), .C2(new_n434), .ZN(new_n594));
  INV_X1    g393(.A(new_n553), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT35), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n577), .A2(new_n578), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n592), .A2(new_n596), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n586), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n435), .A2(KEYINPUT75), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n601), .A2(new_n516), .A3(new_n584), .A4(new_n593), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n553), .B(KEYINPUT83), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n421), .A2(new_n422), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n347), .B1(new_n605), .B2(KEYINPUT37), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT37), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n415), .B2(new_n420), .ZN(new_n608));
  OR3_X1    g407(.A1(new_n606), .A2(KEYINPUT38), .A3(new_n608), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n428), .A2(new_n429), .A3(new_n607), .ZN(new_n610));
  OAI22_X1  g409(.A1(new_n610), .A2(new_n606), .B1(KEYINPUT38), .B2(new_n423), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n591), .A2(new_n515), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n499), .A2(new_n438), .A3(new_n500), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT78), .B1(new_n486), .B2(new_n489), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n494), .A2(new_n488), .A3(new_n491), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n478), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g415(.A(KEYINPUT39), .B(new_n613), .C1(new_n616), .C2(new_n438), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n479), .B1(new_n490), .B2(new_n495), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n619), .A3(new_n439), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n508), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n621), .A2(KEYINPUT84), .A3(KEYINPUT40), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT40), .B1(new_n621), .B2(KEYINPUT84), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n590), .B(new_n594), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n612), .A2(new_n624), .A3(new_n553), .ZN(new_n625));
  INV_X1    g424(.A(new_n598), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(KEYINPUT36), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n579), .A2(new_n581), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(KEYINPUT36), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n604), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  AOI211_X1 g429(.A(new_n260), .B(new_n344), .C1(new_n600), .C2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n325), .A2(KEYINPUT10), .A3(new_n274), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT101), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n274), .A2(new_n320), .A3(new_n321), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n635), .B(new_n636), .C1(new_n325), .C2(new_n274), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n325), .A2(KEYINPUT101), .A3(KEYINPUT10), .A4(new_n274), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n636), .B1(new_n325), .B2(new_n274), .ZN(new_n642));
  INV_X1    g441(.A(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n645), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n631), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n516), .B(KEYINPUT102), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT103), .B(G1gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1324gat));
  INV_X1    g454(.A(new_n594), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  OR3_X1    g456(.A1(new_n229), .A2(KEYINPUT104), .A3(KEYINPUT42), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n229), .B1(KEYINPUT104), .B2(KEYINPUT42), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(G8gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(G8gat), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n661), .B(new_n662), .C1(KEYINPUT42), .C2(new_n657), .ZN(G1325gat));
  INV_X1    g462(.A(new_n651), .ZN(new_n664));
  INV_X1    g463(.A(new_n629), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n664), .A2(G15gat), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(G15gat), .B1(new_n664), .B2(new_n598), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(G1326gat));
  INV_X1    g467(.A(new_n603), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n651), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  AOI21_X1  g471(.A(new_n260), .B1(new_n600), .B2(new_n630), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n650), .A2(new_n305), .A3(new_n341), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT105), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(KEYINPUT105), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n673), .A2(new_n205), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n677), .A2(KEYINPUT45), .A3(new_n652), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT45), .B1(new_n677), .B2(new_n652), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n586), .A2(new_n681), .A3(new_n599), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(new_n586), .B2(new_n599), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n630), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT44), .B1(new_n684), .B2(new_n341), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  INV_X1    g485(.A(new_n341), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n686), .B(new_n687), .C1(new_n600), .C2(new_n630), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n650), .A2(new_n305), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n260), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NOR4_X1   g490(.A1(new_n685), .A2(new_n652), .A3(new_n688), .A4(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n680), .B1(new_n692), .B2(new_n205), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT107), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n680), .B(new_n695), .C1(new_n205), .C2(new_n692), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(G36gat), .A3(new_n656), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  NOR4_X1   g499(.A1(new_n685), .A2(new_n656), .A3(new_n691), .A4(new_n688), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(new_n206), .ZN(G1329gat));
  NOR3_X1   g501(.A1(new_n698), .A2(G43gat), .A3(new_n626), .ZN(new_n703));
  INV_X1    g502(.A(new_n630), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n600), .A2(KEYINPUT106), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n586), .A2(new_n681), .A3(new_n599), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n686), .B1(new_n707), .B2(new_n687), .ZN(new_n708));
  INV_X1    g507(.A(new_n688), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n708), .A2(new_n665), .A3(new_n690), .A4(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n703), .B1(new_n710), .B2(G43gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g511(.A1(new_n708), .A2(new_n595), .A3(new_n690), .A4(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT110), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n684), .A2(new_n341), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n688), .B1(new_n715), .B2(new_n686), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n716), .A2(new_n717), .A3(new_n595), .A4(new_n690), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n714), .A2(new_n718), .A3(G50gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n600), .A2(new_n630), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n255), .A2(new_n259), .ZN(new_n721));
  AND4_X1   g520(.A1(new_n720), .A2(new_n721), .A3(new_n675), .A4(new_n676), .ZN(new_n722));
  INV_X1    g521(.A(G50gat), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(new_n723), .A3(new_n603), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n724), .A2(KEYINPUT48), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n722), .A2(KEYINPUT109), .A3(new_n723), .A4(new_n603), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n673), .A2(new_n723), .A3(new_n675), .A4(new_n676), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(new_n669), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NOR4_X1   g530(.A1(new_n685), .A2(new_n669), .A3(new_n688), .A4(new_n691), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(new_n723), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n726), .A2(new_n735), .ZN(G1331gat));
  NOR2_X1   g535(.A1(new_n344), .A2(new_n721), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n684), .A2(new_n649), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n652), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(new_n262), .ZN(G1332gat));
  NAND4_X1  g539(.A1(new_n684), .A2(new_n649), .A3(new_n594), .A4(new_n737), .ZN(new_n741));
  AND2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  OR3_X1    g541(.A1(new_n741), .A2(KEYINPUT111), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT111), .B1(new_n741), .B2(new_n742), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1333gat));
  NOR2_X1   g546(.A1(new_n738), .A2(G71gat), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n598), .B(KEYINPUT112), .Z(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G71gat), .B1(new_n738), .B2(new_n629), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1334gat));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n669), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g555(.A1(new_n721), .A2(new_n304), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT113), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n649), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT114), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n716), .A2(new_n761), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n762), .A2(new_n312), .A3(new_n652), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n684), .A2(new_n341), .A3(new_n758), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n684), .A2(KEYINPUT51), .A3(new_n341), .A4(new_n758), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(KEYINPUT115), .A3(new_n767), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n767), .A2(KEYINPUT115), .ZN(new_n769));
  INV_X1    g568(.A(new_n652), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .A4(new_n649), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n763), .B1(new_n312), .B2(new_n771), .ZN(G1336gat));
  NAND4_X1  g571(.A1(new_n708), .A2(new_n761), .A3(new_n594), .A4(new_n709), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(G92gat), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n656), .A2(G92gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n649), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n766), .B2(new_n767), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT52), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n768), .A2(new_n769), .A3(new_n649), .A4(new_n775), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT52), .B1(new_n773), .B2(G92gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(G1337gat));
  NOR2_X1   g581(.A1(new_n626), .A2(G99gat), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n769), .A3(new_n649), .A4(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G99gat), .B1(new_n762), .B2(new_n629), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(G1338gat));
  NOR3_X1   g585(.A1(new_n650), .A2(G106gat), .A3(new_n553), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n768), .A2(new_n769), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789));
  NOR4_X1   g588(.A1(new_n685), .A2(new_n760), .A3(new_n688), .A4(new_n553), .ZN(new_n790));
  INV_X1    g589(.A(G106gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n766), .A2(new_n767), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n708), .A2(new_n761), .A3(new_n603), .A4(new_n709), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n793), .A2(new_n787), .B1(new_n794), .B2(G106gat), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n788), .A2(new_n792), .B1(new_n795), .B2(new_n789), .ZN(G1339gat));
  NAND4_X1  g595(.A1(new_n342), .A2(new_n260), .A3(new_n650), .A4(new_n343), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n634), .A2(new_n643), .A3(new_n637), .A4(new_n638), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n641), .A2(KEYINPUT54), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n639), .A2(new_n802), .A3(new_n640), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n648), .A4(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n803), .A2(new_n648), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(new_n801), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT55), .B1(new_n807), .B2(new_n801), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n645), .A2(new_n648), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(new_n812), .A3(new_n721), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n244), .A2(new_n247), .A3(new_n254), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n236), .B1(new_n235), .B2(new_n238), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n240), .A2(new_n241), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n253), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n649), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n341), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n809), .A2(new_n812), .A3(new_n818), .A4(new_n341), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n305), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n799), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n652), .A2(new_n594), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n824), .A2(new_n598), .A3(new_n669), .A4(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(new_n466), .A3(new_n260), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n652), .B1(new_n799), .B2(new_n823), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(new_n582), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n656), .A3(new_n721), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n827), .B1(new_n830), .B2(new_n466), .ZN(G1340gat));
  OAI21_X1  g630(.A(G120gat), .B1(new_n826), .B2(new_n650), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n656), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n649), .A2(new_n468), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(G1341gat));
  OAI21_X1  g634(.A(G127gat), .B1(new_n826), .B2(new_n305), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n305), .A2(G127gat), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n833), .B2(new_n837), .ZN(G1342gat));
  NOR3_X1   g637(.A1(new_n833), .A2(G134gat), .A3(new_n687), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  OAI21_X1  g641(.A(G134gat), .B1(new_n826), .B2(new_n687), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(G1343gat));
  AOI21_X1  g643(.A(new_n553), .B1(new_n799), .B2(new_n823), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n825), .A2(new_n629), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n824), .B2(new_n603), .ZN(new_n849));
  OR3_X1    g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G141gat), .B1(new_n850), .B2(new_n260), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n629), .A2(KEYINPUT118), .A3(new_n595), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n828), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT118), .B1(new_n629), .B2(new_n595), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n854), .A2(new_n594), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n260), .A2(G141gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n851), .A2(new_n852), .A3(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n847), .A2(new_n849), .A3(new_n848), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n445), .B1(new_n860), .B2(new_n721), .ZN(new_n861));
  INV_X1    g660(.A(new_n858), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT58), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n859), .A2(new_n863), .ZN(G1344gat));
  NAND3_X1  g663(.A1(new_n856), .A2(new_n443), .A3(new_n649), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  INV_X1    g665(.A(new_n848), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n813), .A2(new_n819), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n687), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n304), .B1(new_n869), .B2(new_n821), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n797), .B(KEYINPUT116), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT57), .B(new_n595), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n845), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n823), .A2(new_n797), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n669), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n823), .A2(KEYINPUT120), .A3(new_n797), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n649), .B(new_n867), .C1(new_n876), .C2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n866), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  AOI211_X1 g682(.A(KEYINPUT59), .B(new_n443), .C1(new_n860), .C2(new_n649), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n865), .B1(new_n883), .B2(new_n884), .ZN(G1345gat));
  NAND2_X1  g684(.A1(new_n856), .A2(new_n304), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n451), .A2(new_n453), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n305), .A2(new_n887), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n886), .A2(new_n887), .B1(new_n860), .B2(new_n888), .ZN(G1346gat));
  OAI21_X1  g688(.A(KEYINPUT121), .B1(new_n850), .B2(new_n687), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n860), .A2(new_n891), .A3(new_n341), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(G162gat), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(G162gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n856), .A2(new_n894), .A3(new_n341), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1347gat));
  NAND2_X1  g695(.A1(new_n582), .A2(new_n594), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT122), .Z(new_n898));
  AOI211_X1 g697(.A(new_n770), .B(new_n898), .C1(new_n823), .C2(new_n799), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n390), .A3(new_n721), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n770), .A2(new_n656), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n824), .A2(new_n669), .A3(new_n749), .A4(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n260), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(G1348gat));
  NOR3_X1   g703(.A1(new_n902), .A2(new_n391), .A3(new_n650), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT124), .Z(new_n906));
  AOI21_X1  g705(.A(G176gat), .B1(new_n899), .B2(new_n649), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT123), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n906), .A2(new_n908), .ZN(G1349gat));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910));
  OR3_X1    g709(.A1(new_n902), .A2(new_n910), .A3(new_n305), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n902), .B2(new_n305), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(G183gat), .A3(new_n912), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n899), .B(new_n304), .C1(new_n386), .C2(new_n385), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT60), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n913), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1350gat));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n375), .A3(new_n341), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT126), .Z(new_n921));
  OAI21_X1  g720(.A(G190gat), .B1(new_n902), .B2(new_n687), .ZN(new_n922));
  XOR2_X1   g721(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n924), .ZN(G1351gat));
  NOR3_X1   g724(.A1(new_n770), .A2(new_n656), .A3(new_n665), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n845), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n350), .A3(new_n721), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n721), .B(new_n926), .C1(new_n876), .C2(new_n881), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n928), .B1(new_n930), .B2(new_n350), .ZN(G1352gat));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n351), .A3(new_n649), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT62), .Z(new_n933));
  OAI211_X1 g732(.A(new_n649), .B(new_n926), .C1(new_n876), .C2(new_n881), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n351), .B2(new_n935), .ZN(G1353gat));
  INV_X1    g735(.A(G211gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n927), .A2(new_n937), .A3(new_n304), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n304), .B(new_n926), .C1(new_n876), .C2(new_n881), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  INV_X1    g741(.A(G218gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n943), .A3(new_n341), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n341), .B(new_n926), .C1(new_n876), .C2(new_n881), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n946), .B2(new_n943), .ZN(G1355gat));
endmodule


