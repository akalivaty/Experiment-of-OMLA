//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT64), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT65), .B(G238), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n203), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G87), .A2(G250), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n211), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n202), .A2(new_n203), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n211), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(G250), .B1(G257), .B2(G264), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n227), .B1(new_n231), .B2(KEYINPUT0), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n220), .B(new_n232), .C1(KEYINPUT0), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G226), .B(G232), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  INV_X1    g0043(.A(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT67), .B(G107), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G58), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G222), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G77), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n255), .B1(new_n256), .B2(new_n253), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n224), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G274), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT68), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n265), .B2(new_n270), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(G226), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n262), .A2(G190), .A3(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT70), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n201), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n280), .A2(new_n224), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(G1), .B2(new_n225), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n225), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G150), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n283), .A2(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(G20), .B2(new_n204), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n279), .B1(new_n201), .B2(new_n282), .C1(new_n289), .C2(new_n281), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT9), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n262), .A2(new_n274), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n276), .B(new_n291), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n290), .B1(new_n294), .B2(G169), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n293), .A2(G179), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT71), .ZN(new_n302));
  INV_X1    g0102(.A(G232), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n257), .B2(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n253), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G97), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n253), .A2(G226), .A3(new_n254), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n304), .A2(new_n305), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n261), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT13), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n271), .B1(G238), .B2(new_n273), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n310), .B1(new_n309), .B2(new_n311), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT14), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(G179), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(G169), .C1(new_n312), .C2(new_n313), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n284), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n201), .B2(new_n287), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n280), .A2(new_n224), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(KEYINPUT11), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n282), .A2(new_n203), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT72), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(KEYINPUT11), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n278), .A2(new_n203), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT12), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n326), .A2(new_n328), .A3(new_n329), .A4(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(G200), .B1(new_n312), .B2(new_n313), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(new_n314), .B2(G190), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n320), .A2(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT76), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n253), .B2(G20), .ZN(new_n339));
  INV_X1    g0139(.A(G33), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT3), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT3), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G68), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n286), .A2(G159), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G58), .A2(G68), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT73), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(KEYINPUT73), .A2(G58), .A3(G68), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n221), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT74), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT74), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n356), .A3(G20), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n347), .A2(new_n348), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT16), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n355), .A2(new_n357), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n361), .A2(KEYINPUT16), .A3(new_n347), .A4(new_n348), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n324), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n283), .A2(new_n278), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n282), .B2(new_n283), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n253), .A2(G226), .A3(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G87), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n253), .A2(new_n254), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n368), .B(new_n369), .C1(new_n370), .C2(new_n258), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n261), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n271), .B1(G232), .B2(new_n273), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT75), .B1(new_n374), .B2(G179), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  INV_X1    g0176(.A(G179), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n372), .A2(new_n373), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n315), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n375), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT18), .B1(new_n367), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G190), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n374), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n292), .B1(new_n372), .B2(new_n373), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(new_n363), .A3(new_n366), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT17), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n281), .B1(new_n358), .B2(new_n359), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n365), .B1(new_n388), .B2(new_n362), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT17), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n390), .A3(new_n385), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n337), .A2(new_n381), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n367), .A2(new_n380), .A3(KEYINPUT18), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT18), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n375), .A2(new_n378), .A3(new_n379), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n394), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n393), .A2(new_n396), .A3(KEYINPUT76), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n283), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n286), .B1(G20), .B2(G77), .ZN(new_n400));
  XOR2_X1   g0200(.A(KEYINPUT15), .B(G87), .Z(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n400), .B1(new_n284), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n324), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n282), .A2(new_n256), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n404), .B(new_n405), .C1(G77), .C2(new_n277), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n273), .A2(G244), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n344), .A2(G107), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n408), .B1(new_n257), .B2(new_n212), .C1(new_n303), .C2(new_n370), .ZN(new_n409));
  AOI211_X1 g0209(.A(new_n271), .B(new_n407), .C1(new_n409), .C2(new_n261), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n406), .B1(new_n410), .B2(G169), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT69), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n406), .B(KEYINPUT69), .C1(new_n410), .C2(G169), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(new_n377), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n410), .A2(G190), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n405), .B1(G77), .B2(new_n277), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n403), .B2(new_n324), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n417), .B(new_n419), .C1(new_n292), .C2(new_n410), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  NOR4_X1   g0221(.A1(new_n301), .A2(new_n336), .A3(new_n398), .A4(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT5), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n263), .B(G45), .C1(new_n423), .C2(G41), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT68), .B(G41), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n423), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G274), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n253), .A2(G250), .A3(new_n254), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n253), .A2(G257), .A3(G1698), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G294), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n261), .ZN(new_n432));
  INV_X1    g0232(.A(new_n424), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n266), .A2(new_n268), .A3(new_n423), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n261), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT85), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n435), .A2(new_n436), .A3(G264), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n436), .B1(new_n435), .B2(G264), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n427), .B(new_n432), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G200), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n260), .A2(new_n224), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n266), .A2(new_n268), .A3(new_n423), .ZN(new_n442));
  OAI211_X1 g0242(.A(G264), .B(new_n441), .C1(new_n442), .C2(new_n424), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT85), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n435), .A2(new_n436), .A3(G264), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n446), .A2(G190), .A3(new_n427), .A4(new_n432), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT84), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n341), .A2(new_n343), .A3(new_n225), .A4(G87), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT83), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT83), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n253), .A2(new_n452), .A3(new_n225), .A4(G87), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n453), .A3(KEYINPUT22), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n225), .A2(KEYINPUT23), .A3(G107), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT23), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(G20), .B2(new_n207), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n455), .B(new_n457), .C1(G116), .C2(new_n321), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT22), .B1(new_n451), .B2(new_n453), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n449), .B(KEYINPUT24), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n451), .A2(new_n453), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT22), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(new_n454), .A4(new_n458), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n454), .A3(new_n458), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n449), .B1(new_n468), .B2(KEYINPUT24), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n324), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n278), .A2(new_n207), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n471), .A2(KEYINPUT25), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(KEYINPUT25), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n281), .B(new_n277), .C1(G1), .C2(new_n340), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n472), .B(new_n473), .C1(new_n207), .C2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n448), .A2(new_n470), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n446), .A2(G179), .A3(new_n427), .A4(new_n432), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(KEYINPUT86), .B1(new_n439), .B2(G169), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n444), .A2(new_n445), .B1(new_n261), .B2(new_n431), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT86), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(G179), .A4(new_n427), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n470), .A2(new_n476), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n341), .A2(new_n343), .A3(G244), .A4(new_n254), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(KEYINPUT77), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n253), .A2(G244), .A3(new_n254), .A4(new_n487), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n486), .A2(KEYINPUT77), .B1(G33), .B2(G283), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n261), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n435), .A2(G257), .B1(new_n426), .B2(G274), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n377), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT79), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT79), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n494), .A2(new_n498), .A3(new_n377), .A4(new_n495), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n500), .A2(new_n206), .A3(G107), .ZN(new_n501));
  XNOR2_X1  g0301(.A(G97), .B(G107), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n503), .A2(new_n225), .B1(new_n256), .B2(new_n287), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n207), .B1(new_n339), .B2(new_n345), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n324), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n277), .A2(G97), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n340), .A2(G1), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n278), .A2(new_n324), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n507), .B1(new_n509), .B2(G97), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n497), .A2(new_n499), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n494), .A2(new_n495), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT78), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT78), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n494), .A2(new_n516), .A3(new_n495), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n315), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n517), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G190), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n511), .B1(G200), .B2(new_n514), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n513), .A2(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n435), .A2(G270), .B1(new_n426), .B2(G274), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n341), .A2(new_n343), .A3(G257), .A4(new_n254), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n341), .A2(new_n343), .A3(G264), .A4(G1698), .ZN(new_n525));
  INV_X1    g0325(.A(G303), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n524), .B(new_n525), .C1(new_n526), .C2(new_n253), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n261), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n315), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT21), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n523), .A2(G179), .A3(new_n528), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n277), .A2(G116), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n509), .B2(G116), .ZN(new_n534));
  AOI21_X1  g0334(.A(G20), .B1(G33), .B2(G283), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n340), .A2(G97), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT81), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT81), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n280), .A2(new_n224), .B1(G20), .B2(new_n244), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT20), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT81), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT81), .B1(new_n535), .B2(new_n536), .ZN(new_n545));
  OAI211_X1 g0345(.A(KEYINPUT20), .B(new_n542), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n534), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n532), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n527), .A2(new_n261), .ZN(new_n550));
  OAI211_X1 g0350(.A(G270), .B(new_n441), .C1(new_n442), .C2(new_n424), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n427), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G190), .ZN(new_n554));
  INV_X1    g0354(.A(new_n533), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n474), .B2(new_n244), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT20), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n556), .B1(new_n559), .B2(new_n546), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n554), .B(new_n560), .C1(new_n292), .C2(new_n553), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n529), .A2(new_n548), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT21), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT82), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT82), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n565), .B(KEYINPUT21), .C1(new_n529), .C2(new_n548), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n549), .B(new_n561), .C1(new_n564), .C2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n253), .A2(new_n225), .A3(G68), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT19), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n225), .B1(new_n306), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(G87), .B2(new_n208), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n284), .B2(new_n206), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n324), .B1(new_n278), .B2(new_n402), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n509), .A2(G87), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n263), .A2(G45), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n577), .B(G250), .C1(new_n260), .C2(new_n224), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n263), .A2(G45), .A3(G274), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT80), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT80), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n581), .A2(new_n263), .A3(G45), .A4(G274), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n341), .A2(new_n343), .A3(G244), .A4(G1698), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n341), .A2(new_n343), .A3(G238), .A4(new_n254), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(new_n585), .C1(new_n340), .C2(new_n244), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n583), .B1(new_n586), .B2(new_n261), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G190), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n576), .B(new_n588), .C1(new_n292), .C2(new_n587), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n574), .B1(new_n402), .B2(new_n474), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n586), .A2(new_n261), .ZN(new_n591));
  INV_X1    g0391(.A(new_n583), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n377), .A3(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n590), .B(new_n593), .C1(G169), .C2(new_n587), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n567), .A2(new_n595), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n422), .A2(new_n484), .A3(new_n522), .A4(new_n596), .ZN(G372));
  NAND2_X1  g0397(.A1(new_n320), .A2(new_n332), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n416), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n334), .A2(new_n333), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n390), .B1(new_n389), .B2(new_n385), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n389), .A2(new_n390), .A3(new_n385), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n389), .A2(new_n395), .A3(new_n394), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n601), .A2(new_n605), .B1(new_n381), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n299), .B1(new_n607), .B2(new_n296), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n301), .A2(new_n398), .A3(new_n421), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n335), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n580), .A2(new_n582), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT87), .B1(new_n611), .B2(new_n578), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n578), .A2(KEYINPUT87), .A3(new_n580), .A4(new_n582), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n591), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n315), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT88), .B1(new_n616), .B2(new_n593), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT87), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n583), .A2(new_n618), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n619), .A2(new_n613), .B1(new_n586), .B2(new_n261), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n593), .B(KEYINPUT88), .C1(new_n620), .C2(G169), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n590), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n494), .A2(new_n516), .A3(new_n495), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n516), .B1(new_n494), .B2(new_n495), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n625), .A2(new_n626), .A3(G169), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(new_n512), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n589), .A2(new_n594), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n624), .B1(new_n630), .B2(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n588), .A2(new_n575), .A3(new_n574), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n620), .A2(new_n292), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n628), .A2(new_n632), .A3(new_n623), .A4(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n448), .A2(new_n470), .A3(new_n476), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT88), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n619), .A2(new_n613), .ZN(new_n640));
  AOI21_X1  g0440(.A(G169), .B1(new_n640), .B2(new_n591), .ZN(new_n641));
  AOI211_X1 g0441(.A(G179), .B(new_n583), .C1(new_n586), .C2(new_n261), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n621), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n635), .B1(new_n644), .B2(new_n590), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n549), .B1(new_n564), .B2(new_n566), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n638), .B(new_n645), .C1(new_n483), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n520), .A2(new_n521), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n518), .A2(new_n499), .A3(new_n511), .A4(new_n497), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n631), .B(new_n637), .C1(new_n647), .C2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n608), .B1(new_n610), .B2(new_n652), .ZN(G369));
  AND2_X1   g0453(.A1(new_n225), .A2(G13), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n263), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n560), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n567), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n646), .A2(new_n662), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT89), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT89), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n470), .A2(new_n476), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n479), .A2(new_n482), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n638), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT24), .B1(new_n459), .B2(new_n460), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT84), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(new_n466), .A3(new_n461), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n475), .B1(new_n677), .B2(new_n324), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n661), .ZN(new_n679));
  OAI22_X1  g0479(.A1(new_n674), .A2(new_n679), .B1(new_n673), .B2(new_n661), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n670), .A2(G330), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n646), .A2(new_n661), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n484), .A2(new_n683), .B1(new_n483), .B2(new_n661), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n684), .ZN(G399));
  NOR2_X1   g0485(.A1(new_n229), .A2(new_n425), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n222), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n638), .A2(new_n645), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n560), .B1(new_n530), .B2(new_n531), .ZN(new_n693));
  OAI21_X1  g0493(.A(G169), .B1(new_n550), .B2(new_n552), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n563), .B1(new_n694), .B2(new_n560), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n565), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n562), .A2(KEYINPUT82), .A3(new_n563), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n693), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n439), .A2(G169), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n699), .A2(new_n482), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n698), .B1(new_n678), .B2(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT93), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT93), .B1(new_n648), .B2(new_n649), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n692), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n628), .A2(new_n629), .A3(new_n632), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n623), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n632), .B1(new_n645), .B2(new_n628), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n660), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT94), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n651), .A2(new_n661), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT94), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI211_X1 g0515(.A(new_n714), .B(new_n660), .C1(new_n705), .C2(new_n709), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n712), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G330), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n484), .A2(new_n596), .A3(new_n522), .A4(new_n661), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT31), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT90), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n625), .A2(new_n626), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n480), .A2(new_n553), .A3(G179), .A4(new_n587), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n432), .B1(new_n437), .B2(new_n438), .ZN(new_n726));
  INV_X1    g0526(.A(new_n587), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n726), .A2(new_n531), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n519), .A2(new_n728), .A3(KEYINPUT90), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n724), .A2(new_n725), .A3(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n553), .A2(G179), .A3(new_n620), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n439), .A3(new_n514), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n730), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n661), .B1(new_n735), .B2(KEYINPUT92), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT92), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n730), .A2(new_n737), .A3(new_n732), .A4(new_n734), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n720), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n660), .A2(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n730), .A2(new_n734), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT91), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n731), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n730), .A2(KEYINPUT91), .A3(new_n734), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n718), .B1(new_n740), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n717), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n691), .B1(new_n750), .B2(G1), .ZN(G364));
  NAND3_X1  g0551(.A1(new_n667), .A2(G330), .A3(new_n669), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n263), .B1(new_n654), .B2(G45), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n687), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G330), .B2(new_n670), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n224), .B1(G20), .B2(new_n315), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n225), .A2(new_n382), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n377), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n225), .A2(G190), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n292), .A2(G179), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n761), .A2(new_n202), .B1(new_n764), .B2(new_n207), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G179), .A2(G200), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n225), .B1(new_n766), .B2(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n762), .A2(new_n760), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n253), .B1(new_n767), .B2(new_n206), .C1(new_n256), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n759), .A2(new_n763), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n765), .B(new_n769), .C1(G87), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n762), .A2(new_n766), .ZN(new_n773));
  INV_X1    g0573(.A(G159), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT32), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n225), .A2(new_n377), .A3(new_n292), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n779), .A2(new_n382), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n779), .A2(G190), .A3(new_n780), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n777), .B1(new_n203), .B2(new_n781), .C1(new_n201), .C2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G311), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n344), .B1(new_n768), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n761), .ZN(new_n790));
  INV_X1    g0590(.A(new_n764), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G322), .A2(new_n790), .B1(new_n791), .B2(G283), .ZN(new_n792));
  INV_X1    g0592(.A(new_n773), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G303), .A2(new_n771), .B1(new_n793), .B2(G329), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n767), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n789), .B(new_n795), .C1(G294), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT100), .B(G317), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT33), .ZN(new_n799));
  INV_X1    g0599(.A(G326), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n797), .B1(new_n781), .B2(new_n799), .C1(new_n800), .C2(new_n786), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n758), .B1(new_n787), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n757), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n251), .A2(G45), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n229), .A2(new_n253), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n270), .B2(new_n223), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n229), .A2(new_n344), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(G355), .B(KEYINPUT95), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n813), .A2(new_n814), .B1(G116), .B2(new_n228), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT96), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n808), .A2(new_n811), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n807), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n802), .A2(new_n819), .A3(new_n754), .ZN(new_n820));
  INV_X1    g0620(.A(new_n805), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n668), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n756), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  INV_X1    g0624(.A(new_n754), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n758), .A2(new_n804), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(G77), .B2(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n344), .B1(new_n767), .B2(new_n206), .C1(new_n244), .C2(new_n768), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G107), .A2(new_n771), .B1(new_n793), .B2(G311), .ZN(new_n829));
  INV_X1    g0629(.A(G87), .ZN(new_n830));
  INV_X1    g0630(.A(G294), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n830), .B2(new_n764), .C1(new_n831), .C2(new_n761), .ZN(new_n832));
  INV_X1    g0632(.A(new_n781), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n828), .B(new_n832), .C1(G283), .C2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n526), .B2(new_n786), .ZN(new_n835));
  INV_X1    g0635(.A(new_n768), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G143), .A2(new_n790), .B1(new_n836), .B2(G159), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n781), .B2(new_n285), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n785), .B2(G137), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT34), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G68), .A2(new_n791), .B1(new_n793), .B2(G132), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n344), .B1(new_n771), .B2(G50), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(new_n202), .C2(new_n767), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n835), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n827), .B1(new_n844), .B2(new_n757), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n419), .A2(new_n661), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n600), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n846), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n416), .A2(new_n420), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n845), .B1(new_n850), .B2(new_n804), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT26), .B1(new_n649), .B2(new_n595), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n637), .A2(new_n623), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n702), .A2(new_n638), .A3(new_n522), .A4(new_n645), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n660), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT102), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(new_n850), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n483), .A2(new_n646), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n638), .A2(new_n645), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n858), .A2(new_n859), .A3(new_n650), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n637), .A2(new_n852), .A3(new_n623), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n850), .B(new_n661), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT102), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n850), .B(KEYINPUT101), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n857), .A2(new_n863), .B1(new_n864), .B2(new_n713), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n825), .B1(new_n865), .B2(new_n748), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n866), .A2(KEYINPUT103), .B1(new_n748), .B2(new_n865), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n866), .A2(KEYINPUT103), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n851), .B1(new_n867), .B2(new_n868), .ZN(G384));
  XNOR2_X1  g0669(.A(new_n503), .B(KEYINPUT104), .ZN(new_n870));
  OAI211_X1 g0670(.A(G116), .B(new_n226), .C1(new_n870), .C2(KEYINPUT35), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(KEYINPUT35), .B2(new_n870), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT36), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n223), .A2(G77), .A3(new_n351), .A4(new_n352), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(KEYINPUT105), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n874), .A2(KEYINPUT105), .B1(new_n201), .B2(G68), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n263), .B(G13), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n735), .A2(KEYINPUT92), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n879), .A2(KEYINPUT31), .A3(new_n660), .A4(new_n738), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT108), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT108), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n736), .A2(new_n882), .A3(KEYINPUT31), .A4(new_n738), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n740), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n381), .A2(new_n606), .B1(new_n604), .B2(new_n603), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n389), .A2(new_n658), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n889));
  OAI21_X1  g0689(.A(new_n386), .B1(new_n389), .B2(new_n395), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n889), .B1(new_n890), .B2(new_n887), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n367), .A2(new_n380), .ZN(new_n892));
  INV_X1    g0692(.A(new_n658), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n367), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n889), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n892), .A2(new_n894), .A3(new_n386), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n888), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n393), .A2(new_n396), .A3(KEYINPUT76), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n604), .A2(new_n603), .B1(new_n396), .B2(KEYINPUT76), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n887), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n890), .B2(new_n887), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n896), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n332), .A2(new_n660), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n598), .A2(new_n602), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n598), .A2(new_n661), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n850), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n885), .A2(new_n906), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n884), .B2(new_n740), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n894), .B1(new_n392), .B2(new_n397), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n903), .A2(new_n896), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT40), .B1(new_n917), .B2(new_n905), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n912), .A2(KEYINPUT40), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n881), .A2(new_n883), .B1(new_n720), .B2(new_n739), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n919), .A2(new_n610), .A3(new_n920), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n920), .A2(new_n610), .A3(new_n718), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n885), .A2(new_n911), .A3(new_n918), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n398), .A2(new_n887), .B1(new_n903), .B2(new_n896), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n898), .B1(new_n924), .B2(KEYINPUT38), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n920), .A2(new_n925), .A3(new_n910), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT40), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n922), .B1(new_n928), .B2(G330), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n921), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n422), .B(new_n712), .C1(new_n715), .C2(new_n716), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n608), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n599), .A2(new_n661), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n936), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT39), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n917), .B2(new_n905), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n935), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n393), .A2(new_n396), .A3(new_n658), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n416), .A2(new_n660), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n863), .B2(new_n857), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT38), .B1(new_n902), .B2(new_n904), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n936), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n908), .A2(new_n909), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT107), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n933), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n263), .B2(new_n654), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n933), .A2(new_n950), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n878), .B1(new_n952), .B2(new_n953), .ZN(G367));
  NAND2_X1  g0754(.A1(new_n511), .A2(new_n660), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n703), .B2(new_n704), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n628), .A2(new_n660), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(new_n484), .A3(new_n683), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(KEYINPUT42), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n649), .B1(new_n956), .B2(new_n673), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n959), .A2(KEYINPUT42), .B1(new_n661), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n576), .A2(new_n661), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n623), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(new_n645), .B2(new_n964), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n960), .A2(new_n962), .B1(KEYINPUT43), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n968), .B(new_n969), .Z(new_n970));
  INV_X1    g0770(.A(new_n958), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n681), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n970), .B(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n686), .B(KEYINPUT41), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  MUX2_X1   g0775(.A(new_n674), .B(new_n680), .S(new_n682), .Z(new_n976));
  XNOR2_X1  g0776(.A(new_n752), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n750), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT111), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n750), .A2(new_n977), .A3(KEYINPUT111), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n958), .A2(new_n684), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n985));
  OR3_X1    g0785(.A1(new_n958), .A2(new_n684), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n985), .B1(new_n958), .B2(new_n684), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AND3_X1   g0789(.A1(new_n984), .A2(new_n681), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n681), .B1(new_n989), .B2(new_n984), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT110), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(KEYINPUT110), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n980), .A2(new_n981), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n975), .B1(new_n994), .B2(new_n750), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n753), .B(KEYINPUT112), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n973), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n807), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n228), .B2(new_n402), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n810), .A2(new_n241), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n825), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n253), .B1(new_n767), .B2(new_n203), .C1(new_n201), .C2(new_n768), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G77), .A2(new_n791), .B1(new_n793), .B2(G137), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n202), .B2(new_n770), .C1(new_n285), .C2(new_n761), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1002), .B(new_n1004), .C1(G159), .C2(new_n833), .ZN(new_n1005));
  INV_X1    g0805(.A(G143), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n1006), .B2(new_n786), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n785), .A2(G311), .B1(G303), .B2(new_n790), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1008), .A2(KEYINPUT113), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n771), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT46), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n770), .B2(new_n244), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(new_n207), .C2(new_n767), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G283), .A2(new_n836), .B1(new_n793), .B2(G317), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n344), .C1(new_n206), .C2(new_n764), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(G294), .C2(new_n833), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n1008), .B2(KEYINPUT113), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1007), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT47), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n758), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1001), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n821), .B2(new_n967), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n997), .A2(new_n1023), .ZN(G387));
  INV_X1    g0824(.A(new_n981), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT111), .B1(new_n750), .B2(new_n977), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n686), .B1(new_n750), .B2(new_n977), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n680), .A2(new_n821), .ZN(new_n1028));
  OAI21_X1  g0828(.A(KEYINPUT50), .B1(new_n283), .B2(G50), .ZN(new_n1029));
  AOI21_X1  g0829(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n688), .A3(new_n1030), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n283), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n809), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n238), .A2(new_n270), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n688), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n812), .A2(new_n1035), .B1(new_n207), .B2(new_n229), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1033), .A2(new_n1034), .B1(KEYINPUT114), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(KEYINPUT114), .B2(new_n1036), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n825), .B1(new_n1038), .B2(new_n807), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n770), .A2(new_n256), .B1(new_n768), .B2(new_n203), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n761), .A2(new_n201), .B1(new_n773), .B2(new_n285), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n253), .B1(new_n764), .B2(new_n206), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n402), .A2(new_n767), .ZN(new_n1043));
  NOR4_X1   g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n283), .B2(new_n781), .C1(new_n786), .C2(new_n774), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n253), .B1(new_n791), .B2(G116), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G317), .A2(new_n790), .B1(new_n836), .B2(G303), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n781), .B2(new_n788), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n785), .B2(G322), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT48), .ZN(new_n1050));
  INV_X1    g0850(.A(G283), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n770), .A2(new_n831), .B1(new_n767), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1046), .B1(new_n800), .B2(new_n773), .C1(new_n1053), .C2(KEYINPUT49), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1053), .A2(KEYINPUT49), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1045), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1039), .B1(new_n1056), .B2(new_n757), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n977), .A2(new_n996), .B1(new_n1028), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1027), .A2(new_n1058), .ZN(G393));
  OR2_X1    g0859(.A1(new_n990), .A2(new_n991), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(new_n994), .A3(new_n686), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n996), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n785), .A2(G317), .B1(G311), .B2(new_n790), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1066));
  XNOR2_X1  g0866(.A(new_n1065), .B(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n781), .A2(new_n526), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G294), .A2(new_n836), .B1(new_n793), .B2(G322), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1051), .B2(new_n770), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n344), .B1(new_n767), .B2(new_n244), .C1(new_n207), .C2(new_n764), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n785), .A2(G150), .B1(G159), .B2(new_n790), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n781), .A2(new_n201), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G68), .A2(new_n771), .B1(new_n793), .B2(G143), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n283), .B2(new_n768), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n253), .B1(new_n767), .B2(new_n256), .C1(new_n830), .C2(new_n764), .ZN(new_n1078));
  NOR4_X1   g0878(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n757), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n807), .B1(G97), .B2(new_n229), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n247), .A2(new_n809), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n754), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1080), .B(new_n1083), .C1(new_n958), .C2(new_n821), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1062), .A2(new_n1064), .A3(new_n1084), .ZN(G390));
  NAND3_X1  g0885(.A1(new_n885), .A2(G330), .A3(new_n911), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n934), .B1(new_n944), .B2(new_n947), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n937), .A2(new_n939), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n705), .A2(new_n709), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n661), .A3(new_n850), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n943), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n947), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n934), .B1(new_n936), .B2(new_n898), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1086), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(KEYINPUT31), .A2(new_n719), .B1(new_n736), .B2(new_n738), .ZN(new_n1098));
  OAI211_X1 g0898(.A(G330), .B(new_n850), .C1(new_n1098), .C2(new_n746), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(new_n947), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1100), .B(new_n1095), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n885), .A2(G330), .A3(new_n422), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n608), .A3(new_n931), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n943), .B1(new_n710), .B2(new_n850), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n947), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n748), .A2(new_n850), .A3(new_n1106), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n920), .A2(new_n718), .A3(new_n864), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1105), .B(new_n1107), .C1(new_n1108), .C2(new_n1106), .ZN(new_n1109));
  AND4_X1   g0909(.A1(new_n856), .A2(new_n651), .A3(new_n661), .A4(new_n850), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n856), .B1(new_n855), .B2(new_n850), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1092), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n920), .A2(new_n718), .A3(new_n910), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1106), .B1(new_n748), .B2(new_n850), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1104), .B1(new_n1109), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n687), .B1(new_n1102), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n932), .A2(new_n922), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1105), .B1(new_n1099), .B2(new_n947), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n864), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n885), .A2(G330), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1119), .B1(new_n947), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1099), .A2(new_n947), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n944), .B1(new_n1086), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1118), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT116), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1125), .B(KEYINPUT116), .C1(new_n1097), .C2(new_n1101), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1117), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n344), .B1(new_n793), .B2(G125), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n201), .B2(new_n764), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT118), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n833), .A2(G137), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n770), .A2(new_n285), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n796), .A2(G159), .ZN(new_n1137));
  XOR2_X1   g0937(.A(KEYINPUT54), .B(G143), .Z(new_n1138));
  AOI22_X1  g0938(.A1(G132), .A2(new_n790), .B1(new_n836), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1133), .B(new_n1140), .C1(G128), .C2(new_n785), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n344), .B1(new_n767), .B2(new_n256), .C1(new_n830), .C2(new_n770), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n761), .A2(new_n244), .B1(new_n764), .B2(new_n203), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n768), .A2(new_n206), .B1(new_n773), .B2(new_n831), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n207), .B2(new_n781), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G283), .B2(new_n785), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n757), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1148), .B(new_n825), .C1(new_n399), .C2(new_n826), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n1088), .B2(new_n803), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n935), .B1(new_n1112), .B2(new_n1106), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n937), .A2(new_n939), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1096), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1113), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1089), .A2(new_n1107), .A3(new_n1096), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n996), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT117), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1154), .A2(KEYINPUT117), .A3(new_n996), .A4(new_n1155), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1150), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1130), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(G378));
  INV_X1    g0962(.A(KEYINPUT57), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1116), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n1118), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n949), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n290), .A2(new_n893), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n301), .B(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n927), .B1(new_n913), .B2(new_n906), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n927), .B1(new_n936), .B2(new_n945), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1172), .A2(new_n920), .A3(new_n910), .ZN(new_n1173));
  OAI211_X1 g0973(.A(G330), .B(new_n1170), .C1(new_n1171), .C2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1170), .B1(new_n928), .B2(G330), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1166), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1170), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n919), .B2(new_n718), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n949), .A3(new_n1174), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n687), .B1(new_n1165), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT121), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n949), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1179), .A2(new_n1174), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1185), .A2(KEYINPUT121), .A3(new_n1166), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1184), .A2(new_n1186), .B1(new_n1118), .B2(new_n1164), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1182), .B1(new_n1187), .B2(KEYINPUT57), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1178), .A2(new_n803), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n825), .B1(G50), .B2(new_n826), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n253), .A2(new_n425), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G50), .B(new_n1191), .C1(new_n340), .C2(new_n265), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1191), .B1(new_n203), .B2(new_n767), .C1(new_n256), .C2(new_n770), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n402), .A2(new_n768), .B1(new_n207), .B2(new_n761), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n764), .A2(new_n202), .B1(new_n773), .B2(new_n1051), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n206), .B2(new_n781), .C1(new_n786), .C2(new_n244), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1192), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(G132), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n781), .A2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G128), .A2(new_n790), .B1(new_n836), .B2(G137), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1138), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1202), .B1(new_n285), .B2(new_n767), .C1(new_n770), .C2(new_n1203), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1201), .B(new_n1204), .C1(new_n785), .C2(G125), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n774), .B2(new_n764), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT119), .Z(new_n1210));
  INV_X1    g1010(.A(KEYINPUT59), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1210), .B1(new_n1205), .B2(new_n1211), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1199), .B1(new_n1198), .B2(new_n1197), .C1(new_n1207), .C2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1190), .B1(new_n1213), .B2(new_n757), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1189), .A2(KEYINPUT120), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT120), .B1(new_n1189), .B2(new_n1214), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1218), .B2(new_n996), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1188), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n947), .A2(new_n803), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n825), .B1(G68), .B2(new_n826), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n253), .B1(new_n764), .B2(new_n202), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G137), .A2(new_n790), .B1(new_n793), .B2(G128), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n285), .B2(new_n768), .C1(new_n774), .C2(new_n770), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G50), .C2(new_n796), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n1200), .B2(new_n786), .C1(new_n781), .C2(new_n1203), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n344), .B1(new_n764), .B2(new_n256), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT122), .Z(new_n1230));
  OAI22_X1  g1030(.A1(new_n768), .A2(new_n207), .B1(new_n773), .B2(new_n526), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n206), .A2(new_n770), .B1(new_n761), .B2(new_n1051), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1230), .A2(new_n1043), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n244), .B2(new_n781), .C1(new_n786), .C2(new_n831), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1228), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1223), .B1(new_n1235), .B2(new_n757), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT123), .Z(new_n1237));
  AOI22_X1  g1037(.A1(new_n1221), .A2(new_n996), .B1(new_n1222), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1125), .A2(new_n974), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1221), .A2(new_n1118), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(G381));
  NAND3_X1  g1041(.A1(new_n1027), .A2(new_n823), .A3(new_n1058), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1242), .A2(G384), .ZN(new_n1243));
  AOI211_X1 g1043(.A(G381), .B(G390), .C1(new_n1243), .C2(KEYINPUT124), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(KEYINPUT124), .B2(new_n1243), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1188), .A2(new_n1161), .A3(new_n1219), .ZN(new_n1246));
  OR3_X1    g1046(.A1(new_n1245), .A2(G387), .A3(new_n1246), .ZN(G407));
  NAND2_X1  g1047(.A1(new_n659), .A2(G213), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT125), .Z(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(new_n1246), .C2(new_n1250), .ZN(G409));
  INV_X1    g1051(.A(KEYINPUT127), .ZN(new_n1252));
  INV_X1    g1052(.A(G390), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(G387), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1242), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n823), .B1(new_n1027), .B2(new_n1058), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n997), .A2(new_n1023), .A3(G390), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G390), .B1(new_n997), .B2(new_n1023), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1254), .A2(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1261), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1263), .A2(new_n1257), .A3(new_n1252), .A4(new_n1259), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT126), .B1(new_n1221), .B2(new_n1118), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(KEYINPUT60), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  OAI211_X1 g1069(.A(KEYINPUT126), .B(new_n1269), .C1(new_n1221), .C2(new_n1118), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1268), .A2(new_n686), .A3(new_n1125), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1238), .ZN(new_n1272));
  INV_X1    g1072(.A(G384), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1271), .A2(G384), .A3(new_n1238), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1249), .A2(G2897), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1276), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1275), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1271), .B2(new_n1238), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1161), .B1(new_n1188), .B2(new_n1219), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1164), .A2(new_n1118), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1166), .B1(new_n1185), .B2(KEYINPUT121), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT121), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1285), .B(new_n949), .C1(new_n1179), .C2(new_n1174), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n974), .B(new_n1283), .C1(new_n1284), .C2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1217), .B1(new_n1181), .B2(new_n996), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1287), .A2(new_n1288), .A3(new_n1130), .A4(new_n1160), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1250), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1277), .B(new_n1281), .C1(new_n1282), .C2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1282), .A2(new_n1290), .A3(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1291), .B(new_n1292), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G375), .A2(G378), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1290), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1293), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1300), .A2(KEYINPUT62), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1266), .B1(new_n1296), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1281), .A2(new_n1277), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT61), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT63), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1300), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1294), .A2(KEYINPUT63), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1305), .A2(new_n1307), .A3(new_n1265), .A4(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1302), .A2(new_n1309), .ZN(G405));
  NAND2_X1  g1110(.A1(new_n1297), .A2(new_n1246), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1299), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1297), .A2(new_n1246), .A3(new_n1293), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1265), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1265), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(G402));
endmodule


