//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT24), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(G183gat), .A3(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G183gat), .B2(G190gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n213), .B(new_n220), .C1(new_n211), .C2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n209), .A2(new_n210), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n223), .A2(KEYINPUT26), .A3(new_n205), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n205), .A2(KEYINPUT26), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(new_n214), .B2(new_n215), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT65), .B(G190gat), .Z(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT27), .B(G183gat), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n228), .A2(KEYINPUT28), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT28), .B1(new_n228), .B2(new_n229), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n227), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n228), .A2(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT25), .B1(new_n233), .B2(new_n211), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n222), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT66), .B(G134gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G127gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT67), .B(G127gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G134gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n240));
  XOR2_X1   g039(.A(G113gat), .B(G120gat), .Z(new_n241));
  AOI22_X1  g040(.A1(new_n237), .A2(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n235), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n237), .A2(new_n239), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n241), .A2(new_n240), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n251), .A2(new_n222), .A3(new_n232), .A4(new_n234), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n247), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n204), .B1(new_n253), .B2(KEYINPUT32), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT33), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n253), .A2(KEYINPUT68), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT68), .B1(new_n253), .B2(new_n255), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n254), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n253), .B(KEYINPUT32), .C1(new_n255), .C2(new_n204), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n248), .B1(new_n247), .B2(new_n252), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT34), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n262), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G141gat), .ZN(new_n267));
  INV_X1    g066(.A(G148gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT76), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT76), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n273), .A3(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275));
  INV_X1    g074(.A(G155gat), .ZN(new_n276));
  INV_X1    g075(.A(G162gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n275), .B1(new_n278), .B2(KEYINPUT2), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n272), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n269), .A2(new_n282), .A3(new_n270), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n278), .A2(KEYINPUT75), .ZN(new_n284));
  OR3_X1    g083(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .A4(new_n275), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT29), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT83), .ZN(new_n291));
  OR2_X1    g090(.A1(G197gat), .A2(G204gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(G197gat), .A2(G204gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT22), .ZN(new_n294));
  NAND2_X1  g093(.A1(G211gat), .A2(G218gat), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n292), .A2(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(G211gat), .A2(G218gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n295), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n299), .B1(new_n298), .B2(new_n295), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n297), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n302), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(new_n296), .A3(new_n300), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n303), .A2(KEYINPUT71), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT71), .B1(new_n303), .B2(new_n305), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT83), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n289), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n291), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n303), .A2(new_n288), .A3(new_n305), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n280), .A2(new_n286), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n281), .B1(new_n280), .B2(new_n286), .ZN(new_n315));
  INV_X1    g114(.A(G228gat), .ZN(new_n316));
  INV_X1    g115(.A(G233gat), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n311), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT3), .B1(new_n312), .B2(KEYINPUT82), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n303), .A2(new_n305), .A3(new_n321), .A4(new_n288), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n313), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n305), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n290), .A2(new_n325), .ZN(new_n326));
  OAI22_X1  g125(.A1(new_n323), .A2(new_n326), .B1(new_n316), .B2(new_n317), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(KEYINPUT31), .B(G50gat), .Z(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G78gat), .B(G106gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(G22gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n329), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n319), .A2(new_n327), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n330), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n332), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n319), .A2(new_n327), .A3(new_n333), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n333), .B1(new_n319), .B2(new_n327), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n258), .A2(new_n263), .A3(new_n264), .A4(new_n259), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n266), .A2(new_n335), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT87), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n339), .A2(new_n335), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n344), .A2(KEYINPUT87), .A3(new_n266), .A4(new_n340), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n280), .A2(new_n286), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n251), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n246), .A2(new_n313), .A3(KEYINPUT78), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n313), .B2(new_n281), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n315), .A2(KEYINPUT77), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n251), .A4(new_n287), .ZN(new_n356));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n246), .A2(new_n313), .A3(KEYINPUT4), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n352), .A2(new_n356), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT5), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n251), .A2(new_n348), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n349), .A2(new_n351), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n357), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n251), .B(new_n287), .C1(new_n315), .C2(KEYINPUT77), .ZN(new_n366));
  INV_X1    g165(.A(new_n355), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n360), .B(new_n357), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT4), .B1(new_n246), .B2(new_n313), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n351), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(KEYINPUT4), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G1gat), .B(G29gat), .Z(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G57gat), .B(G85gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n365), .A2(new_n373), .A3(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n359), .A2(new_n364), .B1(new_n369), .B2(new_n372), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(new_n379), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n346), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n381), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n383), .B2(new_n379), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n365), .A2(new_n373), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n378), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(KEYINPUT81), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n384), .A2(new_n386), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n385), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n235), .A2(new_n288), .ZN(new_n393));
  NAND2_X1  g192(.A1(G226gat), .A2(G233gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n235), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n325), .A3(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(G8gat), .B(G36gat), .Z(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT73), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n396), .B1(new_n235), .B2(new_n288), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT72), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n235), .A2(KEYINPUT72), .A3(new_n396), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n308), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n398), .B(new_n402), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n235), .A2(KEYINPUT72), .A3(new_n396), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT72), .B1(new_n235), .B2(new_n396), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n395), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n397), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(new_n403), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n412), .A2(new_n308), .B1(new_n414), .B2(new_n325), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n402), .B(KEYINPUT74), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n409), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT30), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n409), .A2(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n343), .A2(new_n345), .A3(new_n392), .A4(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT35), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT85), .B1(new_n383), .B2(new_n379), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n388), .A2(new_n426), .A3(new_n378), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n387), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n391), .ZN(new_n429));
  AND4_X1   g228(.A1(new_n424), .A2(new_n422), .A3(new_n429), .A4(new_n344), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT69), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n266), .A2(new_n431), .A3(new_n340), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n260), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n423), .A2(KEYINPUT35), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n344), .B1(new_n392), .B2(new_n422), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT36), .B1(new_n432), .B2(new_n433), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT36), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n266), .B2(new_n340), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n251), .A2(new_n347), .A3(new_n348), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT78), .B1(new_n246), .B2(new_n313), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT4), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n370), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n356), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n363), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n447), .B(KEYINPUT39), .C1(new_n363), .C2(new_n362), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n449), .A3(new_n363), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n450), .A2(new_n451), .A3(new_n379), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n450), .B2(new_n379), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT40), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n448), .B(KEYINPUT40), .C1(new_n452), .C2(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n419), .A2(new_n421), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n425), .A2(new_n427), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n402), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n398), .B1(new_n407), .B2(new_n408), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n461), .B1(new_n462), .B2(KEYINPUT37), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT37), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n415), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT38), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n395), .A2(new_n397), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n407), .A2(new_n408), .B1(new_n468), .B2(new_n324), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n469), .B2(new_n464), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT38), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n416), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n415), .B2(new_n464), .ZN(new_n473));
  OAI22_X1  g272(.A1(new_n412), .A2(new_n308), .B1(new_n414), .B2(new_n325), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(KEYINPUT86), .A3(KEYINPUT37), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n470), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n466), .A2(new_n476), .A3(new_n409), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n460), .B(new_n344), .C1(new_n429), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n441), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n436), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n481), .B(KEYINPUT13), .Z(new_n482));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n483));
  INV_X1    g282(.A(G29gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n486));
  AOI21_X1  g285(.A(G36gat), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G36gat), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n483), .A2(new_n488), .A3(G29gat), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n490), .B(new_n492), .C1(KEYINPUT88), .C2(new_n494), .ZN(new_n495));
  OAI22_X1  g294(.A1(new_n487), .A2(new_n489), .B1(KEYINPUT15), .B2(new_n491), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n487), .A2(new_n489), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n496), .B(new_n493), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  INV_X1    g300(.A(G1gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT16), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n501), .A2(G1gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G8gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n500), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n506), .B(G8gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n499), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n482), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(KEYINPUT17), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n495), .A2(new_n499), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n510), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n508), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n481), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n519), .A2(KEYINPUT89), .A3(new_n481), .A4(new_n520), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT90), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n521), .B2(new_n524), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n521), .A2(new_n527), .A3(new_n524), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n515), .B(new_n526), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G197gat), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT11), .B(G169gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(KEYINPUT12), .Z(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  OR3_X1    g336(.A1(new_n521), .A2(new_n527), .A3(new_n524), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n528), .ZN(new_n539));
  INV_X1    g338(.A(new_n536), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n539), .A2(new_n540), .A3(new_n526), .A4(new_n515), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G99gat), .B(G106gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT8), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n546), .B1(G99gat), .B2(G106gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT96), .B(G92gat), .ZN(new_n548));
  INV_X1    g347(.A(G85gat), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(G85gat), .A3(G92gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n545), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(G92gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT96), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT96), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(G92gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n560), .A3(new_n549), .ZN(new_n561));
  INV_X1    g360(.A(G99gat), .ZN(new_n562));
  INV_X1    g361(.A(G106gat), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT8), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND4_X1   g363(.A1(new_n545), .A2(new_n561), .A3(new_n555), .A4(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n556), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n516), .A2(new_n518), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n500), .A2(new_n566), .B1(KEYINPUT41), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT97), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n568), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n544), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n568), .A2(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT97), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n577), .A3(new_n543), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT95), .ZN(new_n580));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  NAND3_X1  g381(.A1(new_n574), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n583), .A2(KEYINPUT98), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(KEYINPUT98), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT99), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n574), .A2(new_n578), .ZN(new_n587));
  INV_X1    g386(.A(new_n582), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI211_X1 g388(.A(KEYINPUT99), .B(new_n582), .C1(new_n574), .C2(new_n578), .ZN(new_n590));
  OAI22_X1  g389(.A1(new_n584), .A2(new_n585), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT21), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT9), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n595), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n597), .B(new_n596), .C1(new_n594), .C2(new_n599), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n510), .B1(new_n593), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n593), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n604), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT93), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT92), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n610), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G183gat), .B(G211gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT94), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n613), .B(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n608), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n608), .A2(new_n616), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n603), .B1(new_n556), .B2(new_n565), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n561), .A2(new_n555), .A3(new_n564), .ZN(new_n622));
  INV_X1    g421(.A(new_n545), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n561), .A2(new_n555), .A3(new_n545), .A4(new_n564), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n624), .A2(new_n602), .A3(new_n601), .A4(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n603), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n566), .A2(KEYINPUT100), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n627), .A2(new_n629), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT101), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n635), .A2(new_n638), .A3(new_n633), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n634), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n632), .B1(new_n640), .B2(new_n631), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n632), .B(new_n644), .C1(new_n640), .C2(new_n631), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n592), .A2(new_n619), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n480), .A2(new_n542), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n392), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n502), .ZN(G1324gat));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n655));
  INV_X1    g454(.A(new_n652), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT16), .B(G8gat), .Z(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n458), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(G8gat), .B1(new_n652), .B2(new_n422), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(KEYINPUT102), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(KEYINPUT102), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n655), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n658), .B(KEYINPUT42), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n666), .A2(KEYINPUT103), .A3(new_n663), .A4(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(G1325gat));
  NOR2_X1   g467(.A1(new_n438), .A2(new_n440), .ZN(new_n669));
  OAI21_X1  g468(.A(G15gat), .B1(new_n652), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n435), .B1(new_n478), .B2(new_n441), .ZN(new_n671));
  INV_X1    g470(.A(new_n542), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n434), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n650), .A2(G15gat), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n670), .A2(new_n676), .ZN(G1326gat));
  INV_X1    g476(.A(new_n344), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n656), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT104), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n680), .B(new_n682), .ZN(G1327gat));
  NOR3_X1   g482(.A1(new_n592), .A2(new_n619), .A3(new_n648), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n480), .A2(new_n542), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n392), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n484), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT45), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n619), .B(KEYINPUT105), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n542), .A3(new_n649), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n392), .A2(new_n422), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n678), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n669), .A2(new_n693), .ZN(new_n694));
  AND4_X1   g493(.A1(new_n456), .A2(new_n457), .A3(new_n459), .A4(new_n458), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n344), .B1(new_n477), .B2(new_n429), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n694), .A2(new_n697), .A3(KEYINPUT106), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n441), .B2(new_n478), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n436), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT107), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT106), .B1(new_n694), .B2(new_n697), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n441), .A2(new_n699), .A3(new_n478), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n435), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n592), .A2(KEYINPUT44), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n702), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT44), .B1(new_n671), .B2(new_n592), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n691), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(new_n687), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n689), .B1(new_n712), .B2(new_n484), .ZN(G1328gat));
  NAND2_X1  g512(.A1(new_n458), .A2(new_n488), .ZN(new_n714));
  OR3_X1    g513(.A1(new_n685), .A2(KEYINPUT108), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT108), .B1(new_n685), .B2(new_n714), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT46), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n711), .A2(new_n458), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n488), .B2(new_n719), .ZN(G1329gat));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721));
  INV_X1    g520(.A(G43gat), .ZN(new_n722));
  INV_X1    g521(.A(new_n669), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n711), .B2(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n685), .A2(G43gat), .A3(new_n674), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n725), .ZN(new_n727));
  AOI211_X1 g526(.A(new_n669), .B(new_n691), .C1(new_n709), .C2(new_n710), .ZN(new_n728));
  OAI211_X1 g527(.A(KEYINPUT47), .B(new_n727), .C1(new_n728), .C2(new_n722), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(G1330gat));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  INV_X1    g530(.A(G50gat), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(new_n711), .B2(new_n678), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n678), .A2(new_n732), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT109), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n686), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n731), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  AOI211_X1 g537(.A(new_n344), .B(new_n691), .C1(new_n709), .C2(new_n710), .ZN(new_n739));
  OAI211_X1 g538(.A(KEYINPUT48), .B(new_n736), .C1(new_n739), .C2(new_n732), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(G1331gat));
  NOR2_X1   g540(.A1(new_n705), .A2(new_n706), .ZN(new_n742));
  AOI211_X1 g541(.A(KEYINPUT107), .B(new_n435), .C1(new_n703), .C2(new_n704), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n619), .ZN(new_n745));
  NOR4_X1   g544(.A1(new_n591), .A2(new_n542), .A3(new_n649), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n687), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n458), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT49), .B(G64gat), .Z(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n751), .B2(new_n753), .ZN(G1333gat));
  OAI21_X1  g553(.A(G71gat), .B1(new_n747), .B2(new_n669), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n674), .A2(G71gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n744), .A2(new_n746), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n755), .A2(KEYINPUT50), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n748), .A2(new_n678), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g563(.A1(new_n392), .A2(new_n649), .A3(G85gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n672), .A2(new_n591), .A3(new_n745), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n701), .A2(new_n766), .A3(KEYINPUT51), .A4(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n705), .B2(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n703), .A2(new_n704), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n767), .B1(new_n773), .B2(new_n436), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n766), .B1(new_n774), .B2(KEYINPUT51), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n765), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n672), .A2(new_n745), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n649), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n709), .B2(new_n710), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n687), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n776), .B1(new_n781), .B2(new_n549), .ZN(G1336gat));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n422), .B(new_n779), .C1(new_n709), .C2(new_n710), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n548), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n649), .A2(new_n422), .A3(G92gat), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT111), .Z(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n772), .B2(new_n775), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g590(.A(KEYINPUT112), .B(new_n788), .C1(new_n772), .C2(new_n775), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n774), .A2(KEYINPUT51), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n787), .B1(new_n794), .B2(new_n771), .ZN(new_n795));
  INV_X1    g594(.A(new_n708), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n742), .A2(new_n743), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n710), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n458), .B(new_n778), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n548), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n795), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n785), .A2(new_n793), .B1(new_n801), .B2(new_n783), .ZN(G1337gat));
  NOR2_X1   g601(.A1(new_n649), .A2(G99gat), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n434), .B(new_n803), .C1(new_n772), .C2(new_n775), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n780), .A2(new_n723), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n562), .ZN(G1338gat));
  OAI211_X1 g605(.A(new_n678), .B(new_n778), .C1(new_n797), .C2(new_n798), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n794), .A2(new_n771), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n649), .A2(G106gat), .A3(new_n344), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n807), .A2(G106gat), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n563), .B1(new_n780), .B2(new_n678), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n809), .B1(new_n772), .B2(new_n775), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n811), .ZN(new_n814));
  OAI22_X1  g613(.A1(new_n810), .A2(new_n811), .B1(new_n812), .B2(new_n814), .ZN(G1339gat));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n637), .A2(new_n639), .ZN(new_n817));
  INV_X1    g616(.A(new_n634), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n631), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n638), .B1(new_n635), .B2(new_n633), .ZN(new_n820));
  AOI211_X1 g619(.A(KEYINPUT101), .B(KEYINPUT10), .C1(new_n627), .C2(new_n629), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n818), .B(new_n631), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT54), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n826), .A3(new_n630), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n645), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n816), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(KEYINPUT54), .B(new_n822), .C1(new_n640), .C2(new_n631), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n645), .A4(new_n827), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n542), .A2(new_n647), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n509), .A2(new_n512), .A3(new_n482), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT113), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n481), .B1(new_n519), .B2(new_n520), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n535), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n541), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n648), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n591), .B1(new_n832), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n831), .A2(new_n647), .ZN(new_n840));
  AND4_X1   g639(.A1(new_n591), .A2(new_n837), .A3(new_n840), .A4(new_n829), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n690), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n592), .A2(new_n672), .A3(new_n619), .A4(new_n649), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n674), .A2(new_n678), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n392), .A2(new_n458), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(G113gat), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n848), .A2(new_n849), .A3(new_n672), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n392), .B1(new_n842), .B2(new_n843), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n343), .A2(new_n345), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n853), .A2(KEYINPUT114), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n458), .B1(new_n853), .B2(KEYINPUT114), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n542), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n850), .B1(new_n857), .B2(new_n849), .ZN(G1340gat));
  NOR2_X1   g657(.A1(new_n649), .A2(G120gat), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G120gat), .B1(new_n848), .B2(new_n649), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1341gat));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n238), .A3(new_n690), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT116), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n856), .A2(new_n619), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n238), .ZN(G1342gat));
  AND2_X1   g666(.A1(new_n591), .A2(new_n236), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n856), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT56), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n871), .A3(new_n868), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n848), .B2(new_n592), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(G1343gat));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n669), .A2(new_n847), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n344), .B1(new_n842), .B2(new_n843), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT55), .B1(new_n819), .B2(new_n823), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n647), .B1(new_n881), .B2(new_n828), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n827), .A2(new_n645), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT55), .B1(new_n883), .B2(new_n830), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n880), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n829), .A2(KEYINPUT117), .A3(new_n647), .A4(new_n831), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n542), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n591), .B1(new_n887), .B2(new_n838), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n745), .B1(new_n888), .B2(new_n841), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n344), .B1(new_n889), .B2(new_n843), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n879), .B(new_n542), .C1(new_n878), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G141gat), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n669), .A2(new_n678), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT119), .Z(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n851), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n458), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n897), .B1(new_n896), .B2(new_n895), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n542), .A2(new_n267), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n875), .B(new_n892), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n891), .A2(new_n901), .A3(G141gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n891), .B2(G141gat), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n895), .A2(new_n458), .A3(new_n899), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n900), .B1(new_n905), .B2(new_n875), .ZN(G1344gat));
  OAI21_X1  g705(.A(new_n879), .B1(new_n878), .B2(new_n890), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  AOI211_X1 g707(.A(KEYINPUT59), .B(new_n268), .C1(new_n908), .C2(new_n648), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n889), .A2(new_n843), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT121), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n889), .A2(new_n913), .A3(new_n843), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n344), .A2(KEYINPUT57), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n877), .A2(new_n878), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n876), .A2(new_n649), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n910), .B1(new_n919), .B2(G148gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n648), .A2(new_n268), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n909), .A2(new_n920), .B1(new_n898), .B2(new_n921), .ZN(G1345gat));
  OAI21_X1  g721(.A(G155gat), .B1(new_n907), .B2(new_n690), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n619), .A2(new_n276), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n898), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT122), .ZN(G1346gat));
  OR2_X1    g725(.A1(new_n898), .A2(new_n592), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n592), .A2(new_n277), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n927), .A2(new_n277), .B1(new_n908), .B2(new_n928), .ZN(G1347gat));
  NAND2_X1  g728(.A1(new_n392), .A2(new_n458), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT123), .Z(new_n931));
  NAND2_X1  g730(.A1(new_n846), .A2(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(new_n209), .A3(new_n672), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n687), .B1(new_n842), .B2(new_n843), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(new_n458), .A3(new_n852), .ZN(new_n935));
  AOI21_X1  g734(.A(G169gat), .B1(new_n935), .B2(new_n542), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n933), .A2(new_n936), .ZN(G1348gat));
  OAI21_X1  g736(.A(G176gat), .B1(new_n932), .B2(new_n649), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n210), .A3(new_n648), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1349gat));
  OAI21_X1  g739(.A(G183gat), .B1(new_n932), .B2(new_n690), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n935), .A2(new_n229), .A3(new_n619), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n935), .A2(new_n228), .A3(new_n591), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n844), .A2(new_n591), .A3(new_n845), .A4(new_n931), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(G190gat), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n947), .B1(new_n946), .B2(G190gat), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n949), .A2(new_n950), .A3(KEYINPUT61), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n946), .A2(G190gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT124), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n952), .B1(new_n954), .B2(new_n948), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n945), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g757(.A(KEYINPUT125), .B(new_n945), .C1(new_n951), .C2(new_n955), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1351gat));
  NOR2_X1   g759(.A1(new_n893), .A2(new_n422), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n934), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n542), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n931), .A2(new_n669), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n916), .A2(new_n917), .A3(new_n965), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n542), .A2(G197gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(G1352gat));
  NAND4_X1  g767(.A1(new_n916), .A2(new_n648), .A3(new_n917), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G204gat), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n649), .A2(G204gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n934), .A2(new_n961), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT62), .Z(new_n973));
  NAND2_X1  g772(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n970), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1353gat));
  OR3_X1    g777(.A1(new_n962), .A2(G211gat), .A3(new_n745), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n916), .A2(new_n619), .A3(new_n917), .A4(new_n965), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n980), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n980), .B2(G211gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  AOI21_X1  g782(.A(G218gat), .B1(new_n963), .B2(new_n591), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n591), .A2(G218gat), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT127), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n984), .B1(new_n966), .B2(new_n986), .ZN(G1355gat));
endmodule


