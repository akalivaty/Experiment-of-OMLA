//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT79), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G137), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT24), .B(G110), .Z(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT66), .B(G119), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(new_n195), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT75), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT75), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT66), .A2(G119), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT66), .A2(G119), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G128), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n200), .B1(new_n204), .B2(new_n196), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n194), .B1(new_n199), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n207), .B1(new_n203), .B2(G128), .ZN(new_n208));
  INV_X1    g022(.A(new_n196), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(new_n203), .B2(G128), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n210), .B2(new_n207), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G110), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G140), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G125), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT16), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT77), .ZN(new_n218));
  INV_X1    g032(.A(G125), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n218), .B(G140), .C1(new_n219), .C2(KEYINPUT76), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT77), .B1(new_n214), .B2(G125), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT76), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(new_n214), .A3(G125), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n220), .A2(new_n221), .A3(new_n223), .A4(KEYINPUT16), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n217), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(G146), .B(new_n217), .C1(new_n226), .C2(new_n227), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n213), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G110), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n233), .B(new_n208), .C1(new_n210), .C2(new_n207), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n198), .A2(KEYINPUT75), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n204), .A2(new_n200), .A3(new_n196), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n237), .B2(new_n194), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n219), .A2(G140), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n215), .A3(new_n229), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n238), .A2(new_n231), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n193), .B1(new_n232), .B2(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n237), .A2(new_n194), .B1(new_n211), .B2(G110), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n220), .A2(new_n221), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n244), .A2(KEYINPUT78), .A3(KEYINPUT16), .A4(new_n223), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n224), .A2(new_n225), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(G146), .B1(new_n247), .B2(new_n217), .ZN(new_n248));
  AOI211_X1 g062(.A(new_n229), .B(new_n216), .C1(new_n245), .C2(new_n246), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n243), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n238), .A2(new_n231), .A3(new_n240), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(new_n192), .ZN(new_n252));
  AOI21_X1  g066(.A(G902), .B1(new_n242), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n187), .B1(new_n253), .B2(KEYINPUT80), .ZN(new_n254));
  INV_X1    g068(.A(G902), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n250), .A2(new_n251), .A3(new_n192), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n192), .B1(new_n250), .B2(new_n251), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT80), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT25), .ZN(new_n260));
  INV_X1    g074(.A(G217), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(G234), .B2(new_n255), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n254), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n242), .A2(new_n252), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n262), .A2(G902), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(G472), .A2(G902), .ZN(new_n268));
  INV_X1    g082(.A(G113), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT2), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G113), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OR2_X1    g087(.A1(KEYINPUT66), .A2(G119), .ZN(new_n274));
  NAND2_X1  g088(.A1(KEYINPUT66), .A2(G119), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(G116), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G116), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G119), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n273), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n276), .A2(new_n278), .A3(new_n273), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT65), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(KEYINPUT65), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT11), .ZN(new_n287));
  INV_X1    g101(.A(G134), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(G137), .ZN(new_n289));
  INV_X1    g103(.A(G137), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT11), .A3(G134), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(G137), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G131), .ZN(new_n294));
  INV_X1    g108(.A(G131), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n289), .A2(new_n291), .A3(new_n295), .A4(new_n292), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n229), .A2(G143), .ZN(new_n298));
  INV_X1    g112(.A(G143), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G146), .ZN(new_n300));
  AND2_X1   g114(.A1(KEYINPUT0), .A2(G128), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n298), .B2(new_n300), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT0), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n195), .A3(KEYINPUT64), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(KEYINPUT0), .B2(G128), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n302), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n297), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n292), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n288), .A2(G137), .ZN(new_n312));
  OAI21_X1  g126(.A(G131), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT1), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n298), .A2(new_n300), .A3(new_n314), .A4(G128), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT1), .B1(new_n299), .B2(G146), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n317), .A2(G128), .B1(new_n298), .B2(new_n300), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n296), .B(new_n313), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  AOI211_X1 g133(.A(new_n284), .B(new_n286), .C1(new_n310), .C2(new_n319), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n310), .A2(KEYINPUT65), .A3(new_n283), .A4(new_n319), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n282), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n324));
  INV_X1    g138(.A(G237), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n188), .A3(G210), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n324), .B(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT26), .B(G101), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n276), .A2(new_n278), .A3(new_n273), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(new_n279), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n310), .A2(new_n332), .A3(new_n319), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT68), .B(KEYINPUT31), .Z(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n323), .A2(new_n330), .A3(new_n333), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n310), .A2(new_n319), .ZN(new_n337));
  INV_X1    g151(.A(new_n284), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n285), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n332), .B1(new_n339), .B2(new_n321), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n310), .A2(new_n332), .A3(new_n319), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n340), .A2(new_n329), .A3(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(KEYINPUT68), .A2(KEYINPUT31), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n336), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n332), .B1(new_n310), .B2(new_n319), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT28), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT69), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT69), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n348), .B(KEYINPUT28), .C1(new_n341), .C2(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT70), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n341), .B2(KEYINPUT28), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n333), .A2(KEYINPUT70), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n330), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(KEYINPUT32), .B(new_n268), .C1(new_n344), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT74), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n323), .A2(new_n330), .A3(new_n333), .ZN(new_n360));
  INV_X1    g174(.A(new_n343), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n355), .B1(new_n347), .B2(new_n349), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n362), .B(new_n336), .C1(new_n363), .C2(new_n330), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT74), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT32), .A4(new_n268), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n268), .B1(new_n344), .B2(new_n357), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT72), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n371), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT72), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n367), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n363), .A2(new_n329), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n340), .A2(new_n341), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n329), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n330), .A2(KEYINPUT29), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n356), .A2(new_n346), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT73), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n356), .A2(KEYINPUT73), .A3(new_n346), .A4(new_n380), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n255), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G472), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n267), .B1(new_n375), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G469), .ZN(new_n388));
  XNOR2_X1  g202(.A(G110), .B(G140), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n188), .A2(G227), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n389), .B(new_n390), .Z(new_n391));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n392), .B1(new_n393), .B2(G107), .ZN(new_n394));
  INV_X1    g208(.A(G107), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT3), .A3(G104), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G101), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(G107), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT81), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n393), .A3(G107), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n397), .A2(new_n398), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT82), .B1(new_n393), .B2(G107), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n395), .A3(G104), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n406), .A3(new_n399), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G101), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n316), .A2(new_n318), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT83), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n317), .A2(G128), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n298), .A2(new_n300), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n315), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n415), .A2(new_n416), .A3(new_n403), .A4(new_n408), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n403), .A2(new_n408), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n403), .B2(new_n408), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n410), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT12), .B1(new_n423), .B2(new_n297), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT12), .ZN(new_n425));
  INV_X1    g239(.A(new_n297), .ZN(new_n426));
  AOI211_X1 g240(.A(new_n425), .B(new_n426), .C1(new_n418), .C2(new_n422), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n409), .A2(KEYINPUT84), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT10), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n410), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n403), .A2(new_n408), .A3(new_n419), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n395), .A2(KEYINPUT3), .A3(G104), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT3), .B1(new_n395), .B2(G104), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n400), .B(new_n402), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G101), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT4), .A3(new_n403), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n439), .A3(G101), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n309), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n433), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT10), .B1(new_n411), .B2(new_n417), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n442), .A2(new_n443), .A3(new_n297), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n391), .B1(new_n428), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n418), .A2(new_n430), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n446), .A2(new_n426), .A3(new_n433), .A4(new_n441), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n297), .B1(new_n442), .B2(new_n443), .ZN(new_n448));
  INV_X1    g262(.A(new_n391), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n388), .B1(new_n451), .B2(new_n255), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n447), .B(new_n449), .C1(new_n424), .C2(new_n427), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT85), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n449), .B1(new_n447), .B2(new_n448), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI211_X1 g270(.A(KEYINPUT85), .B(new_n449), .C1(new_n447), .C2(new_n448), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n388), .B(new_n255), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT86), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n433), .A2(new_n441), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n426), .B1(new_n460), .B2(new_n446), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n391), .B1(new_n461), .B2(new_n444), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT85), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n455), .A2(new_n454), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n453), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n388), .A4(new_n255), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n452), .B1(new_n459), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT9), .B(G234), .ZN(new_n469));
  OAI21_X1  g283(.A(G221), .B1(new_n469), .B2(G902), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT87), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G214), .B1(G237), .B2(G902), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n276), .A2(KEYINPUT5), .A3(new_n278), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT5), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n274), .A2(new_n475), .A3(G116), .A4(new_n275), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n476), .A2(G113), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n331), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n429), .A3(new_n432), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n438), .A2(new_n282), .A3(new_n440), .ZN(new_n480));
  XNOR2_X1  g294(.A(G110), .B(G122), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT88), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n479), .A2(new_n480), .ZN(new_n484));
  INV_X1    g298(.A(new_n481), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT88), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n479), .A2(new_n480), .A3(new_n487), .A4(new_n481), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(KEYINPUT89), .A3(new_n485), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n481), .B1(new_n479), .B2(new_n480), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(KEYINPUT89), .A3(KEYINPUT6), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n309), .A2(G125), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n415), .A2(new_n219), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G224), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(G953), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n498), .B(new_n500), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G210), .B1(G237), .B2(G902), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n498), .B(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n409), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n479), .B1(new_n507), .B2(new_n478), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n481), .B(KEYINPUT8), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n483), .A2(new_n488), .ZN(new_n511));
  AOI21_X1  g325(.A(G902), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n502), .A2(new_n503), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n503), .B1(new_n502), .B2(new_n512), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n473), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT90), .ZN(new_n516));
  INV_X1    g330(.A(new_n473), .ZN(new_n517));
  INV_X1    g331(.A(new_n503), .ZN(new_n518));
  INV_X1    g332(.A(new_n501), .ZN(new_n519));
  AND4_X1   g333(.A1(KEYINPUT89), .A2(new_n484), .A3(KEYINPUT6), .A4(new_n485), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT6), .B1(new_n493), .B2(KEYINPUT89), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n519), .B1(new_n522), .B2(new_n489), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n510), .A2(new_n511), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n255), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n518), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n502), .A2(new_n503), .A3(new_n512), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n517), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G475), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n325), .A2(new_n188), .A3(G214), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n299), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n325), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(G131), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n295), .B1(new_n534), .B2(new_n535), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n532), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n538), .A2(new_n532), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n230), .A2(new_n541), .A3(new_n231), .ZN(new_n542));
  NAND2_X1  g356(.A1(KEYINPUT18), .A2(G131), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n536), .B(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n220), .A2(new_n223), .A3(new_n221), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G146), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n240), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT91), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n536), .B(new_n543), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT91), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n548), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G113), .B(G122), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(new_n393), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n542), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT93), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT93), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n542), .A2(new_n554), .A3(new_n559), .A4(new_n556), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n542), .A2(new_n554), .ZN(new_n562));
  INV_X1    g376(.A(new_n556), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n531), .B1(new_n565), .B2(new_n255), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT19), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n239), .A2(new_n215), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT92), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n546), .A2(KEYINPUT19), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n569), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI22_X1  g387(.A1(new_n573), .A2(G146), .B1(new_n538), .B2(new_n537), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n554), .B1(new_n249), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n558), .A2(new_n560), .B1(new_n563), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(G475), .A2(G902), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT20), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n563), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n561), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT20), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n577), .B(KEYINPUT94), .Z(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n566), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n469), .A2(new_n261), .A3(G953), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT95), .B1(new_n277), .B2(G122), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n589));
  INV_X1    g403(.A(G122), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n590), .A3(G116), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n395), .B1(new_n592), .B2(KEYINPUT14), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n592), .B1(G116), .B2(new_n590), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI221_X1 g409(.A(new_n592), .B1(KEYINPUT14), .B2(new_n395), .C1(G116), .C2(new_n590), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT96), .B1(new_n299), .B2(G128), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n195), .A3(G143), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n299), .A2(G128), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n602), .B1(new_n601), .B2(new_n603), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n288), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n601), .A2(new_n603), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT97), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(G134), .A3(new_n604), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n597), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT13), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n603), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n299), .A2(KEYINPUT13), .A3(G128), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n601), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(G134), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n588), .A2(new_n591), .B1(new_n277), .B2(G122), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n617), .A2(new_n395), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n395), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(G134), .B1(new_n609), .B2(new_n604), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n587), .B1(new_n611), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n595), .A2(new_n596), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n605), .A2(new_n288), .A3(new_n606), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n621), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n607), .B(new_n616), .C1(new_n619), .C2(new_n618), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n586), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n623), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(KEYINPUT98), .B(new_n587), .C1(new_n611), .C2(new_n622), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n255), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT99), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n630), .A2(new_n634), .A3(new_n255), .A4(new_n631), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(G478), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(KEYINPUT15), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n638), .B1(new_n632), .B2(KEYINPUT99), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(G952), .ZN(new_n643));
  AOI211_X1 g457(.A(G953), .B(new_n643), .C1(G234), .C2(G237), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT21), .B(G898), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT100), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n255), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT101), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n642), .A2(new_n651), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n516), .A2(new_n530), .A3(new_n585), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n459), .A2(new_n467), .ZN(new_n654));
  INV_X1    g468(.A(new_n452), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT87), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n657), .A3(new_n470), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n387), .A2(new_n472), .A3(new_n653), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G101), .ZN(G3));
  NAND2_X1  g474(.A1(new_n364), .A2(new_n255), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G472), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n368), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n267), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n658), .A2(new_n472), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n528), .A2(new_n650), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT33), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n630), .A2(new_n668), .A3(new_n631), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n623), .A2(new_n628), .A3(KEYINPUT33), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n669), .A2(new_n670), .A3(G478), .A4(new_n255), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n632), .A2(new_n637), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n667), .B1(new_n585), .B2(new_n674), .ZN(new_n675));
  AOI22_X1  g489(.A1(new_n558), .A2(new_n560), .B1(new_n563), .B2(new_n562), .ZN(new_n676));
  OAI21_X1  g490(.A(G475), .B1(new_n676), .B2(G902), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n582), .B1(new_n581), .B2(new_n577), .ZN(new_n678));
  INV_X1    g492(.A(new_n583), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n576), .A2(KEYINPUT20), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n677), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(KEYINPUT102), .A3(new_n673), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n675), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n665), .A2(new_n666), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT34), .B(G104), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G6));
  AOI21_X1  g500(.A(new_n566), .B1(new_n639), .B2(new_n641), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n579), .A2(new_n688), .ZN(new_n689));
  OAI211_X1 g503(.A(KEYINPUT103), .B(KEYINPUT20), .C1(new_n576), .C2(new_n578), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n581), .A2(new_n582), .A3(new_n577), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n665), .A2(new_n666), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT35), .B(G107), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G9));
  NAND2_X1  g510(.A1(new_n250), .A2(new_n251), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n192), .A2(KEYINPUT36), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n265), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n263), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n663), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n653), .A2(new_n658), .A3(new_n472), .A4(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT37), .B(G110), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G12));
  AOI21_X1  g520(.A(new_n515), .B1(new_n375), .B2(new_n386), .ZN(new_n707));
  INV_X1    g521(.A(G900), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n644), .B1(new_n648), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n692), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n640), .B1(new_n636), .B2(new_n638), .ZN(new_n712));
  NOR4_X1   g526(.A1(new_n711), .A2(new_n702), .A3(new_n566), .A4(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n707), .A2(new_n472), .A3(new_n658), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G128), .ZN(G30));
  AOI21_X1  g529(.A(new_n471), .B1(new_n654), .B2(new_n655), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n657), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n468), .A2(KEYINPUT87), .A3(new_n471), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n709), .B(KEYINPUT39), .Z(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n721), .A2(KEYINPUT40), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(KEYINPUT40), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n377), .A2(new_n329), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n341), .A2(new_n345), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n255), .B1(new_n725), .B2(new_n330), .ZN(new_n726));
  OAI21_X1  g540(.A(G472), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n375), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n526), .A2(new_n527), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n681), .A2(new_n642), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n732), .A2(new_n517), .A3(new_n701), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n728), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n722), .A2(new_n723), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G143), .ZN(G45));
  NAND2_X1  g550(.A1(new_n681), .A2(new_n673), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n737), .A2(new_n702), .A3(new_n709), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n707), .A2(new_n472), .A3(new_n658), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  AOI21_X1  g554(.A(new_n666), .B1(new_n675), .B2(new_n682), .ZN(new_n741));
  INV_X1    g555(.A(new_n367), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n374), .A2(new_n372), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n386), .ZN(new_n744));
  INV_X1    g558(.A(new_n267), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n388), .B1(new_n465), .B2(new_n255), .ZN(new_n746));
  AOI211_X1 g560(.A(new_n471), .B(new_n746), .C1(new_n459), .C2(new_n467), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n741), .A2(new_n744), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n387), .A2(KEYINPUT105), .A3(new_n741), .A4(new_n747), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT41), .B(G113), .Z(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT106), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n752), .B(new_n754), .ZN(G15));
  AND3_X1   g569(.A1(new_n263), .A2(new_n266), .A3(new_n650), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n756), .A2(new_n687), .A3(new_n692), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n744), .A2(new_n747), .A3(new_n757), .A4(new_n528), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n746), .B1(new_n459), .B2(new_n467), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n761), .A2(new_n470), .A3(new_n528), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n762), .A2(KEYINPUT107), .A3(new_n744), .A4(new_n757), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G116), .ZN(G18));
  NOR3_X1   g579(.A1(new_n681), .A2(new_n642), .A3(new_n651), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n762), .A2(new_n744), .A3(new_n766), .A4(new_n701), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  NAND2_X1  g582(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n681), .A2(new_n642), .A3(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n769), .A2(new_n528), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n330), .B1(new_n356), .B2(new_n346), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n268), .B1(new_n344), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n662), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n775), .A2(new_n267), .A3(new_n651), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n772), .A2(new_n747), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G122), .ZN(G24));
  NOR2_X1   g592(.A1(new_n737), .A2(new_n709), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n775), .A2(new_n702), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n762), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G125), .ZN(G27));
  AND2_X1   g597(.A1(new_n386), .A2(new_n358), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT32), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n368), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n267), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n729), .A2(new_n517), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n789), .A2(new_n468), .A3(KEYINPUT109), .A4(new_n471), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n716), .B2(new_n788), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n787), .B(new_n779), .C1(new_n790), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT42), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n716), .A2(new_n788), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT109), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n716), .A2(new_n788), .A3(new_n791), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT42), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n387), .A4(new_n779), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT110), .B(G131), .Z(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(G33));
  INV_X1    g617(.A(new_n711), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n798), .A2(new_n387), .A3(new_n687), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  NAND2_X1  g620(.A1(new_n585), .A2(new_n673), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT43), .Z(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n663), .A3(new_n701), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT44), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n451), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n445), .A2(KEYINPUT45), .A3(new_n450), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n812), .A2(G469), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT46), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n388), .A2(new_n255), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n815), .B1(new_n814), .B2(new_n816), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n818), .A3(new_n654), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n470), .ZN(new_n820));
  INV_X1    g634(.A(new_n720), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n810), .A2(new_n788), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n820), .B(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n779), .A2(new_n267), .A3(new_n788), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n744), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n827), .B1(new_n826), .B2(new_n829), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G140), .ZN(G42));
  AOI21_X1  g648(.A(new_n529), .B1(new_n729), .B2(new_n473), .ZN(new_n835));
  AOI211_X1 g649(.A(KEYINPUT90), .B(new_n517), .C1(new_n526), .C2(new_n527), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n681), .A2(new_n712), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(KEYINPUT114), .A3(new_n650), .A4(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n516), .A2(new_n530), .A3(new_n838), .A4(new_n650), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n704), .B1(new_n843), .B2(new_n665), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT115), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n584), .A2(new_n579), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n674), .B1(new_n846), .B2(new_n677), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n516), .A2(new_n530), .A3(new_n650), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n658), .A3(new_n472), .A4(new_n664), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n659), .A2(new_n767), .A3(new_n777), .A4(new_n849), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n750), .A2(new_n751), .B1(new_n760), .B2(new_n763), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n852), .B(new_n704), .C1(new_n843), .C2(new_n665), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n845), .A2(new_n850), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n702), .A2(new_n642), .A3(new_n566), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n744), .A2(new_n804), .A3(new_n788), .A4(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n798), .A2(new_n781), .B1(new_n719), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n794), .A3(new_n800), .A4(new_n805), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n701), .A2(new_n709), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n772), .A2(new_n716), .A3(new_n728), .A4(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n714), .A2(new_n739), .A3(new_n861), .A4(new_n782), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT52), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n862), .A2(KEYINPUT52), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n859), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n762), .A2(new_n779), .A3(new_n780), .ZN(new_n870));
  AOI211_X1 g684(.A(KEYINPUT72), .B(new_n370), .C1(new_n364), .C2(new_n268), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n369), .B1(new_n368), .B2(new_n371), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n359), .B(new_n366), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n386), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n528), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n717), .A2(new_n875), .A3(new_n718), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n870), .B1(new_n876), .B2(new_n713), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n739), .A4(new_n861), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n879), .A2(new_n880), .A3(new_n863), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n879), .B2(new_n863), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n859), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n869), .B1(new_n868), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n868), .ZN(new_n886));
  XOR2_X1   g700(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n887));
  NAND3_X1  g701(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n866), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n745), .A2(new_n644), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n775), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n808), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n747), .ZN(new_n894));
  NOR4_X1   g708(.A1(new_n893), .A2(new_n473), .A3(new_n731), .A4(new_n894), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT50), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n728), .A2(new_n891), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n894), .A2(new_n789), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n899), .A2(new_n681), .A3(new_n673), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n898), .A2(new_n644), .A3(new_n808), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n780), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n761), .B(KEYINPUT113), .Z(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n470), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n826), .B2(KEYINPUT118), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(KEYINPUT118), .B2(new_n826), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n893), .A2(new_n789), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT51), .B1(new_n903), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n826), .B2(new_n905), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n896), .A2(KEYINPUT51), .A3(new_n902), .A4(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n808), .A2(new_n762), .A3(new_n892), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n643), .A2(G953), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n913), .B(new_n914), .C1(new_n899), .C2(new_n683), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT119), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n901), .A2(new_n787), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(KEYINPUT120), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(KEYINPUT120), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(KEYINPUT48), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT48), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n917), .A2(KEYINPUT120), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n912), .A2(new_n916), .A3(new_n920), .A4(new_n922), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n910), .A2(new_n923), .ZN(new_n924));
  OAI22_X1  g738(.A1(new_n890), .A2(new_n924), .B1(G952), .B2(G953), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n904), .B(KEYINPUT49), .ZN(new_n926));
  NOR4_X1   g740(.A1(new_n807), .A2(new_n267), .A3(new_n471), .A4(new_n517), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT112), .Z(new_n928));
  OR3_X1    g742(.A1(new_n928), .A2(new_n728), .A3(new_n731), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n925), .B1(new_n926), .B2(new_n929), .ZN(G75));
  OAI21_X1  g744(.A(KEYINPUT116), .B1(new_n864), .B2(new_n865), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n879), .A2(new_n880), .A3(new_n863), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT53), .B1(new_n933), .B2(new_n859), .ZN(new_n934));
  INV_X1    g748(.A(new_n888), .ZN(new_n935));
  OAI211_X1 g749(.A(G210), .B(G902), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT56), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(KEYINPUT121), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n188), .A2(G952), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n495), .B(new_n501), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT55), .Z(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n255), .B1(new_n886), .B2(new_n888), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT56), .B1(new_n945), .B2(G210), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n946), .B2(KEYINPUT121), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n936), .A2(new_n937), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT121), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(new_n949), .A3(new_n943), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n941), .B1(new_n947), .B2(new_n950), .ZN(G51));
  XNOR2_X1  g765(.A(new_n816), .B(KEYINPUT57), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n465), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n945), .A2(new_n814), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n939), .B1(new_n956), .B2(new_n957), .ZN(G54));
  NAND2_X1  g772(.A1(KEYINPUT58), .A2(G475), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n945), .A2(new_n581), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n581), .B1(new_n945), .B2(new_n960), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n939), .ZN(G60));
  XOR2_X1   g777(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n964));
  NOR2_X1   g778(.A1(new_n637), .A2(new_n255), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  AOI22_X1  g781(.A1(new_n890), .A2(new_n967), .B1(new_n669), .B2(new_n670), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n669), .A2(new_n670), .A3(new_n967), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n953), .B2(new_n954), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n940), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n968), .A2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n886), .B2(new_n888), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n975), .A2(new_n264), .ZN(new_n976));
  INV_X1    g790(.A(new_n974), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n699), .B(new_n977), .C1(new_n934), .C2(new_n935), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n976), .A2(KEYINPUT61), .A3(new_n940), .A4(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n978), .B(new_n940), .C1(new_n264), .C2(new_n975), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n979), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n647), .B2(new_n499), .ZN(new_n984));
  INV_X1    g798(.A(new_n854), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(G953), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n522), .B(new_n489), .C1(G898), .C2(new_n188), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT123), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT124), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n986), .B(new_n989), .ZN(G69));
  OAI211_X1 g804(.A(new_n387), .B(new_n788), .C1(new_n847), .C2(new_n838), .ZN(new_n991));
  OAI221_X1 g805(.A(new_n823), .B1(new_n721), .B2(new_n991), .C1(new_n831), .C2(new_n832), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n877), .A2(new_n739), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n735), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n339), .A2(new_n321), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT125), .Z(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(new_n573), .Z(new_n1000));
  NOR3_X1   g814(.A1(new_n997), .A2(G953), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n822), .A2(new_n772), .A3(new_n787), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n823), .A2(new_n1003), .A3(new_n805), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1004), .A2(new_n801), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1005), .A2(new_n833), .A3(new_n188), .A4(new_n993), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G900), .A2(G953), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1002), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n1001), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G227), .A2(G900), .ZN(new_n1012));
  AND4_X1   g826(.A1(G953), .A2(new_n1011), .A3(new_n1012), .A4(new_n1000), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1010), .A2(new_n1013), .ZN(G72));
  INV_X1    g828(.A(new_n378), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1015), .A2(new_n724), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  XOR2_X1   g831(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1018));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT127), .Z(new_n1021));
  AOI21_X1  g835(.A(new_n939), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n1005), .A2(new_n833), .A3(new_n993), .ZN(new_n1023));
  AOI22_X1  g837(.A1(new_n997), .A2(new_n724), .B1(new_n1023), .B2(new_n1015), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1022), .B1(new_n1024), .B2(new_n854), .ZN(new_n1025));
  AND3_X1   g839(.A1(new_n884), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1025), .A2(new_n1026), .ZN(G57));
endmodule


