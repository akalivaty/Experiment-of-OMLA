//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT86), .Z(new_n188));
  INV_X1    g002(.A(KEYINPUT85), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G122), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT8), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n196), .A3(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n193), .A2(G119), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(KEYINPUT5), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G113), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT5), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n198), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G116), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n198), .B1(new_n205), .B2(G119), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT2), .B(G113), .Z(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT75), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(KEYINPUT75), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n210), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT76), .A2(G101), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT76), .A2(G101), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G107), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT75), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n218), .A2(G107), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n214), .A2(new_n217), .A3(new_n219), .A4(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n213), .A2(new_n219), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G101), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n204), .A2(new_n208), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n204), .A2(new_n208), .B1(new_n224), .B2(new_n226), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n192), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT1), .B1(new_n235), .B2(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT64), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n241), .B(KEYINPUT1), .C1(new_n235), .C2(G146), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(G128), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n234), .A2(new_n236), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n238), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT70), .B(G125), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OR2_X1    g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n244), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G143), .B(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n249), .ZN(new_n253));
  INV_X1    g067(.A(new_n246), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G224), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(KEYINPUT83), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT7), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT84), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n247), .A2(KEYINPUT7), .A3(new_n255), .A4(new_n259), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n230), .A2(new_n261), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n197), .A2(new_n199), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(new_n207), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n221), .B1(new_n222), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n219), .B1(new_n210), .B2(new_n213), .ZN(new_n270));
  OAI21_X1  g084(.A(G101), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n271), .B2(new_n224), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n267), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n227), .A3(new_n191), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n264), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n204), .A2(new_n208), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n224), .A2(new_n226), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n227), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n281), .A2(new_n192), .B1(new_n256), .B2(new_n260), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n262), .B1(new_n282), .B2(new_n263), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n189), .B(new_n190), .C1(new_n277), .C2(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n256), .B(new_n259), .Z(new_n285));
  NAND2_X1  g099(.A1(new_n275), .A2(new_n227), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n191), .B(KEYINPUT82), .Z(new_n287));
  AOI22_X1  g101(.A1(new_n276), .A2(KEYINPUT6), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n286), .A2(KEYINPUT6), .A3(new_n287), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n230), .A2(new_n261), .A3(new_n263), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT84), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n276), .A3(new_n264), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n189), .B1(new_n294), .B2(new_n190), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n188), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n190), .B1(new_n277), .B2(new_n283), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT85), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n298), .A2(new_n187), .A3(new_n290), .A4(new_n284), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT87), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT87), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n304), .A3(new_n301), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n231), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n237), .B1(new_n307), .B2(new_n252), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n224), .A2(new_n226), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n224), .A2(new_n308), .A3(KEYINPUT77), .A4(new_n226), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n245), .A2(new_n279), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT11), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G137), .ZN(new_n318));
  INV_X1    g132(.A(G137), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT11), .A3(G134), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(G137), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  INV_X1    g137(.A(G131), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n318), .A2(new_n320), .A3(new_n324), .A4(new_n321), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n315), .A2(KEYINPUT12), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT12), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n311), .A2(new_n312), .B1(new_n245), .B2(new_n279), .ZN(new_n329));
  INV_X1    g143(.A(new_n326), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n327), .A2(new_n331), .A3(KEYINPUT79), .ZN(new_n332));
  XNOR2_X1  g146(.A(G110), .B(G140), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n257), .A2(G227), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT10), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n313), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n224), .A2(new_n226), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n242), .A2(G128), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n241), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n244), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n237), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT10), .A4(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n224), .A2(KEYINPUT10), .A3(new_n226), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT78), .B1(new_n346), .B2(new_n245), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n234), .A2(new_n236), .B1(new_n248), .B2(new_n249), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n234), .A2(new_n236), .A3(new_n249), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT66), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT66), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n251), .A2(new_n352), .A3(new_n253), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n351), .B(new_n353), .C1(new_n273), .C2(new_n274), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n338), .A2(new_n348), .A3(new_n330), .A4(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n356), .B(new_n328), .C1(new_n329), .C2(new_n330), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n332), .A2(new_n336), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n355), .A2(new_n357), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n361), .A2(KEYINPUT81), .A3(new_n336), .A4(new_n332), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n338), .A2(new_n348), .A3(new_n354), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n326), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n355), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n335), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n360), .A2(new_n362), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G469), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT68), .B(G902), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n327), .A2(new_n331), .A3(KEYINPUT79), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n355), .A2(new_n357), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT80), .B1(new_n361), .B2(new_n332), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n335), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n365), .A2(new_n366), .A3(new_n335), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(G469), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(G469), .A2(G902), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n371), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT9), .B(G234), .ZN(new_n383));
  OAI21_X1  g197(.A(G221), .B1(new_n383), .B2(G902), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G217), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n370), .B2(G234), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT22), .B(G137), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n390), .B(new_n391), .Z(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT16), .ZN(new_n394));
  INV_X1    g208(.A(G125), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n395), .A2(KEYINPUT70), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(KEYINPUT70), .ZN(new_n397));
  OAI21_X1  g211(.A(G140), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n394), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n394), .A2(new_n399), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n246), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n233), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n400), .B1(new_n246), .B2(new_n399), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n405), .B2(KEYINPUT16), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G146), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n407), .A3(KEYINPUT71), .ZN(new_n408));
  OR3_X1    g222(.A1(new_n406), .A2(KEYINPUT71), .A3(G146), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT69), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n231), .A2(G119), .ZN(new_n411));
  INV_X1    g225(.A(G119), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(G128), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n410), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(G128), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n231), .A2(G119), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT69), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(KEYINPUT24), .B(G110), .Z(new_n419));
  NAND3_X1  g233(.A1(new_n231), .A2(KEYINPUT23), .A3(G119), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n415), .B(new_n420), .C1(new_n413), .C2(KEYINPUT23), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n418), .A2(new_n419), .B1(G110), .B2(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n408), .A2(new_n409), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT73), .ZN(new_n424));
  XNOR2_X1  g238(.A(G125), .B(G140), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n233), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT72), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT72), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n428), .A3(new_n233), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n419), .B1(new_n414), .B2(new_n417), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n421), .A2(G110), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n401), .A2(new_n233), .A3(new_n403), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n424), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n431), .A2(new_n432), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(new_n407), .A3(KEYINPUT73), .A4(new_n430), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n393), .B1(new_n423), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n408), .A2(new_n409), .A3(new_n422), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n440), .A2(new_n435), .A3(new_n437), .A4(new_n392), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n370), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT25), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n439), .A2(KEYINPUT25), .A3(new_n370), .A4(new_n441), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n389), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n439), .A2(new_n441), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n388), .A2(G902), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT74), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT74), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n446), .B2(new_n450), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n317), .A2(G137), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n319), .A2(G134), .ZN(new_n457));
  OAI21_X1  g271(.A(G131), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n344), .A2(new_n325), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n326), .A2(new_n351), .A3(new_n353), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(KEYINPUT30), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n325), .A2(new_n458), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n343), .B2(new_n237), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n323), .A2(new_n325), .B1(new_n251), .B2(new_n253), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n461), .A2(new_n267), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n459), .A2(new_n266), .A3(new_n460), .ZN(new_n468));
  INV_X1    g282(.A(G237), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n257), .A3(G210), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT27), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT26), .B(G101), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n467), .A2(new_n468), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT31), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT31), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n467), .A2(new_n476), .A3(new_n468), .A4(new_n473), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n468), .A2(KEYINPUT28), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT28), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n459), .A2(new_n479), .A3(new_n460), .A4(new_n266), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n464), .A2(new_n465), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n478), .A2(new_n480), .B1(new_n267), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n475), .B(new_n477), .C1(new_n482), .C2(new_n473), .ZN(new_n483));
  NOR2_X1   g297(.A1(G472), .A2(G902), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(KEYINPUT32), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n459), .A2(new_n460), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n478), .A2(new_n480), .B1(new_n486), .B2(new_n267), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n473), .A2(KEYINPUT29), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n370), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT29), .ZN(new_n492));
  INV_X1    g306(.A(new_n473), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n467), .A2(new_n468), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n482), .B2(new_n493), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n491), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G472), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n485), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n483), .A2(new_n499), .A3(new_n484), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n483), .B2(new_n484), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT32), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n455), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n469), .A2(new_n257), .A3(G214), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n235), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(new_n324), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n408), .A2(new_n409), .B1(KEYINPUT17), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n512), .A2(KEYINPUT91), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(KEYINPUT89), .A3(new_n324), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT89), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n509), .B2(G131), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n514), .B(new_n516), .C1(new_n324), .C2(new_n510), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(KEYINPUT17), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n512), .B2(KEYINPUT91), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(G113), .B(G122), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(new_n218), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n398), .A2(G146), .A3(new_n400), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n524), .A2(KEYINPUT88), .B1(new_n429), .B2(new_n427), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(KEYINPUT88), .B2(new_n524), .ZN(new_n526));
  NAND2_X1  g340(.A1(KEYINPUT18), .A2(G131), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n509), .B(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n520), .A2(new_n522), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT19), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n425), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n405), .B2(new_n531), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G146), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n534), .B(KEYINPUT90), .Z(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n407), .A3(new_n517), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n529), .ZN(new_n537));
  INV_X1    g351(.A(new_n522), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(G475), .A2(G902), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n507), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n541), .ZN(new_n543));
  AOI211_X1 g357(.A(KEYINPUT20), .B(new_n543), .C1(new_n530), .C2(new_n539), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n520), .A2(new_n529), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n538), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n546), .B2(new_n530), .ZN(new_n547));
  INV_X1    g361(.A(G475), .ZN(new_n548));
  OAI22_X1  g362(.A1(new_n542), .A2(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G952), .ZN(new_n550));
  AOI211_X1 g364(.A(G953), .B(new_n550), .C1(G234), .C2(G237), .ZN(new_n551));
  AOI211_X1 g365(.A(new_n257), .B(new_n370), .C1(G234), .C2(G237), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT21), .B(G898), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n370), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT92), .B1(new_n231), .B2(G143), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(new_n235), .A3(G128), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n235), .A2(G128), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n317), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n194), .A2(new_n196), .A3(G122), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n193), .A2(G122), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n212), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n212), .B1(new_n563), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n562), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT13), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n559), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(KEYINPUT93), .A3(new_n561), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT13), .B1(new_n556), .B2(new_n558), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n572), .B1(new_n573), .B2(new_n560), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n571), .B(new_n574), .C1(new_n569), .C2(new_n559), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n568), .B1(new_n575), .B2(G134), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT14), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n194), .A2(new_n196), .A3(new_n578), .A4(G122), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n579), .A2(new_n564), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n563), .A2(new_n581), .A3(KEYINPUT14), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n563), .B2(KEYINPUT14), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n566), .B1(new_n584), .B2(G107), .ZN(new_n585));
  AOI211_X1 g399(.A(G134), .B(new_n560), .C1(new_n558), .C2(new_n556), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n317), .B1(new_n559), .B2(new_n561), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT94), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n557), .B1(G128), .B2(new_n235), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n231), .A2(KEYINPUT92), .A3(G143), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n561), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G134), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n562), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n585), .A2(KEYINPUT96), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT96), .B1(new_n585), .B2(new_n595), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n577), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n383), .A2(new_n387), .A3(G953), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n579), .A2(new_n564), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n563), .A2(KEYINPUT14), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT95), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n563), .A2(new_n581), .A3(KEYINPUT14), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n565), .B1(new_n607), .B2(new_n212), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n588), .A2(new_n594), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n602), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n585), .A2(KEYINPUT96), .A3(new_n595), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n577), .A3(new_n599), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n555), .B1(new_n601), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT97), .ZN(new_n615));
  INV_X1    g429(.A(G478), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(KEYINPUT15), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n615), .B(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n549), .A2(new_n554), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n306), .A2(new_n386), .A3(new_n506), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT98), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(new_n217), .ZN(G3));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n614), .B2(G478), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n600), .B2(KEYINPUT99), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n599), .B1(new_n612), .B2(new_n577), .ZN(new_n628));
  AOI211_X1 g442(.A(new_n576), .B(new_n600), .C1(new_n610), .C2(new_n611), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n601), .A2(new_n613), .A3(new_n626), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n555), .A2(new_n616), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n630), .A2(new_n623), .A3(new_n631), .A4(new_n632), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT101), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n634), .A2(new_n638), .A3(new_n635), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n637), .A2(new_n549), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n301), .ZN(new_n641));
  INV_X1    g455(.A(new_n187), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n291), .B2(new_n295), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n641), .B1(new_n643), .B2(new_n299), .ZN(new_n644));
  INV_X1    g458(.A(new_n554), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n483), .A2(new_n370), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(G472), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n452), .A2(new_n503), .A3(new_n454), .A4(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n385), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  AOI21_X1  g468(.A(new_n522), .B1(new_n536), .B2(new_n529), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n513), .A2(new_n519), .B1(new_n526), .B2(new_n528), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n655), .B1(new_n656), .B2(new_n522), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT20), .B1(new_n657), .B2(new_n543), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n540), .A2(new_n507), .A3(new_n541), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n530), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n656), .A2(new_n522), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n190), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G475), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n618), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n646), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n651), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  NAND2_X1  g483(.A1(new_n444), .A2(new_n445), .ZN(new_n670));
  INV_X1    g484(.A(new_n438), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n440), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n393), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n670), .A2(new_n388), .B1(new_n674), .B2(new_n448), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n503), .A3(KEYINPUT102), .A4(new_n649), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n483), .A2(new_n484), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT67), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n649), .A2(new_n680), .A3(new_n500), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n678), .B1(new_n681), .B2(new_n675), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n306), .A3(new_n386), .A4(new_n619), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT37), .B(G110), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  NAND3_X1  g500(.A1(new_n680), .A2(new_n504), .A3(new_n500), .ZN(new_n687));
  INV_X1    g501(.A(new_n484), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n475), .A2(new_n477), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n482), .A2(new_n473), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n495), .A2(new_n492), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n555), .B1(new_n487), .B2(new_n489), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n691), .A2(KEYINPUT32), .B1(new_n694), .B2(G472), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n675), .B1(new_n687), .B2(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n696), .A2(new_n384), .A3(new_n382), .ZN(new_n697));
  INV_X1    g511(.A(G900), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n552), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(KEYINPUT103), .ZN(new_n700));
  INV_X1    g514(.A(new_n551), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(KEYINPUT103), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n665), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n697), .A2(new_n644), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT104), .B(G128), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G30));
  XNOR2_X1  g522(.A(new_n703), .B(KEYINPUT39), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n386), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n300), .B(KEYINPUT38), .Z(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n676), .A2(new_n641), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n486), .A2(new_n267), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n468), .A3(new_n493), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n190), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n493), .B1(new_n467), .B2(new_n468), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n485), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n687), .A2(new_n721), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n618), .A2(new_n715), .A3(new_n549), .A4(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n711), .A2(new_n712), .A3(new_n714), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT105), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G143), .ZN(G45));
  AND4_X1   g540(.A1(new_n384), .A2(new_n696), .A3(new_n382), .A4(new_n644), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n637), .A2(new_n549), .A3(new_n639), .A4(new_n703), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n368), .A2(new_n370), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G469), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n371), .ZN(new_n735));
  INV_X1    g549(.A(new_n384), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n734), .A2(KEYINPUT106), .A3(new_n384), .A4(new_n371), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n647), .A2(new_n506), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND4_X1  g555(.A1(new_n737), .A2(new_n666), .A3(new_n506), .A4(new_n738), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G116), .ZN(G18));
  AND4_X1   g557(.A1(new_n384), .A2(new_n644), .A3(new_n734), .A4(new_n371), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n619), .A3(new_n696), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  OAI21_X1  g560(.A(new_n689), .B1(new_n473), .B2(new_n487), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n747), .A2(new_n484), .B1(new_n648), .B2(G472), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(new_n451), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(new_n645), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n549), .A2(new_n618), .A3(new_n644), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n737), .A2(new_n750), .A3(new_n751), .A4(new_n738), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  AOI22_X1  g567(.A1(new_n659), .A2(new_n658), .B1(new_n663), .B2(G475), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n634), .A2(new_n638), .A3(new_n635), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n638), .B1(new_n634), .B2(new_n635), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n676), .A2(new_n748), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n744), .A3(new_n703), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  NOR2_X1   g575(.A1(new_n728), .A2(KEYINPUT42), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n382), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n373), .B1(new_n372), .B2(new_n374), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n361), .A2(KEYINPUT80), .A3(new_n332), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n378), .B1(new_n767), .B2(new_n335), .ZN(new_n768));
  OAI21_X1  g582(.A(G469), .B1(new_n768), .B2(G902), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(KEYINPUT107), .A3(new_n371), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n300), .A2(new_n641), .A3(new_n736), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n764), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n762), .A2(new_n772), .A3(new_n506), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n755), .A2(new_n756), .ZN(new_n774));
  INV_X1    g588(.A(new_n451), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT108), .B1(new_n679), .B2(new_n504), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n498), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n679), .A2(KEYINPUT108), .A3(new_n504), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n774), .A2(new_n779), .A3(new_n549), .A4(new_n703), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n764), .A2(new_n770), .A3(new_n771), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT42), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n773), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n783), .B1(new_n773), .B2(new_n782), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G131), .ZN(G33));
  AOI21_X1  g601(.A(KEYINPUT107), .B1(new_n769), .B2(new_n371), .ZN(new_n788));
  AND4_X1   g602(.A1(KEYINPUT107), .A2(new_n371), .A3(new_n380), .A4(new_n381), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n506), .A3(new_n705), .A4(new_n771), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  NOR2_X1   g606(.A1(new_n300), .A2(new_n641), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n774), .A2(new_n754), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT43), .Z(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n681), .A3(new_n676), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT44), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n768), .A2(KEYINPUT45), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n768), .A2(KEYINPUT45), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(G469), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n381), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(KEYINPUT46), .A3(new_n381), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n371), .A3(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(new_n384), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(new_n709), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n799), .B(new_n809), .C1(new_n798), .C2(new_n797), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G137), .ZN(G39));
  NAND2_X1  g625(.A1(new_n808), .A2(KEYINPUT47), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n807), .A2(new_n384), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n455), .A2(new_n505), .A3(new_n793), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n729), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  NAND3_X1  g633(.A1(new_n451), .A2(new_n301), .A3(new_n384), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n714), .A2(new_n722), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n795), .B1(KEYINPUT49), .B2(new_n735), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n821), .B(new_n822), .C1(KEYINPUT49), .C2(new_n735), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n739), .A2(new_n620), .A3(new_n742), .A4(new_n745), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n728), .A2(new_n758), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n772), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n549), .A2(new_n618), .A3(new_n704), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n697), .A2(new_n793), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n791), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n640), .A2(new_n665), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n554), .B1(new_n303), .B2(new_n305), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n651), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n684), .A3(new_n752), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n825), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n727), .B1(new_n729), .B2(new_n705), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n675), .A2(new_n384), .A3(new_n703), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n687), .B2(new_n721), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n751), .A2(new_n838), .A3(new_n764), .A4(new_n770), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n836), .A2(new_n760), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n836), .A2(KEYINPUT52), .A3(new_n760), .A4(new_n839), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n773), .A2(new_n782), .A3(KEYINPUT53), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n835), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n786), .A2(new_n835), .A3(new_n844), .ZN(new_n847));
  XOR2_X1   g661(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n848));
  AND3_X1   g662(.A1(new_n847), .A2(KEYINPUT111), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT111), .B1(new_n847), .B2(new_n848), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n824), .B(new_n846), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n786), .A2(new_n835), .A3(new_n844), .A4(new_n848), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(KEYINPUT54), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT112), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n851), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n735), .A2(new_n736), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n796), .A2(new_n551), .A3(new_n860), .A4(new_n793), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n758), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n793), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n863), .A2(new_n455), .A3(new_n701), .A4(new_n722), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n774), .A2(new_n549), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n796), .A2(new_n551), .A3(new_n749), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n713), .A2(new_n641), .A3(new_n860), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT113), .ZN(new_n870));
  NOR2_X1   g684(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n812), .A2(new_n815), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n734), .A2(new_n736), .A3(new_n371), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n868), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n793), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(KEYINPUT114), .B(KEYINPUT50), .C1(new_n868), .C2(new_n870), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n875), .A2(new_n880), .A3(KEYINPUT51), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n779), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n861), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT48), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n879), .A2(new_n744), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n550), .B(G953), .C1(new_n864), .C2(new_n757), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n794), .B(new_n868), .C1(new_n876), .C2(new_n877), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n867), .A2(new_n874), .A3(new_n881), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT115), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(KEYINPUT115), .B(new_n891), .C1(new_n892), .C2(new_n893), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n890), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n859), .A2(new_n898), .A3(KEYINPUT116), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(G952), .B2(G953), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT116), .B1(new_n859), .B2(new_n898), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n823), .B1(new_n900), .B2(new_n901), .ZN(G75));
  NOR2_X1   g716(.A1(new_n257), .A2(G952), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n288), .A2(new_n289), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n285), .ZN(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n370), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n642), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n910), .A2(new_n188), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n907), .A2(new_n912), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n903), .B(new_n913), .C1(new_n914), .C2(new_n915), .ZN(G51));
  NOR3_X1   g730(.A1(new_n909), .A2(new_n370), .A3(new_n802), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT119), .Z(new_n918));
  XNOR2_X1  g732(.A(new_n368), .B(KEYINPUT118), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n851), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n381), .B(KEYINPUT57), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n903), .B1(new_n918), .B2(new_n924), .ZN(G54));
  NAND3_X1  g739(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n926), .A2(KEYINPUT120), .A3(new_n657), .ZN(new_n927));
  INV_X1    g741(.A(new_n903), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n926), .B2(new_n657), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT120), .B1(new_n926), .B2(new_n657), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(G60));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n630), .A2(new_n631), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT59), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n933), .B1(new_n921), .B2(new_n939), .ZN(new_n940));
  AOI211_X1 g754(.A(KEYINPUT121), .B(new_n938), .C1(new_n920), .C2(new_n851), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n928), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n851), .A2(new_n854), .A3(new_n857), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n857), .B1(new_n851), .B2(new_n854), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n935), .B1(new_n945), .B2(new_n937), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n932), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n847), .A2(new_n848), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT111), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n847), .A2(KEYINPUT111), .A3(new_n848), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n824), .B1(new_n952), .B2(new_n846), .ZN(new_n953));
  INV_X1    g767(.A(new_n851), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n939), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT121), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n921), .A2(new_n933), .A3(new_n939), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n856), .A2(new_n858), .A3(new_n937), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n934), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n958), .A2(new_n960), .A3(KEYINPUT122), .A4(new_n928), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n947), .A2(new_n961), .ZN(G63));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT60), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n908), .A2(new_n674), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n909), .A2(new_n964), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n928), .B(new_n966), .C1(new_n967), .C2(new_n447), .ZN(new_n968));
  XNOR2_X1  g782(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n968), .A2(KEYINPUT124), .A3(new_n969), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n972), .B(new_n973), .C1(new_n974), .C2(new_n968), .ZN(G66));
  INV_X1    g789(.A(G224), .ZN(new_n976));
  OAI21_X1  g790(.A(G953), .B1(new_n553), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n825), .A2(new_n834), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n904), .B1(G898), .B2(new_n257), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G69));
  NAND2_X1  g795(.A1(new_n810), .A2(new_n818), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n809), .A2(new_n751), .A3(new_n779), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n983), .A2(new_n760), .A3(new_n791), .A4(new_n836), .ZN(new_n984));
  INV_X1    g798(.A(new_n786), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n257), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n461), .A2(new_n466), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT125), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(new_n533), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(G900), .B2(G953), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n257), .B1(G227), .B2(G900), .ZN(new_n992));
  AOI22_X1  g806(.A1(new_n987), .A2(new_n991), .B1(KEYINPUT127), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n725), .A2(new_n760), .A3(new_n836), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT62), .ZN(new_n995));
  INV_X1    g809(.A(new_n831), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n996), .A2(KEYINPUT126), .ZN(new_n997));
  NOR4_X1   g811(.A1(new_n710), .A2(new_n505), .A3(new_n455), .A4(new_n794), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(new_n831), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n810), .B(new_n818), .C1(new_n997), .C2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n257), .B1(new_n995), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n990), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n993), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n992), .A2(KEYINPUT127), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1004), .B(new_n1005), .Z(G72));
  NOR4_X1   g820(.A1(new_n995), .A2(new_n1001), .A3(new_n834), .A4(new_n825), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT63), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n719), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n494), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n986), .A2(new_n978), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1011), .B1(new_n1012), .B2(new_n1009), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1011), .A2(new_n719), .A3(new_n1009), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n852), .A2(new_n853), .A3(new_n1014), .ZN(new_n1015));
  AND4_X1   g829(.A1(new_n928), .A2(new_n1010), .A3(new_n1013), .A4(new_n1015), .ZN(G57));
endmodule


