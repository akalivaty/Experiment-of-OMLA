//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1224, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0007(.A1(G97), .A2(G107), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  NAND2_X1  g0018(.A1(new_n206), .A2(G50), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n212), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n229));
  AND3_X1   g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n213), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n223), .B1(new_n224), .B2(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n218), .B(new_n232), .C1(new_n224), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G222), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G223), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n257), .B1(new_n258), .B2(new_n255), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT70), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT70), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n266), .B(new_n211), .C1(G41), .C2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  OAI211_X1 g0068(.A(G1), .B(G13), .C1(new_n252), .C2(new_n268), .ZN(new_n269));
  AND3_X1   g0069(.A1(new_n265), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n264), .A2(KEYINPUT69), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n274), .B(new_n211), .C1(G41), .C2(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n270), .A2(G226), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n263), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT71), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n263), .A2(KEYINPUT71), .A3(new_n277), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G179), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n212), .A2(G33), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n285), .B1(new_n286), .B2(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n221), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n293), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n211), .A2(G20), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G50), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n298), .A2(new_n300), .B1(G50), .B2(new_n295), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n280), .A2(new_n304), .A3(new_n281), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n284), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n282), .A2(G190), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT9), .B1(new_n294), .B2(new_n302), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  AOI211_X1 g0109(.A(new_n309), .B(new_n301), .C1(new_n291), .C2(new_n293), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n280), .A2(G200), .A3(new_n281), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n307), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n312), .B2(KEYINPUT72), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n313), .A2(new_n315), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n306), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n289), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n299), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n298), .A2(new_n320), .B1(new_n295), .B2(new_n319), .ZN(new_n321));
  INV_X1    g0121(.A(new_n293), .ZN(new_n322));
  AND2_X1   g0122(.A1(KEYINPUT3), .A2(G33), .ZN(new_n323));
  NOR2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT7), .B1(new_n325), .B2(new_n212), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n253), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n254), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(G68), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT75), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n253), .A2(new_n212), .A3(new_n254), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT7), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n327), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(KEYINPUT75), .A3(G68), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT16), .ZN(new_n338));
  INV_X1    g0138(.A(G159), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n288), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n341));
  AOI211_X1 g0141(.A(new_n338), .B(new_n340), .C1(new_n341), .C2(G20), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n322), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT76), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n334), .A2(new_n344), .A3(new_n327), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n328), .A2(KEYINPUT76), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(G68), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n340), .B1(new_n341), .B2(G20), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n338), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n321), .B1(new_n343), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G226), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G1698), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G223), .B2(G1698), .ZN(new_n354));
  INV_X1    g0154(.A(G87), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n354), .A2(new_n325), .B1(new_n252), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n262), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n265), .A2(G232), .A3(new_n269), .A4(new_n267), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n272), .A2(new_n276), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n283), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n356), .A2(new_n262), .B1(new_n272), .B2(new_n276), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n304), .B1(new_n362), .B2(new_n358), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT18), .B1(new_n351), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT18), .ZN(new_n366));
  INV_X1    g0166(.A(new_n364), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n348), .A2(KEYINPUT16), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n331), .B2(new_n336), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT16), .B1(new_n347), .B2(new_n348), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n369), .A2(new_n370), .A3(new_n322), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n366), .B(new_n367), .C1(new_n371), .C2(new_n321), .ZN(new_n372));
  INV_X1    g0172(.A(G200), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n360), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(G190), .B2(new_n360), .ZN(new_n375));
  INV_X1    g0175(.A(new_n321), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT75), .B1(new_n335), .B2(G68), .ZN(new_n377));
  AOI211_X1 g0177(.A(new_n330), .B(new_n203), .C1(new_n334), .C2(new_n327), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n342), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n293), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n375), .B(new_n376), .C1(new_n380), .C2(new_n370), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT17), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n350), .A2(new_n293), .A3(new_n379), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n384), .A2(KEYINPUT17), .A3(new_n376), .A4(new_n375), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n365), .A2(new_n372), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n212), .A2(G33), .A3(G77), .ZN(new_n387));
  INV_X1    g0187(.A(G50), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n387), .B1(new_n212), .B2(G68), .C1(new_n288), .C2(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n389), .A2(KEYINPUT11), .A3(new_n293), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT11), .B1(new_n389), .B2(new_n293), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n322), .A2(G68), .A3(new_n295), .A4(new_n299), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT74), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n211), .A2(new_n203), .A3(G13), .A4(G20), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT73), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT12), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT12), .B1(new_n395), .B2(new_n396), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n393), .B(new_n394), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n393), .B1(new_n397), .B2(new_n398), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT74), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n392), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT14), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n352), .A2(new_n256), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(G232), .B2(new_n256), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n407), .B2(new_n325), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n262), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n265), .A2(G238), .A3(new_n269), .A4(new_n267), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n359), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(KEYINPUT13), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n408), .A2(new_n262), .B1(new_n272), .B2(new_n276), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(new_n410), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n404), .B(G169), .C1(new_n412), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(KEYINPUT13), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n413), .A3(new_n410), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(G179), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(new_n418), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n404), .B1(new_n421), .B2(G169), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n403), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n417), .A2(G190), .A3(new_n418), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n402), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n373), .B1(new_n417), .B2(new_n418), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n297), .A2(G77), .A3(new_n299), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G77), .B2(new_n295), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n319), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n431), .B1(new_n290), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n430), .B1(new_n433), .B2(new_n293), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n255), .A2(G232), .A3(new_n256), .ZN(new_n435));
  INV_X1    g0235(.A(G107), .ZN(new_n436));
  INV_X1    g0236(.A(G238), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n435), .B1(new_n436), .B2(new_n255), .C1(new_n259), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n262), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n270), .A2(G244), .B1(new_n272), .B2(new_n276), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G190), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n434), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n373), .B1(new_n439), .B2(new_n440), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n434), .B1(new_n441), .B2(new_n304), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n439), .A2(new_n283), .A3(new_n440), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n423), .A2(new_n428), .A3(new_n445), .A4(new_n448), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n318), .A2(new_n386), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(G257), .B(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n452));
  OAI211_X1 g0252(.A(G250), .B(new_n256), .C1(new_n323), .C2(new_n324), .ZN(new_n453));
  INV_X1    g0253(.A(G294), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n452), .B(new_n453), .C1(new_n252), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n211), .A2(G45), .ZN(new_n456));
  OR2_X1    g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  NAND2_X1  g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n262), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n455), .A2(new_n262), .B1(new_n460), .B2(G264), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n272), .A2(new_n459), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n283), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n455), .A2(new_n262), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(G264), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n304), .ZN(new_n467));
  INV_X1    g0267(.A(G116), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n290), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT82), .B1(new_n212), .B2(G107), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT23), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT23), .ZN(new_n472));
  OAI211_X1 g0272(.A(KEYINPUT82), .B(new_n472), .C1(new_n212), .C2(G107), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n469), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n212), .B(G87), .C1(new_n323), .C2(new_n324), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n475), .A2(KEYINPUT22), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(KEYINPUT22), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT24), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n475), .B(KEYINPUT22), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT24), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(new_n474), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n322), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n252), .A2(G1), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n296), .A2(new_n293), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT25), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n295), .A2(new_n486), .A3(G107), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n295), .B2(G107), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n485), .A2(G107), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n463), .B(new_n467), .C1(new_n483), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n466), .A2(new_n373), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n461), .A2(new_n442), .A3(new_n462), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n478), .A2(KEYINPUT24), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n481), .B1(new_n480), .B2(new_n474), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n293), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n498), .A3(new_n490), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n456), .A2(G250), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT80), .B1(new_n262), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT80), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n269), .A2(new_n502), .A3(G250), .A4(new_n456), .ZN(new_n503));
  INV_X1    g0303(.A(new_n456), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n501), .A2(new_n503), .B1(new_n272), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n506));
  OAI211_X1 g0306(.A(G238), .B(new_n256), .C1(new_n323), .C2(new_n324), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(new_n507), .C1(new_n252), .C2(new_n468), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n262), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n505), .A2(new_n509), .A3(G190), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n373), .B1(new_n505), .B2(new_n509), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n255), .A2(new_n212), .A3(G68), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT19), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n212), .B1(new_n405), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G87), .B2(new_n209), .ZN(new_n516));
  INV_X1    g0316(.A(G97), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n514), .B1(new_n290), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n513), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n293), .B1(new_n296), .B2(new_n432), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n485), .A2(G87), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n512), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n505), .A2(new_n509), .ZN(new_n524));
  INV_X1    g0324(.A(new_n432), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n485), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n304), .A2(new_n524), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n505), .A2(new_n509), .A3(KEYINPUT81), .A4(new_n283), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT81), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n524), .B2(G179), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n492), .A2(new_n499), .A3(new_n523), .A4(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n295), .A2(G97), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n485), .B2(G97), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n345), .A2(G107), .A3(new_n346), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT77), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n288), .A2(new_n258), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  AND2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n540), .B2(new_n208), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n436), .A2(KEYINPUT6), .A3(G97), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n536), .B(new_n538), .C1(new_n543), .C2(new_n212), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n212), .B1(new_n541), .B2(new_n542), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT77), .B1(new_n545), .B2(new_n537), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n535), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT78), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n547), .A2(new_n548), .A3(new_n293), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n547), .B2(new_n293), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n534), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(G244), .B(new_n256), .C1(new_n323), .C2(new_n324), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT79), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT4), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n255), .A2(G244), .A3(new_n256), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G283), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n255), .A2(G250), .A3(G1698), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n555), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n262), .ZN(new_n561));
  XNOR2_X1  g0361(.A(KEYINPUT5), .B(G41), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n504), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(G257), .A3(new_n269), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n462), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n304), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n565), .B1(new_n262), .B2(new_n560), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n283), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n551), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n561), .A2(new_n442), .A3(new_n566), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(G200), .B2(new_n569), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n575), .B(new_n534), .C1(new_n549), .C2(new_n550), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n460), .A2(G270), .B1(new_n272), .B2(new_n459), .ZN(new_n577));
  OAI211_X1 g0377(.A(G264), .B(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n578));
  OAI211_X1 g0378(.A(G257), .B(new_n256), .C1(new_n323), .C2(new_n324), .ZN(new_n579));
  INV_X1    g0379(.A(G303), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n255), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n262), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n292), .A2(new_n221), .B1(G20), .B2(new_n468), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n558), .B(new_n212), .C1(G33), .C2(new_n517), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT20), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(KEYINPUT20), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n296), .A2(new_n468), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n485), .A2(G116), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n583), .A2(new_n593), .A3(G169), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n583), .A2(G200), .ZN(new_n597));
  INV_X1    g0397(.A(new_n593), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n577), .A2(G190), .A3(new_n582), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n577), .A2(G179), .A3(new_n582), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n593), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n583), .A2(new_n593), .A3(KEYINPUT21), .A4(G169), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n596), .A2(new_n600), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n532), .A2(new_n573), .A3(new_n576), .A4(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n451), .A2(new_n606), .ZN(G372));
  INV_X1    g0407(.A(new_n306), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n365), .A2(new_n372), .ZN(new_n609));
  INV_X1    g0409(.A(new_n448), .ZN(new_n610));
  OAI21_X1  g0410(.A(G169), .B1(new_n412), .B2(new_n415), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT14), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n419), .A3(new_n416), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n428), .A2(new_n610), .B1(new_n613), .B2(new_n403), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n383), .A2(new_n385), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n609), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n315), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(new_n312), .A3(new_n307), .A4(new_n311), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n313), .A2(new_n315), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n608), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n505), .A2(new_n509), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n283), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n527), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n522), .A2(new_n512), .B1(new_n527), .B2(new_n623), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n483), .A2(new_n491), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n467), .A2(new_n463), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n596), .A2(new_n602), .A3(new_n603), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n499), .B(new_n625), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n534), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n547), .A2(new_n293), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT78), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n547), .A2(new_n548), .A3(new_n293), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n576), .B1(new_n635), .B2(new_n571), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n624), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n551), .A2(new_n625), .A3(new_n572), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n531), .A2(new_n523), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(KEYINPUT26), .A3(new_n551), .A4(new_n572), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n621), .B1(new_n451), .B2(new_n646), .ZN(G369));
  NAND3_X1  g0447(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G213), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g0452(.A(KEYINPUT83), .B(G343), .Z(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n598), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n629), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n604), .B2(new_n656), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G330), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n492), .A2(new_n499), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n626), .A2(new_n655), .ZN(new_n663));
  OAI22_X1  g0463(.A1(new_n662), .A2(new_n663), .B1(new_n492), .B2(new_n655), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n629), .A2(new_n655), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n662), .ZN(new_n667));
  INV_X1    g0467(.A(new_n655), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n492), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n665), .A2(new_n670), .ZN(G399));
  NOR2_X1   g0471(.A1(new_n215), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n220), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n673), .ZN(new_n677));
  XOR2_X1   g0477(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n678));
  XNOR2_X1  g0478(.A(new_n677), .B(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n668), .B1(new_n638), .B2(new_n644), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  XOR2_X1   g0481(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n642), .A2(new_n551), .A3(new_n572), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(KEYINPUT26), .ZN(new_n686));
  OAI211_X1 g0486(.A(KEYINPUT29), .B(new_n655), .C1(new_n686), .C2(new_n637), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n461), .A2(new_n509), .A3(new_n505), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(KEYINPUT30), .A3(new_n569), .A4(new_n601), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n601), .A2(new_n569), .A3(new_n461), .A4(new_n622), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n583), .A2(new_n524), .A3(new_n283), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n561), .A2(new_n566), .B1(new_n461), .B2(new_n462), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n690), .A2(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT85), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n689), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n690), .A2(new_n691), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n692), .A2(new_n693), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n697), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  OAI211_X1 g0499(.A(KEYINPUT31), .B(new_n668), .C1(new_n696), .C2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(new_n698), .A3(new_n689), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n668), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n700), .B(new_n704), .C1(new_n606), .C2(new_n668), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n683), .A2(new_n687), .B1(G330), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n679), .B1(new_n706), .B2(G1), .ZN(G364));
  NOR2_X1   g0507(.A1(new_n373), .A2(G179), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(G20), .A3(G190), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n580), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n212), .A2(new_n283), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n442), .A3(G200), .ZN(new_n712));
  INV_X1    g0512(.A(G317), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n713), .A2(KEYINPUT33), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(KEYINPUT33), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n212), .A2(G190), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G179), .A2(G200), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n710), .B(new_n716), .C1(G329), .C2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G190), .A2(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n711), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G311), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n325), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n711), .A2(G190), .A3(G200), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n725), .B1(G326), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n711), .A2(G190), .A3(new_n373), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n212), .B1(new_n718), .B2(G190), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n730), .A2(G322), .B1(new_n732), .B2(G294), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n717), .A2(new_n708), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT89), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G283), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n721), .A2(new_n728), .A3(new_n733), .A4(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n735), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n436), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n255), .B1(new_n712), .B2(new_n203), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n355), .A2(new_n709), .B1(new_n723), .B2(new_n258), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n726), .A2(new_n388), .B1(new_n731), .B2(new_n517), .ZN(new_n742));
  OR4_X1    g0542(.A1(new_n739), .A2(new_n740), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  XOR2_X1   g0543(.A(KEYINPUT88), .B(KEYINPUT32), .Z(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n719), .B2(new_n339), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n720), .A2(G159), .A3(new_n744), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n746), .B(new_n747), .C1(new_n202), .C2(new_n729), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n737), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n221), .B1(G20), .B2(new_n304), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n215), .A2(new_n325), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n752), .A2(G355), .B1(new_n468), .B2(new_n215), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n215), .A2(new_n255), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(new_n676), .B2(G45), .ZN(new_n755));
  INV_X1    g0555(.A(G45), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n249), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n753), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT87), .Z(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n750), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n214), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n211), .B1(new_n764), .B2(G45), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n672), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n751), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT90), .ZN(new_n769));
  INV_X1    g0569(.A(new_n761), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n658), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n661), .A2(new_n767), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G330), .B2(new_n658), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(G396));
  OAI22_X1  g0575(.A1(new_n443), .A2(new_n444), .B1(new_n434), .B2(new_n655), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n448), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n446), .A2(new_n447), .A3(new_n655), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n680), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n705), .A2(G330), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n767), .B1(new_n781), .B2(new_n782), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n750), .A2(new_n759), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G283), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n712), .A2(new_n788), .B1(new_n723), .B2(new_n468), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT91), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(new_n580), .B2(new_n726), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT92), .Z(new_n793));
  NAND2_X1  g0593(.A1(new_n735), .A2(G87), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G311), .A2(new_n720), .B1(new_n732), .B2(G97), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n794), .B(new_n795), .C1(new_n454), .C2(new_n729), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n325), .B1(new_n709), .B2(new_n436), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT93), .Z(new_n798));
  NOR2_X1   g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n712), .ZN(new_n800));
  INV_X1    g0600(.A(new_n723), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n800), .A2(G150), .B1(new_n801), .B2(G159), .ZN(new_n802));
  INV_X1    g0602(.A(G137), .ZN(new_n803));
  INV_X1    g0603(.A(G143), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n802), .B1(new_n803), .B2(new_n726), .C1(new_n804), .C2(new_n729), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT34), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n735), .A2(G68), .ZN(new_n808));
  INV_X1    g0608(.A(G132), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n255), .B1(new_n719), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n709), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n810), .B1(G50), .B2(new_n811), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n808), .B(new_n812), .C1(new_n202), .C2(new_n731), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n806), .B2(new_n805), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n793), .A2(new_n799), .B1(new_n807), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n750), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n767), .B1(G77), .B2(new_n787), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n760), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n779), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT94), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n785), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G384));
  NOR2_X1   g0622(.A1(new_n764), .A2(new_n211), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT39), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n348), .B1(new_n377), .B2(new_n378), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n338), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n321), .B1(new_n343), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n381), .B1(new_n827), .B2(new_n651), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n364), .ZN(new_n829));
  OAI21_X1  g0629(.A(KEYINPUT37), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n384), .A2(new_n376), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n367), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n652), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT37), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n381), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n827), .A2(new_n651), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n830), .A2(new_n835), .B1(new_n386), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n837), .A2(KEYINPUT97), .A3(KEYINPUT38), .ZN(new_n838));
  INV_X1    g0638(.A(new_n381), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n364), .B1(new_n384), .B2(new_n376), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT96), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT37), .A4(new_n833), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n832), .A2(new_n833), .A3(new_n381), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n651), .B1(new_n384), .B2(new_n376), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT37), .B1(new_n845), .B2(new_n842), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n386), .A2(new_n845), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT38), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n830), .A2(new_n835), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n386), .A2(new_n836), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT38), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT97), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n824), .B(new_n838), .C1(new_n850), .C2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n613), .A2(new_n403), .A3(new_n655), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT95), .Z(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT38), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n851), .B2(new_n852), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n856), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n609), .A2(new_n652), .ZN(new_n865));
  INV_X1    g0665(.A(new_n862), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n403), .A2(new_n668), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n423), .A2(new_n428), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n403), .B(new_n668), .C1(new_n613), .C2(new_n427), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n641), .A2(new_n643), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n655), .B(new_n780), .C1(new_n872), .C2(new_n637), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n873), .B2(new_n778), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n865), .B1(new_n866), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n864), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n682), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n450), .B(new_n687), .C1(new_n680), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n621), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n876), .B(new_n879), .ZN(new_n880));
  AND4_X1   g0680(.A1(KEYINPUT97), .A2(new_n851), .A3(new_n852), .A4(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT97), .B1(new_n837), .B2(KEYINPUT38), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n843), .A2(new_n847), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n386), .A2(new_n845), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n881), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n779), .B1(new_n868), .B2(new_n869), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n605), .A2(new_n642), .A3(new_n492), .A4(new_n499), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n889), .A2(new_n636), .A3(new_n668), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n701), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n704), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n888), .B(KEYINPUT40), .C1(new_n890), .C2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n704), .B(new_n891), .C1(new_n606), .C2(new_n668), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(new_n888), .C1(new_n860), .C2(new_n861), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n887), .A2(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n450), .A2(new_n895), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n660), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n898), .B2(new_n899), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n823), .B1(new_n880), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n880), .B2(new_n901), .ZN(new_n903));
  INV_X1    g0703(.A(new_n543), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n904), .A2(KEYINPUT35), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(KEYINPUT35), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n905), .A2(G116), .A3(new_n222), .A4(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT36), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n258), .B1(G58), .B2(G68), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n220), .A2(new_n909), .B1(new_n388), .B2(G68), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n214), .A2(G1), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n903), .B(new_n908), .C1(new_n910), .C2(new_n911), .ZN(G367));
  OAI211_X1 g0712(.A(new_n573), .B(new_n576), .C1(new_n635), .C2(new_n655), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n551), .A2(new_n572), .A3(new_n668), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n667), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT42), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n913), .A2(new_n492), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n668), .B1(new_n920), .B2(new_n573), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT100), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT100), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n919), .B2(new_n921), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n917), .A2(new_n918), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT43), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n522), .A2(new_n655), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(new_n624), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT98), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n625), .A2(new_n928), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n927), .B1(new_n934), .B2(KEYINPUT99), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(KEYINPUT99), .B2(new_n934), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n923), .A2(new_n925), .A3(new_n926), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT101), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n922), .A2(KEYINPUT100), .B1(new_n918), .B2(new_n917), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT101), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n939), .A2(new_n940), .A3(new_n925), .A4(new_n936), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n925), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n936), .B1(KEYINPUT43), .B2(new_n934), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n938), .A2(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n665), .A2(new_n915), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n672), .B(KEYINPUT41), .Z(new_n946));
  NAND2_X1  g0746(.A1(new_n913), .A2(new_n914), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n670), .ZN(new_n948));
  XOR2_X1   g0748(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n670), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT45), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n661), .A2(KEYINPUT103), .A3(new_n664), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n953), .B1(new_n950), .B2(new_n952), .ZN(new_n955));
  INV_X1    g0755(.A(new_n666), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n916), .B1(new_n664), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n661), .B(new_n957), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n954), .A2(new_n955), .A3(new_n706), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n946), .B1(new_n959), .B2(new_n706), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n944), .A2(new_n945), .B1(new_n960), .B2(new_n766), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n938), .A2(new_n941), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n942), .A2(new_n943), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n945), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT104), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n960), .A2(new_n766), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n964), .A2(new_n965), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT104), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n944), .A2(new_n945), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n754), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n240), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n762), .B1(new_n216), .B2(new_n432), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n731), .A2(new_n203), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n325), .B(new_n977), .C1(G159), .C2(new_n800), .ZN(new_n978));
  INV_X1    g0778(.A(new_n734), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n811), .A2(G58), .B1(new_n979), .B2(G77), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G50), .A2(new_n801), .B1(new_n720), .B2(G137), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G143), .A2(new_n727), .B1(new_n730), .B2(G150), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n811), .A2(G116), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT46), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n436), .B2(new_n731), .C1(new_n724), .C2(new_n726), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n325), .B1(new_n734), .B2(new_n517), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G303), .B2(new_n730), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n800), .A2(G294), .B1(new_n720), .B2(G317), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(new_n788), .C2(new_n723), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n983), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT47), .Z(new_n992));
  OAI221_X1 g0792(.A(new_n767), .B1(new_n975), .B2(new_n976), .C1(new_n992), .C2(new_n816), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT105), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n934), .A2(new_n770), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n973), .A2(new_n997), .ZN(G387));
  INV_X1    g0798(.A(new_n767), .ZN(new_n999));
  INV_X1    g0799(.A(new_n674), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n1000), .A2(new_n752), .B1(new_n436), .B2(new_n215), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n237), .A2(new_n756), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n319), .A2(new_n388), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT50), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n674), .B(new_n756), .C1(new_n203), .C2(new_n258), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n754), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1001), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n999), .B1(new_n1007), .B2(new_n762), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n664), .B2(new_n770), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n709), .A2(new_n258), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n325), .B(new_n1010), .C1(G150), .C2(new_n720), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n517), .B2(new_n738), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT106), .Z(new_n1013));
  OAI22_X1  g0813(.A1(new_n712), .A2(new_n289), .B1(new_n723), .B2(new_n203), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G50), .B2(new_n730), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n727), .A2(G159), .B1(new_n732), .B2(new_n525), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G311), .A2(new_n800), .B1(new_n727), .B2(G322), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT107), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n729), .A2(new_n713), .B1(new_n723), .B2(new_n580), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT108), .Z(new_n1023));
  AND2_X1   g0823(.A1(new_n1023), .A2(KEYINPUT48), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n811), .A2(G294), .B1(new_n732), .B2(G283), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n1023), .B2(KEYINPUT48), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(KEYINPUT49), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n734), .A2(new_n468), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n255), .B(new_n1029), .C1(G326), .C2(new_n720), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1027), .A2(KEYINPUT49), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1017), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1009), .B1(new_n1033), .B2(new_n750), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n766), .B2(new_n958), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n706), .A2(new_n958), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n672), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n706), .A2(new_n958), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1035), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(KEYINPUT109), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT109), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1041), .B(new_n1035), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1042), .ZN(G393));
  NOR2_X1   g0843(.A1(new_n950), .A2(new_n952), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n661), .A2(new_n664), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1036), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n672), .B(new_n959), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n766), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n762), .B1(new_n517), .B2(new_n216), .C1(new_n245), .C2(new_n974), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT110), .Z(new_n1051));
  AOI21_X1  g0851(.A(new_n325), .B1(new_n720), .B2(G143), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n794), .B(new_n1052), .C1(new_n203), .C2(new_n709), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT111), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n731), .A2(new_n258), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n712), .A2(new_n388), .B1(new_n723), .B2(new_n289), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n729), .A2(new_n339), .B1(new_n726), .B2(new_n286), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1057), .A2(KEYINPUT51), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(KEYINPUT51), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1055), .B(new_n1056), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n729), .A2(new_n724), .B1(new_n726), .B2(new_n713), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT52), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G294), .A2(new_n801), .B1(new_n720), .B2(G322), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n580), .B2(new_n712), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n325), .B1(new_n731), .B2(new_n468), .C1(new_n709), .C2(new_n788), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n739), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1054), .A2(new_n1060), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1051), .B(new_n767), .C1(new_n816), .C2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT112), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n770), .B2(new_n947), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1048), .A2(new_n1049), .A3(new_n1070), .ZN(G390));
  OAI211_X1 g0871(.A(new_n888), .B(G330), .C1(new_n890), .C2(new_n892), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT113), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT113), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n895), .A2(new_n1074), .A3(G330), .A4(new_n888), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n873), .A2(new_n778), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n870), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n856), .A2(new_n863), .B1(new_n1078), .B2(new_n858), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n655), .B(new_n777), .C1(new_n686), .C2(new_n637), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n778), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n870), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n887), .A2(new_n858), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1076), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n887), .A2(new_n1082), .A3(new_n858), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n705), .A2(G330), .A3(new_n780), .A4(new_n870), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n860), .A2(new_n861), .A3(new_n824), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n887), .B2(new_n824), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n874), .A2(new_n859), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1085), .B(new_n1086), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1084), .A2(new_n1090), .A3(new_n766), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT114), .Z(new_n1092));
  NAND2_X1  g0892(.A1(new_n1084), .A2(new_n1090), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n450), .A2(G330), .A3(new_n895), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n878), .A2(new_n621), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n705), .A2(G330), .A3(new_n780), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n871), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n1075), .A3(new_n1073), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n1077), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n895), .A2(G330), .A3(new_n780), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1081), .B1(new_n871), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n1086), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1095), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1093), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1084), .A2(new_n1090), .A3(new_n1103), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n672), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n255), .B1(new_n734), .B2(new_n388), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1108), .A2(KEYINPUT115), .B1(G125), .B2(new_n720), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(KEYINPUT115), .B2(new_n1108), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT116), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n800), .A2(G137), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n811), .A2(G150), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1112), .B1(new_n723), .B2(new_n1113), .C1(new_n1114), .C2(KEYINPUT53), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1114), .A2(KEYINPUT53), .B1(new_n727), .B2(G128), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1116), .B1(new_n809), .B2(new_n729), .C1(new_n339), .C2(new_n731), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n1111), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n255), .B(new_n1055), .C1(G87), .C2(new_n811), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G116), .A2(new_n730), .B1(new_n727), .B2(G283), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n723), .A2(new_n517), .B1(new_n719), .B2(new_n454), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G107), .B2(new_n800), .ZN(new_n1122));
  AND4_X1   g0922(.A1(new_n808), .A2(new_n1119), .A3(new_n1120), .A4(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n750), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n999), .B1(new_n289), .B2(new_n786), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(new_n1088), .C2(new_n760), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1092), .A2(new_n1107), .A3(new_n1126), .ZN(G378));
  INV_X1    g0927(.A(new_n1095), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1106), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n303), .A2(new_n652), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n620), .B2(new_n306), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1132), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n608), .B(new_n1134), .C1(new_n618), .C2(new_n619), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1131), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n318), .A2(new_n1134), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n620), .A2(new_n306), .A3(new_n1132), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n1138), .A3(new_n1130), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n898), .B2(G330), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n896), .A2(new_n897), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n894), .B(new_n838), .C1(new_n850), .C2(new_n855), .ZN(new_n1143));
  AND4_X1   g0943(.A1(G330), .A2(new_n1142), .A3(new_n1143), .A4(new_n1140), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n876), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n864), .A2(new_n875), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n898), .A2(G330), .A3(new_n1140), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1142), .A2(new_n1143), .A3(G330), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1140), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1146), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1145), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1129), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT57), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n673), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n1145), .B2(new_n1151), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1129), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT118), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT118), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1156), .A2(new_n1159), .A3(new_n1129), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1155), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1152), .A2(new_n766), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n767), .B1(G50), .B2(new_n787), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(G33), .A2(G41), .ZN(new_n1164));
  AOI211_X1 g0964(.A(G50), .B(new_n1164), .C1(new_n325), .C2(new_n268), .ZN(new_n1165));
  NOR4_X1   g0965(.A1(new_n1010), .A2(new_n977), .A3(G41), .A4(new_n255), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n800), .A2(G97), .B1(new_n801), .B2(new_n525), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n979), .A2(G58), .B1(new_n720), .B2(G283), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G107), .A2(new_n730), .B1(new_n727), .B2(G116), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT58), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1165), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n800), .A2(G132), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n709), .B2(new_n1113), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n727), .A2(G125), .B1(new_n732), .B2(G150), .ZN(new_n1175));
  INV_X1    g0975(.A(G128), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1175), .B1(new_n1176), .B2(new_n729), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1174), .B(new_n1177), .C1(G137), .C2(new_n801), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1164), .B1(new_n734), .B2(new_n339), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G124), .B2(new_n720), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT117), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT59), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1183), .B1(new_n1178), .B2(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1172), .B1(new_n1171), .B2(new_n1170), .C1(new_n1180), .C2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1163), .B1(new_n1186), .B2(new_n750), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1140), .B2(new_n760), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1162), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1161), .A2(new_n1190), .ZN(G375));
  INV_X1    g0991(.A(new_n946), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1098), .A2(new_n1077), .B1(new_n1101), .B2(new_n1086), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1095), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1104), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n767), .B1(G68), .B2(new_n787), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n712), .A2(new_n1113), .B1(new_n723), .B2(new_n286), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n325), .B(new_n1197), .C1(G58), .C2(new_n979), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n709), .A2(new_n339), .B1(new_n719), .B2(new_n1176), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT121), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n729), .A2(new_n803), .B1(new_n731), .B2(new_n388), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G132), .B2(new_n727), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1198), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n325), .B1(new_n723), .B2(new_n436), .C1(new_n468), .C2(new_n712), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G294), .B2(new_n727), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n811), .A2(G97), .B1(new_n720), .B2(G303), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT119), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT119), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n735), .A2(G77), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1205), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n729), .A2(new_n788), .B1(new_n731), .B2(new_n432), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT120), .Z(new_n1212));
  OAI21_X1  g1012(.A(new_n1203), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1196), .B1(new_n1213), .B2(new_n750), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n759), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1214), .B1(new_n870), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1193), .B2(new_n765), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1195), .A2(new_n1218), .ZN(G381));
  NOR2_X1   g1019(.A1(G375), .A2(G378), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1040), .A2(new_n774), .A3(new_n1042), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(new_n1221), .A2(G390), .A3(G381), .A4(G384), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1220), .A2(new_n973), .A3(new_n997), .A4(new_n1222), .ZN(G407));
  NAND2_X1  g1023(.A1(new_n653), .A2(G213), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1220), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(G407), .A2(G213), .A3(new_n1226), .ZN(G409));
  INV_X1    g1027(.A(G390), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G387), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1221), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n774), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT124), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1231), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT124), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1221), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n973), .A2(new_n997), .A3(G390), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1229), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(G390), .B1(new_n973), .B2(new_n997), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n996), .B(new_n1228), .C1(new_n967), .C2(new_n972), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1236), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT63), .ZN(new_n1244));
  INV_X1    g1044(.A(G378), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1190), .B1(new_n946), .B2(new_n1153), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1161), .A2(G378), .A3(new_n1190), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1225), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT60), .B1(new_n1193), .B2(new_n1095), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1194), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1193), .A2(KEYINPUT60), .A3(new_n1095), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n672), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT122), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n673), .B1(new_n1250), .B2(new_n1194), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(KEYINPUT122), .A3(new_n1252), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1217), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(new_n821), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1249), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1243), .B1(new_n1244), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1249), .A2(KEYINPUT63), .A3(new_n1259), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1257), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT122), .B1(new_n1256), .B2(new_n1252), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1218), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n821), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1258), .A2(G384), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1225), .A2(G2897), .ZN(new_n1269));
  XOR2_X1   g1069(.A(new_n1269), .B(KEYINPUT123), .Z(new_n1270));
  XNOR2_X1  g1070(.A(new_n1268), .B(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1249), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT61), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1261), .A2(new_n1262), .A3(new_n1273), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1275), .A2(new_n1273), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1243), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1274), .B1(new_n1277), .B2(new_n1278), .ZN(G405));
  AND3_X1   g1079(.A1(new_n1161), .A2(G378), .A3(new_n1190), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G378), .B1(new_n1161), .B2(new_n1190), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1259), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT125), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1259), .B(new_n1284), .C1(new_n1280), .C2(new_n1281), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1128), .A2(new_n1106), .B1(new_n1145), .B2(new_n1151), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n672), .B1(new_n1287), .B2(KEYINPUT57), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1156), .A2(new_n1159), .A3(new_n1129), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1159), .B1(new_n1156), .B2(new_n1129), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1245), .B1(new_n1291), .B2(new_n1189), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n1268), .A3(new_n1248), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT126), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1292), .A2(new_n1268), .A3(KEYINPUT126), .A4(new_n1248), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1286), .A2(new_n1297), .A3(new_n1243), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT127), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1286), .A2(new_n1297), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1278), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1286), .A2(new_n1297), .A3(new_n1243), .A4(KEYINPUT127), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1300), .A2(new_n1302), .A3(new_n1303), .ZN(G402));
endmodule


