//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955;
  AND2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G141gat), .B(G148gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT2), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n210));
  OR2_X1    g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n206), .A2(new_n209), .B1(new_n204), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT80), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT79), .B(KEYINPUT2), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n204), .B1(new_n205), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G155gat), .B(G162gat), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n220), .A2(new_n211), .A3(new_n209), .A4(new_n212), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT80), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT3), .ZN(new_n224));
  INV_X1    g023(.A(G127gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(G134gat), .ZN(new_n226));
  INV_X1    g025(.A(G134gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G127gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G113gat), .B2(G120gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G113gat), .A2(G120gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  OAI22_X1  g031(.A1(new_n226), .A2(new_n228), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G113gat), .ZN(new_n234));
  INV_X1    g033(.A(G120gat), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT1), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n227), .A2(G127gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n225), .A2(G134gat), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n236), .A2(new_n231), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n219), .A2(new_n216), .A3(new_n221), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n217), .A2(new_n224), .A3(new_n240), .A4(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n233), .A2(new_n239), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n215), .A2(KEYINPUT81), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT81), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n222), .B2(new_n240), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n246), .A3(KEYINPUT4), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n222), .B2(new_n240), .ZN(new_n249));
  NAND2_X1  g048(.A1(G225gat), .A2(G233gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n242), .A2(new_n247), .A3(new_n249), .A4(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT5), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n222), .A2(new_n240), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT81), .B1(new_n215), .B2(new_n243), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n222), .A2(new_n245), .A3(new_n240), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n254), .B1(new_n258), .B2(new_n251), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n251), .A2(new_n248), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(new_n256), .B2(new_n257), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n222), .A2(new_n248), .A3(new_n240), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n242), .A3(new_n264), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n259), .A2(KEYINPUT82), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT82), .B1(new_n259), .B2(new_n265), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n253), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G1gat), .B(G29gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT0), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G57gat), .ZN(new_n271));
  INV_X1    g070(.A(G85gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n268), .A2(KEYINPUT6), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n253), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n223), .B1(new_n222), .B2(KEYINPUT3), .ZN(new_n278));
  AOI211_X1 g077(.A(KEYINPUT80), .B(new_n216), .C1(new_n219), .C2(new_n221), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n241), .A2(new_n240), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n260), .B1(new_n244), .B2(new_n246), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n281), .A2(new_n282), .A3(new_n263), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n244), .A2(new_n246), .B1(new_n222), .B2(new_n240), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT5), .B1(new_n284), .B2(new_n250), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n277), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n259), .A2(new_n265), .A3(KEYINPUT82), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n276), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n288), .A2(KEYINPUT84), .A3(new_n273), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT84), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(new_n268), .B2(new_n274), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n253), .B(new_n273), .C1(new_n266), .C2(new_n267), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT83), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n273), .A2(new_n253), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(new_n286), .B2(new_n287), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT83), .B1(new_n298), .B2(KEYINPUT6), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n275), .B1(new_n292), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n302));
  XNOR2_X1  g101(.A(G64gat), .B(G92gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(G8gat), .B(G36gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n305), .B(new_n306), .Z(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G197gat), .B(G204gat), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n309), .B1(KEYINPUT22), .B2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G211gat), .B(G218gat), .Z(new_n314));
  AND2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n313), .A2(new_n314), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318));
  INV_X1    g117(.A(G169gat), .ZN(new_n319));
  INV_X1    g118(.A(G176gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT26), .ZN(new_n322));
  NAND2_X1  g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n318), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n331));
  INV_X1    g130(.A(G183gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT68), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n335), .B(new_n337), .C1(new_n338), .C2(G183gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT69), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(KEYINPUT27), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n338), .A2(KEYINPUT69), .ZN(new_n343));
  OAI211_X1 g142(.A(KEYINPUT70), .B(G183gat), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n333), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(KEYINPUT27), .B(G183gat), .Z(new_n349));
  NAND2_X1  g148(.A1(new_n335), .A2(new_n337), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n329), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT64), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT24), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n318), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n358), .B1(new_n318), .B2(new_n359), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT65), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n357), .B(KEYINPUT65), .C1(new_n360), .C2(new_n361), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT23), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT25), .B1(new_n321), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT66), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n320), .ZN(new_n369));
  NAND2_X1  g168(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n369), .A2(KEYINPUT23), .A3(new_n319), .A4(new_n370), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n367), .A2(new_n371), .A3(new_n327), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n364), .A2(new_n365), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT23), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n366), .B1(G169gat), .B2(G176gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n326), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n374), .B(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n355), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n350), .B2(G183gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT25), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n373), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G226gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n354), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(KEYINPUT29), .ZN(new_n389));
  INV_X1    g188(.A(new_n329), .ZN(new_n390));
  OAI21_X1  g189(.A(G183gat), .B1(new_n342), .B2(new_n343), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n339), .B1(new_n391), .B2(new_n330), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n346), .B1(new_n392), .B2(new_n344), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n390), .B1(new_n393), .B2(new_n352), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT25), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n379), .B2(new_n382), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n367), .A2(new_n371), .A3(new_n327), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(new_n363), .B2(new_n362), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n396), .B1(new_n398), .B2(new_n365), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n389), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n317), .B1(new_n388), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT75), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n394), .A2(new_n399), .A3(new_n386), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n313), .B(new_n314), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n354), .A2(new_n385), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n403), .B(new_n404), .C1(new_n405), .C2(new_n389), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(KEYINPUT75), .B(new_n317), .C1(new_n388), .C2(new_n400), .ZN(new_n408));
  AOI211_X1 g207(.A(new_n302), .B(new_n308), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n308), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT78), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT78), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n407), .A2(new_n408), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n307), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n413), .B(new_n410), .C1(new_n415), .C2(new_n302), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT30), .B1(new_n414), .B2(new_n307), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n301), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n404), .B1(new_n421), .B2(new_n241), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(G228gat), .B2(G233gat), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n404), .A2(KEYINPUT85), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n316), .B2(KEYINPUT85), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT3), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n426), .B2(new_n215), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n404), .A2(new_n421), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n215), .B1(new_n428), .B2(new_n216), .ZN(new_n429));
  OAI211_X1 g228(.A(G228gat), .B(G233gat), .C1(new_n429), .C2(new_n422), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G22gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n427), .A2(G22gat), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G78gat), .B(G106gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT31), .ZN(new_n437));
  INV_X1    g236(.A(G50gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n439), .A2(KEYINPUT86), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n439), .B(KEYINPUT86), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n433), .A2(new_n442), .A3(new_n434), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n286), .A2(new_n287), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n273), .B1(new_n446), .B2(new_n253), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n409), .A2(new_n411), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n448), .B2(new_n419), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT40), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n242), .A2(new_n247), .A3(new_n249), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n251), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n454), .A3(new_n273), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT39), .B1(new_n258), .B2(new_n251), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(new_n451), .B2(new_n251), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n454), .B1(new_n453), .B2(new_n273), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT88), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n450), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n459), .A2(new_n458), .ZN(new_n463));
  OAI211_X1 g262(.A(KEYINPUT88), .B(KEYINPUT40), .C1(new_n463), .C2(new_n456), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n445), .B1(new_n449), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n293), .A2(new_n295), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n275), .B1(new_n467), .B2(new_n447), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n308), .B1(new_n407), .B2(new_n408), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n307), .B1(new_n414), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n401), .A2(new_n406), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT38), .B1(new_n473), .B2(KEYINPUT37), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n407), .A2(KEYINPUT37), .A3(new_n408), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT38), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n472), .A2(KEYINPUT89), .A3(new_n474), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n470), .A2(new_n477), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n420), .A2(new_n445), .B1(new_n466), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n240), .B1(new_n354), .B2(new_n385), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT72), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n405), .A2(new_n243), .ZN(new_n486));
  NAND2_X1  g285(.A1(G227gat), .A2(G233gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT72), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(new_n240), .C1(new_n354), .C2(new_n385), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT34), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT73), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n490), .A2(KEYINPUT34), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT73), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n490), .A2(new_n495), .A3(KEYINPUT34), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT32), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n485), .A2(new_n489), .A3(new_n486), .ZN(new_n499));
  INV_X1    g298(.A(new_n487), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT33), .B1(new_n499), .B2(new_n500), .ZN(new_n502));
  XOR2_X1   g301(.A(G15gat), .B(G43gat), .Z(new_n503));
  XNOR2_X1  g302(.A(G71gat), .B(G99gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n501), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  AOI221_X4 g306(.A(new_n498), .B1(KEYINPUT33), .B2(new_n505), .C1(new_n499), .C2(new_n500), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n497), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n499), .A2(new_n500), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT33), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n506), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n501), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n493), .B1(KEYINPUT73), .B2(new_n491), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n501), .B1(new_n502), .B2(new_n506), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .A4(new_n496), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT36), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT36), .B1(new_n509), .B2(new_n517), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT74), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n517), .A3(KEYINPUT36), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n517), .A3(new_n444), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT35), .B1(new_n420), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n418), .A2(new_n409), .A3(new_n411), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(new_n468), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n530), .A3(new_n468), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n529), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n483), .A2(new_n526), .B1(new_n528), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT94), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT16), .ZN(new_n541));
  AOI21_X1  g340(.A(G1gat), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n540), .B(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NOR3_X1   g345(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n547));
  INV_X1    g346(.A(G29gat), .ZN(new_n548));
  INV_X1    g347(.A(G36gat), .ZN(new_n549));
  OAI22_X1  g348(.A1(new_n546), .A2(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G43gat), .B(G50gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(KEYINPUT15), .A3(new_n551), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n551), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(KEYINPUT15), .B2(new_n551), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n545), .B1(new_n547), .B2(KEYINPUT93), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(KEYINPUT93), .B2(new_n547), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n552), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n544), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n559), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n543), .A3(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(KEYINPUT18), .A3(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n543), .B(new_n557), .Z(new_n566));
  XOR2_X1   g365(.A(new_n564), .B(KEYINPUT13), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT18), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n558), .A2(new_n562), .ZN(new_n570));
  INV_X1    g369(.A(new_n564), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n565), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(KEYINPUT91), .B(KEYINPUT11), .Z(new_n574));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G169gat), .B(G197gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT92), .B(KEYINPUT12), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n568), .A3(new_n572), .ZN(new_n582));
  INV_X1    g381(.A(new_n580), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT95), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n581), .A2(new_n584), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G71gat), .B(G78gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT96), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(G57gat), .B(G64gat), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n593), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n593), .B(new_n592), .C1(new_n596), .C2(new_n595), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n543), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT97), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n605));
  XNOR2_X1  g404(.A(G127gat), .B(G155gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n604), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n608), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT7), .ZN(new_n616));
  NAND2_X1  g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  INV_X1    g416(.A(G92gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(KEYINPUT8), .A2(new_n617), .B1(new_n272), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G99gat), .B(G106gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(new_n559), .B2(new_n557), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n560), .ZN(new_n624));
  AND2_X1   g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n622), .A2(new_n557), .B1(KEYINPUT41), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G134gat), .B(G162gat), .Z(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT98), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n627), .B(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n631));
  XNOR2_X1  g430(.A(G190gat), .B(G218gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n630), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n614), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n601), .A2(KEYINPUT10), .A3(new_n622), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n640), .A2(KEYINPUT99), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n601), .A2(new_n622), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n601), .A2(new_n622), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n640), .A2(KEYINPUT99), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n641), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G176gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(G204gat), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n642), .A2(new_n644), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(G230gat), .A3(G233gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n649), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n648), .B(KEYINPUT100), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n654), .ZN(new_n659));
  INV_X1    g458(.A(new_n652), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(KEYINPUT101), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT101), .B1(new_n659), .B2(new_n660), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n655), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n639), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n536), .A2(new_n591), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n301), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  INV_X1    g469(.A(new_n531), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT103), .Z(new_n677));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678));
  OAI221_X1 g477(.A(new_n677), .B1(new_n678), .B2(new_n674), .C1(new_n539), .C2(new_n672), .ZN(G1325gat));
  INV_X1    g478(.A(new_n518), .ZN(new_n680));
  AOI21_X1  g479(.A(G15gat), .B1(new_n667), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n526), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(G15gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT104), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n667), .B2(new_n684), .ZN(G1326gat));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n445), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  NOR2_X1   g487(.A1(new_n536), .A2(new_n591), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n614), .A2(new_n664), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n638), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n548), .A3(new_n668), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n691), .A2(new_n585), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n420), .A2(new_n445), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n466), .A2(new_n482), .ZN(new_n701));
  INV_X1    g500(.A(new_n524), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n525), .B1(new_n523), .B2(KEYINPUT74), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n509), .A2(new_n517), .A3(new_n444), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n705), .A2(new_n301), .A3(new_n417), .A4(new_n419), .ZN(new_n706));
  AND4_X1   g505(.A1(new_n530), .A2(new_n468), .A3(new_n448), .A4(new_n419), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n532), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n706), .A2(KEYINPUT35), .B1(new_n708), .B2(new_n529), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n704), .B1(new_n709), .B2(KEYINPUT106), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n528), .A2(new_n535), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n699), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n712), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT107), .A4(new_n704), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n638), .A2(KEYINPUT44), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n714), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n638), .B1(new_n704), .B2(new_n711), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI211_X1 g522(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n536), .C2(new_n638), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n698), .B1(new_n719), .B2(new_n725), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n726), .A2(new_n668), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n696), .B1(new_n727), .B2(new_n548), .ZN(G1328gat));
  NOR3_X1   g527(.A1(new_n693), .A2(G36gat), .A3(new_n531), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT46), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n726), .A2(new_n671), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(new_n549), .ZN(G1329gat));
  INV_X1    g531(.A(G43gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n694), .A2(new_n733), .A3(new_n680), .ZN(new_n734));
  AOI211_X1 g533(.A(new_n526), .B(new_n698), .C1(new_n719), .C2(new_n725), .ZN(new_n735));
  OAI211_X1 g534(.A(KEYINPUT47), .B(new_n734), .C1(new_n735), .C2(new_n733), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT108), .B1(new_n735), .B2(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n725), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(new_n682), .A3(new_n697), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(new_n740), .A3(G43gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n737), .A2(new_n741), .A3(new_n734), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n742), .A2(KEYINPUT109), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT109), .B1(new_n742), .B2(new_n743), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n736), .B1(new_n744), .B2(new_n745), .ZN(G1330gat));
  AOI21_X1  g545(.A(new_n438), .B1(new_n726), .B2(new_n445), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n693), .A2(G50gat), .A3(new_n444), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  OAI22_X1  g548(.A1(new_n747), .A2(new_n748), .B1(KEYINPUT110), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(KEYINPUT110), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1331gat));
  AND2_X1   g551(.A1(new_n714), .A2(new_n717), .ZN(new_n753));
  INV_X1    g552(.A(new_n664), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n587), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n639), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n668), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g560(.A1(new_n758), .A2(new_n531), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  AND2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n762), .B2(new_n763), .ZN(G1333gat));
  OAI21_X1  g565(.A(G71gat), .B1(new_n758), .B2(new_n526), .ZN(new_n767));
  INV_X1    g566(.A(G71gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n680), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n758), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g570(.A1(new_n759), .A2(new_n445), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g572(.A1(new_n614), .A2(new_n587), .A3(new_n638), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n710), .B2(new_n713), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT51), .Z(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n754), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(new_n272), .A3(new_n668), .ZN(new_n779));
  AOI211_X1 g578(.A(new_n614), .B(new_n756), .C1(new_n719), .C2(new_n725), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n668), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(new_n272), .ZN(G1336gat));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n618), .A3(new_n671), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n618), .B1(new_n780), .B2(new_n671), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(KEYINPUT51), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n775), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n671), .A2(new_n664), .A3(new_n618), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n786), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n785), .A2(new_n786), .B1(new_n792), .B2(new_n784), .ZN(G1337gat));
  AOI21_X1  g592(.A(G99gat), .B1(new_n778), .B2(new_n680), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n682), .A2(G99gat), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n780), .B2(new_n795), .ZN(G1338gat));
  INV_X1    g595(.A(G106gat), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n780), .B2(new_n445), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n754), .A2(G106gat), .A3(new_n444), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n798), .B1(new_n789), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  INV_X1    g600(.A(new_n799), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n777), .B2(new_n802), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n800), .A2(new_n801), .B1(new_n798), .B2(new_n803), .ZN(G1339gat));
  INV_X1    g603(.A(new_n614), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n647), .A2(new_n806), .A3(new_n657), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(new_n660), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n649), .B(KEYINPUT54), .C1(new_n647), .C2(new_n657), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT55), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(new_n809), .A3(KEYINPUT55), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n587), .A2(new_n811), .A3(new_n655), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n570), .A2(new_n571), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n814), .A2(KEYINPUT112), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n566), .A2(new_n567), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(KEYINPUT112), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n818), .A2(new_n578), .B1(new_n573), .B2(new_n580), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n664), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n637), .B1(new_n813), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n637), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n812), .A2(new_n655), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n822), .A2(new_n823), .A3(new_n810), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n805), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n665), .A2(new_n585), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT113), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n825), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n445), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n301), .A2(new_n671), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n518), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n591), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT114), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n587), .A2(new_n234), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n836), .B2(new_n839), .ZN(G1340gat));
  NOR2_X1   g639(.A1(new_n836), .A2(new_n754), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(new_n235), .ZN(G1341gat));
  NOR2_X1   g641(.A1(new_n836), .A2(new_n805), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(new_n225), .ZN(G1342gat));
  NOR2_X1   g643(.A1(new_n836), .A2(new_n638), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n227), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n847), .B(new_n848), .C1(new_n227), .C2(new_n845), .ZN(G1343gat));
  AOI21_X1  g648(.A(new_n823), .B1(KEYINPUT116), .B2(new_n811), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n810), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n850), .A2(new_n586), .A3(new_n589), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n637), .B1(new_n853), .B2(new_n820), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n805), .B1(new_n854), .B2(new_n824), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(new_n826), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT57), .B1(new_n856), .B2(new_n444), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n682), .A2(new_n834), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT115), .ZN(new_n859));
  INV_X1    g658(.A(new_n830), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n829), .B1(new_n825), .B2(new_n826), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n445), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n857), .A2(new_n859), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(G141gat), .B1(new_n865), .B2(new_n591), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n862), .A2(new_n445), .A3(new_n858), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(G141gat), .A3(new_n591), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n866), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n865), .A2(new_n585), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n869), .B1(new_n872), .B2(G141gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n873), .B2(new_n867), .ZN(G1344gat));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n875), .B(G148gat), .C1(new_n865), .C2(new_n754), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n666), .A2(new_n590), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n855), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n878), .B(new_n863), .C1(new_n881), .C2(new_n444), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n862), .A2(new_n883), .A3(KEYINPUT57), .A4(new_n445), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n444), .B1(new_n855), .B2(new_n880), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT118), .B1(new_n885), .B2(KEYINPUT57), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n828), .A2(KEYINPUT57), .A3(new_n445), .A4(new_n830), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT117), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n882), .A2(new_n884), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n664), .A3(new_n859), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G148gat), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n877), .B1(new_n891), .B2(KEYINPUT59), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT119), .B(new_n875), .C1(new_n890), .C2(G148gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n876), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OR3_X1    g693(.A1(new_n868), .A2(G148gat), .A3(new_n754), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1345gat));
  OAI21_X1  g695(.A(G155gat), .B1(new_n865), .B2(new_n805), .ZN(new_n897));
  INV_X1    g696(.A(new_n868), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n207), .A3(new_n614), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n865), .B2(new_n638), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n208), .A3(new_n637), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n527), .A2(new_n531), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT120), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n831), .A2(new_n668), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n587), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n301), .A2(new_n671), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT121), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n909), .A2(new_n518), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n832), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n591), .A2(new_n319), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n907), .B1(new_n914), .B2(new_n915), .ZN(G1348gat));
  AOI21_X1  g715(.A(G176gat), .B1(new_n906), .B2(new_n664), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT123), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n754), .B1(new_n369), .B2(new_n370), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n914), .B2(new_n919), .ZN(G1349gat));
  AOI21_X1  g719(.A(new_n332), .B1(new_n914), .B2(new_n614), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n805), .A2(new_n349), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n906), .B2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT60), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(KEYINPUT60), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n924), .A2(KEYINPUT60), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n923), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n925), .A2(new_n928), .ZN(G1350gat));
  AOI21_X1  g728(.A(new_n334), .B1(new_n914), .B2(new_n637), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT61), .Z(new_n931));
  NAND4_X1  g730(.A1(new_n906), .A2(new_n335), .A3(new_n337), .A4(new_n637), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1351gat));
  NOR4_X1   g732(.A1(new_n831), .A2(new_n444), .A3(new_n682), .A4(new_n908), .ZN(new_n934));
  AOI21_X1  g733(.A(G197gat), .B1(new_n934), .B2(new_n587), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n682), .A2(new_n909), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT125), .Z(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(G197gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n938), .A2(new_n939), .A3(new_n591), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n935), .B1(new_n940), .B2(new_n889), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT126), .Z(G1352gat));
  XOR2_X1   g741(.A(KEYINPUT127), .B(G204gat), .Z(new_n943));
  NAND3_X1  g742(.A1(new_n934), .A2(new_n664), .A3(new_n943), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT62), .Z(new_n945));
  AND3_X1   g744(.A1(new_n889), .A2(new_n664), .A3(new_n937), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n943), .B2(new_n946), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n934), .A2(new_n310), .A3(new_n614), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n682), .A2(new_n909), .A3(new_n805), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n310), .B1(new_n889), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n950), .A2(KEYINPUT63), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(KEYINPUT63), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(G1354gat));
  AOI21_X1  g752(.A(G218gat), .B1(new_n934), .B2(new_n637), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n938), .A2(new_n311), .A3(new_n638), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n889), .ZN(G1355gat));
endmodule


