

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U549 ( .A(KEYINPUT65), .B(n538), .Z(n648) );
  XNOR2_X1 U550 ( .A(n519), .B(KEYINPUT17), .ZN(n885) );
  NOR2_X1 U551 ( .A1(n700), .A2(n921), .ZN(n702) );
  OR2_X1 U552 ( .A1(n711), .A2(n710), .ZN(n707) );
  INV_X1 U553 ( .A(KEYINPUT107), .ZN(n708) );
  AND2_X1 U554 ( .A1(n827), .A2(n817), .ZN(n512) );
  AND2_X1 U555 ( .A1(n512), .A2(n819), .ZN(n513) );
  AND2_X1 U556 ( .A1(G8), .A2(n740), .ZN(n514) );
  OR2_X1 U557 ( .A1(n782), .A2(n781), .ZN(n515) );
  NAND2_X1 U558 ( .A1(n748), .A2(n746), .ZN(n516) );
  AND2_X1 U559 ( .A1(n777), .A2(n776), .ZN(n517) );
  INV_X1 U560 ( .A(KEYINPUT64), .ZN(n701) );
  XNOR2_X1 U561 ( .A(n702), .B(n701), .ZN(n711) );
  XNOR2_X1 U562 ( .A(n709), .B(n708), .ZN(n713) );
  NOR2_X1 U563 ( .A1(n741), .A2(n514), .ZN(n742) );
  NAND2_X1 U564 ( .A1(n516), .A2(n742), .ZN(n772) );
  AND2_X1 U565 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U566 ( .A1(G164), .A2(G1384), .ZN(n784) );
  NOR2_X1 U567 ( .A1(n649), .A2(n541), .ZN(n642) );
  XOR2_X1 U568 ( .A(n597), .B(KEYINPUT15), .Z(n710) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XOR2_X1 U570 ( .A(KEYINPUT66), .B(n518), .Z(n519) );
  NAND2_X1 U571 ( .A1(n885), .A2(G138), .ZN(n526) );
  INV_X1 U572 ( .A(G2105), .ZN(n520) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n888) );
  NAND2_X1 U574 ( .A1(G114), .A2(n888), .ZN(n522) );
  NOR2_X1 U575 ( .A1(G2104), .A2(n520), .ZN(n890) );
  NAND2_X1 U576 ( .A1(G126), .A2(n890), .ZN(n521) );
  AND2_X1 U577 ( .A1(n522), .A2(n521), .ZN(n524) );
  AND2_X1 U578 ( .A1(n520), .A2(G2104), .ZN(n884) );
  NAND2_X1 U579 ( .A1(n884), .A2(G102), .ZN(n523) );
  AND2_X1 U580 ( .A1(n524), .A2(n523), .ZN(n525) );
  AND2_X1 U581 ( .A1(n526), .A2(n525), .ZN(G164) );
  XOR2_X1 U582 ( .A(G2443), .B(G2446), .Z(n528) );
  XNOR2_X1 U583 ( .A(G2427), .B(G2451), .ZN(n527) );
  XNOR2_X1 U584 ( .A(n528), .B(n527), .ZN(n534) );
  XOR2_X1 U585 ( .A(G2430), .B(G2454), .Z(n530) );
  XNOR2_X1 U586 ( .A(G1341), .B(G1348), .ZN(n529) );
  XNOR2_X1 U587 ( .A(n530), .B(n529), .ZN(n532) );
  XOR2_X1 U588 ( .A(G2435), .B(G2438), .Z(n531) );
  XNOR2_X1 U589 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U590 ( .A(n534), .B(n533), .Z(n535) );
  AND2_X1 U591 ( .A1(G14), .A2(n535), .ZN(G401) );
  INV_X1 U592 ( .A(G651), .ZN(n541) );
  NOR2_X1 U593 ( .A1(G543), .A2(n541), .ZN(n536) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n536), .Z(n653) );
  NAND2_X1 U595 ( .A1(G64), .A2(n653), .ZN(n540) );
  XNOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .ZN(n537) );
  XNOR2_X1 U597 ( .A(n537), .B(KEYINPUT67), .ZN(n649) );
  NOR2_X1 U598 ( .A1(G651), .A2(n649), .ZN(n538) );
  NAND2_X1 U599 ( .A1(G52), .A2(n648), .ZN(n539) );
  NAND2_X1 U600 ( .A1(n540), .A2(n539), .ZN(n547) );
  NOR2_X1 U601 ( .A1(G651), .A2(G543), .ZN(n639) );
  NAND2_X1 U602 ( .A1(G90), .A2(n639), .ZN(n543) );
  NAND2_X1 U603 ( .A1(G77), .A2(n642), .ZN(n542) );
  NAND2_X1 U604 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U605 ( .A(KEYINPUT9), .B(n544), .Z(n545) );
  XNOR2_X1 U606 ( .A(KEYINPUT70), .B(n545), .ZN(n546) );
  NOR2_X1 U607 ( .A1(n547), .A2(n546), .ZN(G171) );
  AND2_X1 U608 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U609 ( .A1(n888), .A2(G111), .ZN(n549) );
  NAND2_X1 U610 ( .A1(G135), .A2(n885), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n890), .A2(G123), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT18), .B(n550), .Z(n551) );
  NOR2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n884), .A2(G99), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n1001) );
  XNOR2_X1 U617 ( .A(G2096), .B(n1001), .ZN(n555) );
  OR2_X1 U618 ( .A1(G2100), .A2(n555), .ZN(G156) );
  INV_X1 U619 ( .A(G82), .ZN(G220) );
  NAND2_X1 U620 ( .A1(n888), .A2(G113), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G101), .A2(n884), .ZN(n556) );
  XOR2_X1 U622 ( .A(n556), .B(KEYINPUT23), .Z(n557) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n685) );
  NAND2_X1 U624 ( .A1(n890), .A2(G125), .ZN(n687) );
  NAND2_X1 U625 ( .A1(G137), .A2(n885), .ZN(n689) );
  NAND2_X1 U626 ( .A1(n687), .A2(n689), .ZN(n559) );
  NOR2_X1 U627 ( .A1(n685), .A2(n559), .ZN(G160) );
  NAND2_X1 U628 ( .A1(n639), .A2(G89), .ZN(n560) );
  XOR2_X1 U629 ( .A(KEYINPUT4), .B(n560), .Z(n563) );
  NAND2_X1 U630 ( .A1(n642), .A2(G76), .ZN(n561) );
  XOR2_X1 U631 ( .A(KEYINPUT82), .B(n561), .Z(n562) );
  NOR2_X1 U632 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U633 ( .A(KEYINPUT83), .B(n564), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n565), .B(KEYINPUT5), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G63), .A2(n653), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G51), .A2(n648), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n569) );
  XOR2_X1 U638 ( .A(KEYINPUT6), .B(KEYINPUT84), .Z(n568) );
  XNOR2_X1 U639 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U641 ( .A(KEYINPUT7), .B(n572), .ZN(G168) );
  XOR2_X1 U642 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U644 ( .A(n573), .B(KEYINPUT74), .ZN(n574) );
  XNOR2_X1 U645 ( .A(KEYINPUT10), .B(n574), .ZN(G223) );
  INV_X1 U646 ( .A(G223), .ZN(n837) );
  NAND2_X1 U647 ( .A1(n837), .A2(G567), .ZN(n575) );
  XOR2_X1 U648 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  XOR2_X1 U649 ( .A(G860), .B(KEYINPUT78), .Z(n609) );
  NAND2_X1 U650 ( .A1(G68), .A2(n642), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n639), .A2(G81), .ZN(n576) );
  XNOR2_X1 U652 ( .A(n576), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n578), .A2(n577), .ZN(n581) );
  XOR2_X1 U654 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n579) );
  XNOR2_X1 U655 ( .A(KEYINPUT13), .B(n579), .ZN(n580) );
  XNOR2_X1 U656 ( .A(n581), .B(n580), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n653), .A2(G56), .ZN(n582) );
  XNOR2_X1 U658 ( .A(KEYINPUT14), .B(n582), .ZN(n583) );
  NAND2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U660 ( .A(n585), .B(KEYINPUT77), .ZN(n587) );
  NAND2_X1 U661 ( .A1(G43), .A2(n648), .ZN(n586) );
  NAND2_X1 U662 ( .A1(n587), .A2(n586), .ZN(n921) );
  OR2_X1 U663 ( .A1(n609), .A2(n921), .ZN(G153) );
  INV_X1 U664 ( .A(G171), .ZN(G301) );
  NAND2_X1 U665 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U666 ( .A1(G92), .A2(n639), .ZN(n596) );
  NAND2_X1 U667 ( .A1(G79), .A2(n642), .ZN(n588) );
  XNOR2_X1 U668 ( .A(n588), .B(KEYINPUT80), .ZN(n591) );
  NAND2_X1 U669 ( .A1(G54), .A2(n648), .ZN(n589) );
  XOR2_X1 U670 ( .A(KEYINPUT81), .B(n589), .Z(n590) );
  NAND2_X1 U671 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G66), .A2(n653), .ZN(n592) );
  XNOR2_X1 U673 ( .A(KEYINPUT79), .B(n592), .ZN(n593) );
  NOR2_X1 U674 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n597) );
  INV_X1 U676 ( .A(G868), .ZN(n665) );
  NAND2_X1 U677 ( .A1(n710), .A2(n665), .ZN(n598) );
  NAND2_X1 U678 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U679 ( .A1(G91), .A2(n639), .ZN(n601) );
  NAND2_X1 U680 ( .A1(G78), .A2(n642), .ZN(n600) );
  NAND2_X1 U681 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U682 ( .A(KEYINPUT71), .B(n602), .ZN(n606) );
  NAND2_X1 U683 ( .A1(G65), .A2(n653), .ZN(n604) );
  NAND2_X1 U684 ( .A1(G53), .A2(n648), .ZN(n603) );
  AND2_X1 U685 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n606), .A2(n605), .ZN(G299) );
  NOR2_X1 U687 ( .A1(G286), .A2(n665), .ZN(n608) );
  NOR2_X1 U688 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U689 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U690 ( .A1(n609), .A2(G559), .ZN(n610) );
  INV_X1 U691 ( .A(n710), .ZN(n926) );
  NAND2_X1 U692 ( .A1(n610), .A2(n926), .ZN(n611) );
  XNOR2_X1 U693 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U694 ( .A1(G868), .A2(n921), .ZN(n614) );
  NAND2_X1 U695 ( .A1(G868), .A2(n926), .ZN(n612) );
  NOR2_X1 U696 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U697 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U698 ( .A1(G559), .A2(n926), .ZN(n615) );
  XNOR2_X1 U699 ( .A(n921), .B(n615), .ZN(n662) );
  NOR2_X1 U700 ( .A1(n662), .A2(G860), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G93), .A2(n639), .ZN(n617) );
  NAND2_X1 U702 ( .A1(G80), .A2(n642), .ZN(n616) );
  NAND2_X1 U703 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U704 ( .A1(G55), .A2(n648), .ZN(n618) );
  XNOR2_X1 U705 ( .A(KEYINPUT85), .B(n618), .ZN(n619) );
  NOR2_X1 U706 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n653), .A2(G67), .ZN(n621) );
  NAND2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n664) );
  XOR2_X1 U709 ( .A(n664), .B(KEYINPUT86), .Z(n623) );
  XNOR2_X1 U710 ( .A(n624), .B(n623), .ZN(G145) );
  NAND2_X1 U711 ( .A1(n653), .A2(G60), .ZN(n625) );
  XNOR2_X1 U712 ( .A(n625), .B(KEYINPUT68), .ZN(n627) );
  NAND2_X1 U713 ( .A1(G47), .A2(n648), .ZN(n626) );
  NAND2_X1 U714 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U715 ( .A(KEYINPUT69), .B(n628), .ZN(n632) );
  NAND2_X1 U716 ( .A1(G85), .A2(n639), .ZN(n630) );
  NAND2_X1 U717 ( .A1(G72), .A2(n642), .ZN(n629) );
  AND2_X1 U718 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U719 ( .A1(n632), .A2(n631), .ZN(G290) );
  NAND2_X1 U720 ( .A1(G88), .A2(n639), .ZN(n634) );
  NAND2_X1 U721 ( .A1(G75), .A2(n642), .ZN(n633) );
  NAND2_X1 U722 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U723 ( .A1(G62), .A2(n653), .ZN(n636) );
  NAND2_X1 U724 ( .A1(G50), .A2(n648), .ZN(n635) );
  NAND2_X1 U725 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U726 ( .A1(n638), .A2(n637), .ZN(G166) );
  NAND2_X1 U727 ( .A1(G61), .A2(n653), .ZN(n641) );
  NAND2_X1 U728 ( .A1(G86), .A2(n639), .ZN(n640) );
  NAND2_X1 U729 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U730 ( .A1(n642), .A2(G73), .ZN(n643) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U732 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U733 ( .A1(n648), .A2(G48), .ZN(n646) );
  NAND2_X1 U734 ( .A1(n647), .A2(n646), .ZN(G305) );
  NAND2_X1 U735 ( .A1(G49), .A2(n648), .ZN(n651) );
  NAND2_X1 U736 ( .A1(G87), .A2(n649), .ZN(n650) );
  NAND2_X1 U737 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U738 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U739 ( .A1(G651), .A2(G74), .ZN(n654) );
  NAND2_X1 U740 ( .A1(n655), .A2(n654), .ZN(G288) );
  XNOR2_X1 U741 ( .A(KEYINPUT19), .B(KEYINPUT87), .ZN(n657) );
  XNOR2_X1 U742 ( .A(G290), .B(G166), .ZN(n656) );
  XNOR2_X1 U743 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U744 ( .A(n658), .B(G299), .ZN(n659) );
  XNOR2_X1 U745 ( .A(n659), .B(n664), .ZN(n660) );
  XNOR2_X1 U746 ( .A(n660), .B(G305), .ZN(n661) );
  XNOR2_X1 U747 ( .A(n661), .B(G288), .ZN(n905) );
  XOR2_X1 U748 ( .A(n662), .B(n905), .Z(n663) );
  NAND2_X1 U749 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U750 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U751 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2084), .A2(G2078), .ZN(n670) );
  XNOR2_X1 U753 ( .A(KEYINPUT88), .B(KEYINPUT20), .ZN(n668) );
  XNOR2_X1 U754 ( .A(n668), .B(KEYINPUT89), .ZN(n669) );
  XNOR2_X1 U755 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U756 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U757 ( .A(n672), .B(KEYINPUT90), .ZN(n673) );
  XNOR2_X1 U758 ( .A(n673), .B(KEYINPUT21), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n674), .A2(G2072), .ZN(n675) );
  XOR2_X1 U760 ( .A(KEYINPUT91), .B(n675), .Z(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U762 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  XOR2_X1 U763 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  XNOR2_X1 U766 ( .A(n677), .B(KEYINPUT92), .ZN(n678) );
  NOR2_X1 U767 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U768 ( .A1(G96), .A2(n679), .ZN(n842) );
  NAND2_X1 U769 ( .A1(n842), .A2(G2106), .ZN(n683) );
  NAND2_X1 U770 ( .A1(G108), .A2(G120), .ZN(n680) );
  NOR2_X1 U771 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U772 ( .A1(G69), .A2(n681), .ZN(n841) );
  NAND2_X1 U773 ( .A1(G567), .A2(n841), .ZN(n682) );
  NAND2_X1 U774 ( .A1(n683), .A2(n682), .ZN(n917) );
  NAND2_X1 U775 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U776 ( .A1(n917), .A2(n684), .ZN(n840) );
  NAND2_X1 U777 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U778 ( .A(G166), .ZN(G303) );
  INV_X1 U779 ( .A(G40), .ZN(n686) );
  NOR2_X1 U780 ( .A1(n686), .A2(n685), .ZN(n688) );
  AND2_X1 U781 ( .A1(n688), .A2(n687), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n783) );
  NAND2_X1 U783 ( .A1(KEYINPUT101), .A2(n783), .ZN(n694) );
  INV_X1 U784 ( .A(KEYINPUT101), .ZN(n692) );
  AND2_X1 U785 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U786 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n703) );
  AND2_X1 U788 ( .A1(n784), .A2(G1996), .ZN(n695) );
  AND2_X1 U789 ( .A1(n703), .A2(n695), .ZN(n697) );
  XOR2_X1 U790 ( .A(KEYINPUT26), .B(KEYINPUT106), .Z(n696) );
  XNOR2_X1 U791 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n703), .A2(n784), .ZN(n732) );
  NAND2_X1 U793 ( .A1(n732), .A2(G1341), .ZN(n698) );
  NAND2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n700) );
  AND2_X1 U795 ( .A1(n703), .A2(n784), .ZN(n726) );
  NOR2_X1 U796 ( .A1(n726), .A2(G1348), .ZN(n705) );
  NOR2_X1 U797 ( .A1(G2067), .A2(n732), .ZN(n704) );
  NOR2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U801 ( .A1(n713), .A2(n712), .ZN(n718) );
  INV_X1 U802 ( .A(G299), .ZN(n927) );
  NAND2_X1 U803 ( .A1(n726), .A2(G2072), .ZN(n714) );
  XNOR2_X1 U804 ( .A(n714), .B(KEYINPUT27), .ZN(n716) );
  INV_X1 U805 ( .A(G1956), .ZN(n947) );
  NOR2_X1 U806 ( .A1(n947), .A2(n726), .ZN(n715) );
  NOR2_X1 U807 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U808 ( .A1(n927), .A2(n719), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n718), .A2(n717), .ZN(n723) );
  NOR2_X1 U810 ( .A1(n927), .A2(n719), .ZN(n721) );
  XNOR2_X1 U811 ( .A(KEYINPUT28), .B(KEYINPUT105), .ZN(n720) );
  XNOR2_X1 U812 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n725) );
  XOR2_X1 U814 ( .A(KEYINPUT29), .B(KEYINPUT108), .Z(n724) );
  XNOR2_X1 U815 ( .A(n725), .B(n724), .ZN(n730) );
  XOR2_X1 U816 ( .A(G1961), .B(KEYINPUT104), .Z(n942) );
  NOR2_X1 U817 ( .A1(n726), .A2(n942), .ZN(n728) );
  XNOR2_X1 U818 ( .A(G2078), .B(KEYINPUT25), .ZN(n973) );
  NOR2_X1 U819 ( .A1(n732), .A2(n973), .ZN(n727) );
  NOR2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n731) );
  NAND2_X1 U821 ( .A1(G171), .A2(n731), .ZN(n729) );
  NAND2_X1 U822 ( .A1(n730), .A2(n729), .ZN(n748) );
  NOR2_X1 U823 ( .A1(G171), .A2(n731), .ZN(n737) );
  NAND2_X1 U824 ( .A1(G8), .A2(n732), .ZN(n782) );
  NOR2_X1 U825 ( .A1(G1966), .A2(n782), .ZN(n741) );
  NOR2_X1 U826 ( .A1(G2084), .A2(n732), .ZN(n740) );
  NOR2_X1 U827 ( .A1(n741), .A2(n740), .ZN(n733) );
  NAND2_X1 U828 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U829 ( .A(KEYINPUT30), .B(n734), .ZN(n735) );
  NOR2_X1 U830 ( .A1(G168), .A2(n735), .ZN(n736) );
  NOR2_X1 U831 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U832 ( .A(n738), .B(KEYINPUT31), .ZN(n739) );
  XNOR2_X1 U833 ( .A(n739), .B(KEYINPUT109), .ZN(n746) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n932) );
  AND2_X1 U835 ( .A1(n772), .A2(n932), .ZN(n755) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n782), .ZN(n744) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n732), .ZN(n743) );
  NOR2_X1 U838 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U839 ( .A1(n745), .A2(G303), .ZN(n749) );
  AND2_X1 U840 ( .A1(n746), .A2(n749), .ZN(n747) );
  NAND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n752) );
  INV_X1 U842 ( .A(n749), .ZN(n750) );
  OR2_X1 U843 ( .A1(n750), .A2(G286), .ZN(n751) );
  AND2_X1 U844 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U845 ( .A1(n753), .A2(G8), .ZN(n754) );
  XNOR2_X1 U846 ( .A(n754), .B(KEYINPUT32), .ZN(n771) );
  NAND2_X1 U847 ( .A1(n755), .A2(n771), .ZN(n762) );
  INV_X1 U848 ( .A(KEYINPUT33), .ZN(n760) );
  INV_X1 U849 ( .A(n932), .ZN(n757) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n764) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U852 ( .A1(n764), .A2(n756), .ZN(n933) );
  OR2_X1 U853 ( .A1(n757), .A2(n933), .ZN(n758) );
  OR2_X1 U854 ( .A1(n782), .A2(n758), .ZN(n759) );
  AND2_X1 U855 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U856 ( .A(n763), .B(KEYINPUT110), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n764), .A2(KEYINPUT33), .ZN(n765) );
  NOR2_X1 U858 ( .A1(n782), .A2(n765), .ZN(n766) );
  NOR2_X1 U859 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U860 ( .A(G1981), .B(G305), .Z(n918) );
  NAND2_X1 U861 ( .A1(n768), .A2(n918), .ZN(n777) );
  NOR2_X1 U862 ( .A1(G2090), .A2(G303), .ZN(n769) );
  XOR2_X1 U863 ( .A(KEYINPUT111), .B(n769), .Z(n770) );
  NAND2_X1 U864 ( .A1(G8), .A2(n770), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n775), .A2(n782), .ZN(n776) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n780) );
  XNOR2_X1 U869 ( .A(KEYINPUT24), .B(KEYINPUT103), .ZN(n778) );
  XNOR2_X1 U870 ( .A(n778), .B(KEYINPUT102), .ZN(n779) );
  XNOR2_X1 U871 ( .A(n780), .B(n779), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n517), .A2(n515), .ZN(n820) );
  NOR2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n832) );
  NAND2_X1 U874 ( .A1(n884), .A2(G104), .ZN(n785) );
  XNOR2_X1 U875 ( .A(n785), .B(KEYINPUT94), .ZN(n787) );
  NAND2_X1 U876 ( .A1(G140), .A2(n885), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(n788), .ZN(n795) );
  NAND2_X1 U879 ( .A1(n890), .A2(G128), .ZN(n789) );
  XNOR2_X1 U880 ( .A(KEYINPUT95), .B(n789), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n888), .A2(G116), .ZN(n790) );
  XOR2_X1 U882 ( .A(KEYINPUT96), .B(n790), .Z(n791) );
  NOR2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U884 ( .A(n793), .B(KEYINPUT35), .ZN(n794) );
  NOR2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U886 ( .A(KEYINPUT36), .B(n796), .ZN(n901) );
  XNOR2_X1 U887 ( .A(KEYINPUT37), .B(G2067), .ZN(n829) );
  NOR2_X1 U888 ( .A1(n901), .A2(n829), .ZN(n994) );
  NAND2_X1 U889 ( .A1(n832), .A2(n994), .ZN(n827) );
  NAND2_X1 U890 ( .A1(G95), .A2(n884), .ZN(n798) );
  NAND2_X1 U891 ( .A1(G119), .A2(n890), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n888), .A2(G107), .ZN(n800) );
  NAND2_X1 U894 ( .A1(G131), .A2(n885), .ZN(n799) );
  NAND2_X1 U895 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U897 ( .A(n803), .B(KEYINPUT97), .ZN(n876) );
  NAND2_X1 U898 ( .A1(G1991), .A2(n876), .ZN(n804) );
  XOR2_X1 U899 ( .A(KEYINPUT98), .B(n804), .Z(n815) );
  NAND2_X1 U900 ( .A1(G105), .A2(n884), .ZN(n805) );
  XNOR2_X1 U901 ( .A(n805), .B(KEYINPUT38), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G117), .A2(n888), .ZN(n807) );
  NAND2_X1 U903 ( .A1(G129), .A2(n890), .ZN(n806) );
  NAND2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U905 ( .A1(G141), .A2(n885), .ZN(n808) );
  XNOR2_X1 U906 ( .A(KEYINPUT99), .B(n808), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U908 ( .A1(n812), .A2(n811), .ZN(n879) );
  NAND2_X1 U909 ( .A1(G1996), .A2(n879), .ZN(n813) );
  XOR2_X1 U910 ( .A(KEYINPUT100), .B(n813), .Z(n814) );
  NOR2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n1011) );
  INV_X1 U912 ( .A(n832), .ZN(n816) );
  NOR2_X1 U913 ( .A1(n1011), .A2(n816), .ZN(n823) );
  INV_X1 U914 ( .A(n823), .ZN(n817) );
  XOR2_X1 U915 ( .A(G1986), .B(KEYINPUT93), .Z(n818) );
  XNOR2_X1 U916 ( .A(G290), .B(n818), .ZN(n923) );
  NAND2_X1 U917 ( .A1(n923), .A2(n832), .ZN(n819) );
  NAND2_X1 U918 ( .A1(n820), .A2(n513), .ZN(n835) );
  NOR2_X1 U919 ( .A1(G1991), .A2(n876), .ZN(n1004) );
  NOR2_X1 U920 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U921 ( .A1(n1004), .A2(n821), .ZN(n822) );
  NOR2_X1 U922 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U923 ( .A1(G1996), .A2(n879), .ZN(n997) );
  NOR2_X1 U924 ( .A1(n824), .A2(n997), .ZN(n825) );
  XNOR2_X1 U925 ( .A(n825), .B(KEYINPUT39), .ZN(n826) );
  XNOR2_X1 U926 ( .A(n826), .B(KEYINPUT112), .ZN(n828) );
  NAND2_X1 U927 ( .A1(n828), .A2(n827), .ZN(n830) );
  NAND2_X1 U928 ( .A1(n901), .A2(n829), .ZN(n993) );
  NAND2_X1 U929 ( .A1(n830), .A2(n993), .ZN(n831) );
  XOR2_X1 U930 ( .A(KEYINPUT113), .B(n831), .Z(n833) );
  NAND2_X1 U931 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U932 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n836), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U936 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U938 ( .A1(n840), .A2(n839), .ZN(G188) );
  NOR2_X1 U939 ( .A1(n842), .A2(n841), .ZN(G325) );
  XOR2_X1 U940 ( .A(KEYINPUT114), .B(G325), .Z(G261) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  INV_X1 U943 ( .A(G108), .ZN(G238) );
  INV_X1 U944 ( .A(G69), .ZN(G235) );
  XOR2_X1 U945 ( .A(G2678), .B(G2090), .Z(n844) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U947 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U948 ( .A(n845), .B(G2100), .Z(n847) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U951 ( .A(G2096), .B(KEYINPUT115), .Z(n849) );
  XNOR2_X1 U952 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n848) );
  XNOR2_X1 U953 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U954 ( .A(n851), .B(n850), .Z(G227) );
  XOR2_X1 U955 ( .A(G1976), .B(G1971), .Z(n853) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1961), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U958 ( .A(n854), .B(G2474), .Z(n856) );
  XNOR2_X1 U959 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U960 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U961 ( .A(KEYINPUT41), .B(G1981), .Z(n858) );
  XNOR2_X1 U962 ( .A(G1966), .B(G1956), .ZN(n857) );
  XNOR2_X1 U963 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U964 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U965 ( .A1(G124), .A2(n890), .ZN(n861) );
  XNOR2_X1 U966 ( .A(n861), .B(KEYINPUT116), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U968 ( .A1(G112), .A2(n888), .ZN(n863) );
  NAND2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n884), .A2(G100), .ZN(n866) );
  NAND2_X1 U971 ( .A1(G136), .A2(n885), .ZN(n865) );
  NAND2_X1 U972 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U973 ( .A1(n868), .A2(n867), .ZN(G162) );
  NAND2_X1 U974 ( .A1(G118), .A2(n888), .ZN(n870) );
  NAND2_X1 U975 ( .A1(G130), .A2(n890), .ZN(n869) );
  NAND2_X1 U976 ( .A1(n870), .A2(n869), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n884), .A2(G106), .ZN(n872) );
  NAND2_X1 U978 ( .A1(G142), .A2(n885), .ZN(n871) );
  NAND2_X1 U979 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U980 ( .A(n873), .B(KEYINPUT45), .Z(n874) );
  NOR2_X1 U981 ( .A1(n875), .A2(n874), .ZN(n877) );
  XNOR2_X1 U982 ( .A(n877), .B(n876), .ZN(n900) );
  XOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n878) );
  XNOR2_X1 U984 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U985 ( .A(n880), .B(KEYINPUT46), .Z(n882) );
  XNOR2_X1 U986 ( .A(G164), .B(KEYINPUT120), .ZN(n881) );
  XNOR2_X1 U987 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U988 ( .A(n1001), .B(n883), .ZN(n898) );
  NAND2_X1 U989 ( .A1(n884), .A2(G103), .ZN(n887) );
  NAND2_X1 U990 ( .A1(G139), .A2(n885), .ZN(n886) );
  NAND2_X1 U991 ( .A1(n887), .A2(n886), .ZN(n896) );
  NAND2_X1 U992 ( .A1(n888), .A2(G115), .ZN(n889) );
  XNOR2_X1 U993 ( .A(KEYINPUT119), .B(n889), .ZN(n893) );
  NAND2_X1 U994 ( .A1(n890), .A2(G127), .ZN(n891) );
  XOR2_X1 U995 ( .A(KEYINPUT118), .B(n891), .Z(n892) );
  NOR2_X1 U996 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U997 ( .A(n894), .B(KEYINPUT47), .ZN(n895) );
  NOR2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n1007) );
  XNOR2_X1 U999 ( .A(G160), .B(n1007), .ZN(n897) );
  XNOR2_X1 U1000 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U1001 ( .A(n900), .B(n899), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n901), .B(G162), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n904), .ZN(G395) );
  XOR2_X1 U1005 ( .A(n905), .B(G286), .Z(n907) );
  XNOR2_X1 U1006 ( .A(G171), .B(n926), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1008 ( .A(n908), .B(n921), .Z(n909) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(KEYINPUT122), .B(KEYINPUT49), .ZN(n910) );
  XNOR2_X1 U1012 ( .A(n911), .B(n910), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n917), .ZN(n912) );
  XNOR2_X1 U1014 ( .A(KEYINPUT121), .B(n912), .ZN(n913) );
  NOR2_X1 U1015 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(n917), .ZN(G319) );
  INV_X1 U1020 ( .A(G96), .ZN(G221) );
  XOR2_X1 U1021 ( .A(G16), .B(KEYINPUT56), .Z(n941) );
  XNOR2_X1 U1022 ( .A(G1966), .B(G168), .ZN(n919) );
  NAND2_X1 U1023 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1024 ( .A(n920), .B(KEYINPUT57), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(G1341), .B(n921), .ZN(n922) );
  NOR2_X1 U1026 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n939) );
  XNOR2_X1 U1028 ( .A(n926), .B(G1348), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(n927), .B(G1956), .ZN(n928) );
  NAND2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(G1961), .B(G301), .ZN(n930) );
  NOR2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n937) );
  AND2_X1 U1033 ( .A1(G303), .A2(G1971), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n991) );
  XOR2_X1 U1039 ( .A(n942), .B(G5), .Z(n944) );
  XNOR2_X1 U1040 ( .A(G21), .B(G1966), .ZN(n943) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n956) );
  XOR2_X1 U1042 ( .A(G4), .B(KEYINPUT126), .Z(n946) );
  XNOR2_X1 U1043 ( .A(G1348), .B(KEYINPUT59), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(n946), .B(n945), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(G20), .B(n947), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(G1341), .B(G19), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(G6), .B(G1981), .ZN(n948) );
  NOR2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n954), .B(KEYINPUT60), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G22), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G23), .B(G1976), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n960) );
  XOR2_X1 U1056 ( .A(G1986), .B(G24), .Z(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(KEYINPUT58), .B(n961), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1060 ( .A(KEYINPUT61), .B(n964), .Z(n965) );
  NOR2_X1 U1061 ( .A1(G16), .A2(n965), .ZN(n988) );
  XNOR2_X1 U1062 ( .A(G1996), .B(G32), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(G33), .B(G2072), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n972) );
  XOR2_X1 U1065 ( .A(G1991), .B(G25), .Z(n968) );
  NAND2_X1 U1066 ( .A1(n968), .A2(G28), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(G26), .B(G2067), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1070 ( .A(G27), .B(n973), .Z(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(KEYINPUT123), .B(n976), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(n977), .B(KEYINPUT53), .ZN(n981) );
  XOR2_X1 U1074 ( .A(KEYINPUT124), .B(G34), .Z(n979) );
  XNOR2_X1 U1075 ( .A(G2084), .B(KEYINPUT54), .ZN(n978) );
  XNOR2_X1 U1076 ( .A(n979), .B(n978), .ZN(n980) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(G35), .B(G2090), .ZN(n982) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(KEYINPUT55), .B(n984), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(KEYINPUT125), .B(n985), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(G29), .A2(n986), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(G11), .A2(n989), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(n992), .B(KEYINPUT127), .ZN(n1020) );
  INV_X1 U1087 ( .A(G29), .ZN(n1018) );
  INV_X1 U1088 ( .A(n993), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n1006) );
  XOR2_X1 U1090 ( .A(G160), .B(G2084), .Z(n1000) );
  XOR2_X1 U1091 ( .A(G2090), .B(G162), .Z(n996) );
  NOR2_X1 U1092 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1093 ( .A(KEYINPUT51), .B(n998), .ZN(n999) );
  NOR2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1014) );
  XOR2_X1 U1098 ( .A(G2072), .B(n1007), .Z(n1009) );
  XOR2_X1 U1099 ( .A(G164), .B(G2078), .Z(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(KEYINPUT50), .B(n1010), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1104 ( .A(KEYINPUT52), .B(n1015), .Z(n1016) );
  NOR2_X1 U1105 ( .A1(KEYINPUT55), .A2(n1016), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1021), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

