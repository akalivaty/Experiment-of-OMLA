//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n192), .A3(new_n196), .A4(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  OR2_X1    g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  AOI22_X1  g018(.A1(new_n200), .A2(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n200), .A2(new_n202), .A3(new_n204), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT66), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n204), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(new_n202), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n200), .A2(new_n202), .A3(new_n204), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n198), .A2(new_n207), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n189), .A2(G137), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n191), .A2(G134), .ZN(new_n216));
  OAI21_X1  g030(.A(G131), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n197), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n200), .A3(new_n202), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n199), .A3(G143), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n201), .B(G146), .C1(new_n219), .C2(KEYINPUT1), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT67), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n221), .A2(new_n226), .A3(new_n222), .A4(new_n223), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n218), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT2), .ZN(new_n229));
  INV_X1    g043(.A(G113), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT65), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(KEYINPUT2), .B2(G113), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n231), .A2(new_n233), .B1(KEYINPUT2), .B2(G113), .ZN(new_n234));
  XNOR2_X1  g048(.A(G116), .B(G119), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n214), .A2(new_n228), .A3(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n187), .B1(new_n237), .B2(KEYINPUT28), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n225), .A2(new_n227), .ZN(new_n239));
  INV_X1    g053(.A(new_n218), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n235), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n234), .B(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n198), .A2(new_n207), .A3(new_n213), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT28), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(KEYINPUT72), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n238), .A2(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(new_n218), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n195), .A2(new_n197), .B1(new_n210), .B2(new_n212), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n236), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n245), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT71), .B1(new_n253), .B2(KEYINPUT28), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n255));
  AOI211_X1 g069(.A(new_n255), .B(new_n246), .C1(new_n245), .C2(new_n252), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n248), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT73), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n250), .B2(new_n251), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT64), .ZN(new_n268));
  NOR4_X1   g082(.A1(new_n214), .A2(new_n228), .A3(KEYINPUT68), .A4(new_n266), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n214), .A2(new_n228), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(KEYINPUT30), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n268), .B(new_n236), .C1(new_n269), .C2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n264), .A3(new_n245), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT31), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n273), .A2(new_n264), .A3(new_n245), .A4(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n278));
  INV_X1    g092(.A(new_n252), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT28), .B1(new_n237), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n255), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n253), .A2(KEYINPUT71), .A3(KEYINPUT28), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n278), .B(new_n263), .C1(new_n283), .C2(new_n248), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n265), .A2(new_n275), .A3(new_n277), .A4(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT32), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n248), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n271), .A2(new_n243), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT28), .B1(new_n291), .B2(new_n237), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n263), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n273), .A2(new_n245), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n263), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n254), .A2(new_n256), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n300), .A2(new_n290), .A3(new_n301), .A4(new_n264), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n302), .A3(new_n295), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n257), .B2(new_n264), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n297), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G472), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n285), .A2(KEYINPUT32), .A3(new_n286), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n289), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G217), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(G234), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G110), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G128), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n317));
  OAI22_X1  g131(.A1(new_n317), .A2(KEYINPUT23), .B1(new_n219), .B2(G119), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT76), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n316), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n317), .A2(KEYINPUT23), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n314), .A2(G128), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(KEYINPUT76), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .A4(KEYINPUT77), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n315), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n315), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(KEYINPUT23), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n313), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT80), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT24), .B(G110), .Z(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT75), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n323), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(KEYINPUT80), .B(new_n313), .C1(new_n326), .C2(new_n328), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n331), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G140), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT78), .A3(G125), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n340));
  INV_X1    g154(.A(G125), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(G140), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(G140), .ZN(new_n343));
  OAI211_X1 g157(.A(KEYINPUT16), .B(new_n339), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT16), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n345), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n338), .A2(G125), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n338), .A2(G125), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n349), .B1(new_n350), .B2(new_n340), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n351), .A2(new_n345), .A3(KEYINPUT16), .A4(new_n339), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G146), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(KEYINPUT81), .A3(G146), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n341), .A2(G140), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n349), .A2(new_n359), .A3(new_n199), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n337), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n348), .A2(new_n199), .A3(new_n352), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  OR3_X1    g177(.A1(new_n326), .A2(new_n313), .A3(new_n328), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n363), .B(new_n364), .C1(new_n334), .C2(new_n333), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT22), .B(G137), .ZN(new_n367));
  INV_X1    g181(.A(G953), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n368), .A2(G221), .A3(G234), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n367), .B(new_n369), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n361), .A2(new_n365), .A3(new_n370), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n310), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n372), .A2(KEYINPUT25), .A3(new_n310), .A4(new_n373), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n312), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n311), .A2(G902), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n372), .A2(new_n373), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G214), .B1(G237), .B2(G902), .ZN(new_n384));
  INV_X1    g198(.A(G952), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n385), .A2(KEYINPUT95), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(KEYINPUT95), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n368), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(G234), .B2(G237), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT21), .B(G898), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n391), .B(KEYINPUT96), .Z(new_n392));
  AOI211_X1 g206(.A(new_n310), .B(new_n368), .C1(G234), .C2(G237), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n390), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(G210), .B1(G237), .B2(G902), .ZN(new_n396));
  XOR2_X1   g210(.A(G110), .B(G122), .Z(new_n397));
  INV_X1    g211(.A(G101), .ZN(new_n398));
  INV_X1    g212(.A(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G107), .ZN(new_n400));
  INV_X1    g214(.A(G107), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT3), .A3(G104), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT3), .B1(new_n401), .B2(G104), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n398), .B(new_n400), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT82), .A2(KEYINPUT4), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G101), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(G101), .A3(new_n407), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n243), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n234), .A2(new_n235), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n235), .A2(KEYINPUT5), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n314), .A2(G116), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n415), .B(G113), .C1(KEYINPUT5), .C2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT83), .B1(new_n399), .B2(G107), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n401), .B2(G104), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n401), .A3(G104), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n399), .A2(KEYINPUT84), .A3(G107), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n418), .A2(new_n420), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G101), .ZN(new_n425));
  AND4_X1   g239(.A1(new_n414), .A2(new_n417), .A3(new_n405), .A4(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n397), .B1(new_n413), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n417), .A2(new_n414), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n405), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT3), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n399), .B2(G107), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n433), .A2(new_n402), .B1(new_n399), .B2(G107), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n406), .B1(new_n434), .B2(new_n398), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n398), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n412), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n236), .ZN(new_n438));
  INV_X1    g252(.A(new_n397), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n431), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n224), .A2(new_n341), .ZN(new_n442));
  OAI21_X1  g256(.A(G125), .B1(new_n205), .B2(new_n206), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n442), .B2(new_n443), .ZN(new_n447));
  INV_X1    g261(.A(G224), .ZN(new_n448));
  OAI22_X1  g262(.A1(new_n446), .A2(new_n447), .B1(new_n448), .B2(G953), .ZN(new_n449));
  INV_X1    g263(.A(new_n447), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n448), .A2(G953), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n451), .A3(new_n445), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n454), .B(new_n397), .C1(new_n413), .C2(new_n426), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n441), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n441), .A2(new_n453), .A3(KEYINPUT86), .A4(new_n455), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n397), .B(KEYINPUT8), .Z(new_n461));
  NOR2_X1   g275(.A1(new_n428), .A2(new_n430), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(new_n426), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n442), .A2(new_n443), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT7), .B1(new_n448), .B2(G953), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n463), .A2(new_n440), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n310), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n396), .B1(new_n460), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n396), .ZN(new_n471));
  AOI211_X1 g285(.A(new_n471), .B(new_n468), .C1(new_n458), .C2(new_n459), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n384), .B(new_n395), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G469), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n429), .A2(new_n249), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n224), .B1(new_n425), .B2(new_n405), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n198), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT12), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n207), .A2(new_n213), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n437), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT10), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n225), .B2(new_n227), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n430), .ZN(new_n483));
  INV_X1    g297(.A(new_n198), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n481), .B1(new_n429), .B2(new_n249), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n480), .A2(new_n483), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(G110), .B(G140), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n368), .A2(G227), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n487), .B(new_n488), .Z(new_n489));
  INV_X1    g303(.A(KEYINPUT12), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n490), .B(new_n198), .C1(new_n475), .C2(new_n476), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n478), .A2(new_n486), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n198), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n489), .B1(new_n495), .B2(new_n486), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n474), .B(new_n310), .C1(new_n493), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(G469), .A2(G902), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n478), .A2(new_n486), .A3(new_n491), .ZN(new_n499));
  INV_X1    g313(.A(new_n489), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n486), .A3(new_n489), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(G469), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G221), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT9), .B(G234), .Z(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(new_n310), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  INV_X1    g324(.A(G237), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n368), .A3(G214), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(new_n201), .ZN(new_n513));
  NAND2_X1  g327(.A1(KEYINPUT18), .A2(G131), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n339), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n359), .A2(KEYINPUT78), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n349), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(KEYINPUT87), .B(new_n360), .C1(new_n518), .C2(new_n199), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n351), .A2(new_n339), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT87), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(G146), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n519), .A2(KEYINPUT88), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT88), .B1(new_n519), .B2(new_n522), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n515), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n513), .A2(KEYINPUT89), .A3(G131), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n512), .A2(new_n201), .ZN(new_n528));
  AOI21_X1  g342(.A(G143), .B1(new_n259), .B2(G214), .ZN(new_n529));
  OAI21_X1  g343(.A(G131), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT89), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n513), .A2(G131), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n527), .A2(new_n532), .A3(KEYINPUT17), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n536), .A2(new_n362), .A3(new_n354), .A4(new_n537), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT90), .B(G104), .Z(new_n539));
  XNOR2_X1  g353(.A(G113), .B(G122), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n526), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n343), .A2(new_n350), .A3(KEYINPUT19), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(new_n520), .B2(KEYINPUT19), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n533), .A2(new_n535), .B1(new_n199), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n357), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT81), .B1(new_n353), .B2(G146), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n541), .B1(new_n548), .B2(new_n526), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n510), .B1(new_n542), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT20), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT20), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n552), .B(new_n510), .C1(new_n542), .C2(new_n549), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n541), .B1(new_n526), .B2(new_n538), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n310), .B1(new_n542), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n551), .A2(new_n553), .B1(G475), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(G116), .B(G122), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G107), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n401), .ZN(new_n560));
  XNOR2_X1  g374(.A(G128), .B(G143), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n559), .A2(new_n560), .B1(new_n189), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT91), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT13), .B1(new_n201), .B2(G128), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n201), .A2(G128), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT13), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n219), .B2(G143), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n201), .A2(KEYINPUT13), .A3(G128), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n219), .A2(G143), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT91), .A4(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n566), .A2(new_n571), .A3(G134), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT92), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n566), .A2(new_n571), .A3(KEYINPUT92), .A4(G134), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n562), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n561), .B(new_n189), .ZN(new_n577));
  INV_X1    g391(.A(G116), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(KEYINPUT14), .A3(G122), .ZN(new_n579));
  OAI211_X1 g393(.A(G107), .B(new_n579), .C1(new_n558), .C2(KEYINPUT14), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n580), .A3(new_n560), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n506), .A2(G217), .A3(new_n368), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT93), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n506), .A2(KEYINPUT93), .A3(G217), .A4(new_n368), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n582), .A2(new_n587), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n582), .A2(KEYINPUT94), .A3(new_n587), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(G478), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n594), .A2(KEYINPUT15), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n593), .A2(new_n310), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n595), .B1(new_n593), .B2(new_n310), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n556), .A2(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n473), .A2(new_n509), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n308), .A2(new_n383), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  INV_X1    g416(.A(new_n287), .ZN(new_n603));
  INV_X1    g417(.A(G472), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n285), .B2(new_n310), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n382), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n509), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n585), .A2(KEYINPUT98), .A3(new_n586), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT98), .B1(new_n585), .B2(new_n586), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n582), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT33), .B1(new_n611), .B2(KEYINPUT99), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(KEYINPUT99), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n613), .A2(KEYINPUT100), .A3(new_n591), .A4(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n591), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n616), .B1(new_n617), .B2(new_n612), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n594), .A2(G902), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n593), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT97), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n593), .A2(new_n624), .A3(new_n621), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n619), .A2(new_n620), .A3(new_n623), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n593), .A2(new_n310), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n594), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n555), .A2(G475), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n526), .A2(new_n538), .A3(new_n541), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n548), .A2(new_n526), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n631), .B1(new_n632), .B2(new_n541), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n552), .B1(new_n633), .B2(new_n510), .ZN(new_n634));
  INV_X1    g448(.A(new_n553), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n473), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n606), .A2(new_n607), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n598), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n556), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n473), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n606), .A2(new_n607), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT101), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n645), .B(new_n647), .ZN(G9));
  NOR2_X1   g462(.A1(new_n603), .A2(new_n605), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n371), .A2(KEYINPUT36), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n366), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n361), .A2(new_n365), .A3(new_n651), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n380), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n653), .A2(KEYINPUT102), .A3(new_n380), .A4(new_n654), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n378), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n600), .A2(new_n649), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT103), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n662), .B(new_n664), .ZN(G12));
  OAI21_X1  g479(.A(new_n384), .B1(new_n470), .B2(new_n472), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n389), .B(KEYINPUT104), .Z(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n668), .B2(new_n393), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n556), .A2(new_n642), .A3(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n660), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n308), .A2(new_n672), .A3(new_n607), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n308), .A2(new_n672), .A3(KEYINPUT105), .A4(new_n607), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  NAND2_X1  g492(.A1(new_n460), .A2(new_n469), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n471), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n460), .A2(new_n396), .A3(new_n469), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT38), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n669), .B(new_n685), .Z(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n509), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n660), .B1(new_n689), .B2(KEYINPUT40), .ZN(new_n690));
  INV_X1    g504(.A(new_n384), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n684), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n307), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT32), .B1(new_n285), .B2(new_n286), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n274), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n291), .A2(new_n237), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n696), .B1(new_n263), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n698), .B2(G902), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  AOI211_X1 g514(.A(new_n598), .B(new_n556), .C1(new_n689), .C2(KEYINPUT40), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n692), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  NOR2_X1   g517(.A1(new_n660), .A2(new_n666), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n637), .A2(new_n669), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n308), .A2(new_n607), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  NOR2_X1   g521(.A1(new_n493), .A2(new_n496), .ZN(new_n708));
  OAI21_X1  g522(.A(G469), .B1(new_n708), .B2(G902), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n508), .A3(new_n497), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n709), .A2(KEYINPUT107), .A3(new_n508), .A4(new_n497), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n308), .A2(new_n383), .A3(new_n638), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NOR2_X1   g532(.A1(new_n714), .A2(new_n666), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n308), .A2(new_n719), .A3(new_n383), .A4(new_n644), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NOR2_X1   g535(.A1(new_n660), .A2(new_n599), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n308), .A2(new_n719), .A3(new_n395), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NAND2_X1  g538(.A1(new_n293), .A2(new_n263), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n275), .A2(new_n725), .A3(new_n277), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n726), .A2(new_n286), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n382), .A2(new_n605), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n473), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n636), .B2(new_n642), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n556), .A2(KEYINPUT108), .A3(new_n598), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n728), .A2(new_n729), .A3(new_n715), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  NOR3_X1   g549(.A1(new_n605), .A2(new_n660), .A3(new_n727), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n705), .A3(new_n719), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n680), .A2(new_n384), .A3(new_n681), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n495), .A2(KEYINPUT110), .A3(new_n486), .A4(new_n489), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT110), .B1(new_n499), .B2(new_n500), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n742), .B1(new_n502), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n497), .B1(new_n744), .B2(new_n474), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n498), .B(KEYINPUT109), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n508), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n739), .B1(new_n740), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n470), .A2(new_n472), .A3(new_n691), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n501), .A2(new_n751), .A3(new_n502), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n474), .B1(new_n752), .B2(new_n741), .ZN(new_n753));
  INV_X1    g567(.A(new_n497), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n507), .B1(new_n755), .B2(new_n746), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n750), .A2(new_n756), .A3(KEYINPUT111), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n749), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n308), .A3(new_n383), .A4(new_n705), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n382), .B1(new_n695), .B2(new_n306), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n762), .A2(KEYINPUT42), .A3(new_n705), .A4(new_n758), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  INV_X1    g579(.A(new_n671), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n758), .A2(new_n308), .A3(new_n383), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  INV_X1    g582(.A(new_n629), .ZN(new_n769));
  OR3_X1    g583(.A1(new_n769), .A2(KEYINPUT43), .A3(new_n636), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n556), .A2(KEYINPUT114), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n556), .A2(KEYINPUT114), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n772), .A3(new_n629), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT43), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n649), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n661), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n778), .B1(new_n777), .B2(new_n775), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n750), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT115), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n752), .A2(new_n741), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT45), .ZN(new_n784));
  NAND2_X1  g598(.A1(KEYINPUT45), .A2(G469), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n503), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n503), .A2(KEYINPUT112), .A3(new_n785), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n784), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n746), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT46), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n747), .B1(new_n791), .B2(new_n792), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n754), .B1(new_n797), .B2(KEYINPUT46), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n507), .B(new_n687), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n779), .A2(new_n800), .A3(new_n750), .A4(new_n780), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n782), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  INV_X1    g617(.A(KEYINPUT47), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n796), .A2(new_n798), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n804), .B1(new_n805), .B2(new_n508), .ZN(new_n806));
  AOI211_X1 g620(.A(KEYINPUT47), .B(new_n507), .C1(new_n796), .C2(new_n798), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n308), .A2(new_n383), .A3(new_n740), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n705), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  NAND2_X1  g625(.A1(new_n709), .A2(new_n497), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n773), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n695), .A2(new_n815), .A3(new_n699), .A4(new_n684), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n382), .A2(new_n507), .A3(new_n691), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT116), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n816), .B(new_n818), .C1(new_n814), .C2(new_n813), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n770), .A2(new_n774), .A3(new_n667), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n728), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n812), .A2(new_n508), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n750), .B(new_n822), .C1(new_n808), .C2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n715), .A2(KEYINPUT119), .A3(new_n750), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n714), .B2(new_n740), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n390), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n700), .A2(new_n382), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n556), .A3(new_n769), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n828), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n736), .A3(new_n821), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n728), .A2(new_n715), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n684), .A2(new_n691), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n820), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(KEYINPUT50), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT50), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n820), .A2(new_n834), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n831), .B(new_n833), .C1(new_n837), .C2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n824), .A2(KEYINPUT51), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT51), .B1(new_n824), .B2(new_n841), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n842), .A2(new_n843), .A3(new_n388), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n822), .A2(new_n719), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n706), .A2(new_n737), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n691), .B1(new_n680), .B2(new_n681), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n731), .B2(new_n732), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n695), .B2(new_n699), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n660), .A3(new_n670), .A4(new_n756), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n677), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n734), .A2(new_n716), .A3(new_n720), .A4(new_n723), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n761), .B2(new_n763), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n556), .B1(new_n628), .B2(new_n626), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n729), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT117), .B1(new_n637), .B2(new_n473), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n606), .A2(new_n607), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n645), .A3(new_n601), .A4(new_n662), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n758), .A2(new_n705), .A3(new_n736), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n767), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n660), .A2(new_n740), .A3(new_n599), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n308), .A2(new_n863), .A3(new_n607), .A4(new_n670), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n860), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n677), .A2(new_n846), .A3(new_n850), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n852), .A2(new_n854), .A3(new_n865), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n852), .A2(new_n865), .A3(new_n867), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n853), .A2(KEYINPUT118), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n764), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT53), .B1(new_n853), .B2(KEYINPUT118), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n868), .A2(new_n869), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n844), .A2(new_n845), .A3(new_n872), .A4(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n829), .A2(new_n856), .A3(new_n830), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n832), .A2(new_n762), .A3(new_n821), .ZN(new_n885));
  XNOR2_X1  g699(.A(KEYINPUT120), .B(KEYINPUT48), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n883), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n819), .B1(new_n888), .B2(new_n889), .ZN(G75));
  AOI21_X1  g704(.A(new_n310), .B1(new_n879), .B2(new_n881), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT56), .B1(new_n891), .B2(G210), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n441), .A2(new_n455), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(new_n453), .Z(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT55), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  OR3_X1    g710(.A1(new_n892), .A2(KEYINPUT121), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n368), .A2(G952), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n892), .B2(KEYINPUT121), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n896), .B1(new_n892), .B2(KEYINPUT121), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(G51));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n746), .B(KEYINPUT57), .Z(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n852), .A2(new_n865), .A3(new_n867), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n853), .A2(KEYINPUT118), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n906), .A2(KEYINPUT53), .A3(new_n764), .A4(new_n874), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT54), .B1(new_n870), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n904), .B1(new_n909), .B2(new_n882), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n902), .B1(new_n910), .B2(new_n708), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n903), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n708), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(KEYINPUT122), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n793), .B(KEYINPUT123), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n891), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n911), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n898), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(G54));
  NAND3_X1  g735(.A1(new_n891), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  INV_X1    g736(.A(new_n633), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n898), .ZN(G60));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT59), .Z(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n872), .B2(new_n882), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n619), .A2(new_n623), .A3(new_n625), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n912), .B2(new_n913), .ZN(new_n931));
  OAI221_X1 g745(.A(new_n920), .B1(new_n929), .B2(new_n930), .C1(new_n928), .C2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(G63));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT124), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n870), .B2(new_n908), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n372), .A2(new_n373), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n939), .B(new_n920), .C1(new_n655), .C2(new_n937), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G66));
  INV_X1    g756(.A(new_n392), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n943), .B2(new_n448), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n860), .A2(new_n853), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n944), .B1(new_n945), .B2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n893), .B1(G898), .B2(new_n368), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  NAND2_X1  g762(.A1(new_n637), .A2(new_n643), .ZN(new_n949));
  AND4_X1   g763(.A1(new_n762), .A2(new_n688), .A3(new_n750), .A4(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n677), .A2(new_n846), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n702), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n951), .A2(KEYINPUT62), .A3(new_n702), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n802), .A3(new_n810), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n368), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n268), .B1(new_n272), .B2(new_n269), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT125), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n544), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n368), .A2(G900), .ZN(new_n963));
  AOI211_X1 g777(.A(new_n382), .B(new_n848), .C1(new_n306), .C2(new_n695), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n799), .A2(new_n964), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n764), .A2(new_n810), .A3(new_n767), .A4(new_n965), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n802), .A2(KEYINPUT126), .A3(new_n951), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT126), .B1(new_n802), .B2(new_n951), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n963), .B1(new_n969), .B2(new_n368), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n962), .B1(new_n970), .B2(new_n961), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n368), .B1(G227), .B2(G900), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n972), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n974), .B(new_n962), .C1(new_n970), .C2(new_n961), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(G72));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  INV_X1    g792(.A(new_n945), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n969), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n298), .B(KEYINPUT127), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n980), .A2(new_n263), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n299), .A2(new_n274), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n978), .B(new_n983), .C1(new_n870), .C2(new_n871), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n978), .B1(new_n957), .B2(new_n979), .ZN(new_n985));
  INV_X1    g799(.A(new_n981), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n985), .A2(new_n264), .A3(new_n986), .ZN(new_n987));
  AND4_X1   g801(.A1(new_n920), .A2(new_n982), .A3(new_n984), .A4(new_n987), .ZN(G57));
endmodule


