//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G128), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n196), .A2(KEYINPUT64), .A3(new_n197), .A4(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n189), .A2(KEYINPUT0), .A3(G128), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n191), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT11), .B1(new_n202), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(G137), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G131), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n205), .A2(G134), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(new_n203), .B2(new_n206), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n201), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n217));
  INV_X1    g031(.A(G119), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G116), .ZN(new_n219));
  INV_X1    g033(.A(G116), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT69), .A3(G119), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(G116), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g038(.A(KEYINPUT2), .B(G113), .Z(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n222), .A3(new_n223), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n208), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT66), .B1(new_n202), .B2(G137), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n205), .A3(G134), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n202), .A2(KEYINPUT67), .A3(G137), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n232), .A2(new_n233), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G131), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n193), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n189), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n193), .A2(new_n195), .A3(new_n245), .A4(G128), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n214), .B(new_n238), .C1(new_n244), .C2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n216), .A2(new_n230), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT28), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n216), .A2(new_n251), .A3(new_n230), .A4(new_n248), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n191), .A2(new_n199), .A3(new_n200), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT65), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n191), .A2(new_n199), .A3(new_n256), .A4(new_n200), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n215), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n248), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n229), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n262));
  INV_X1    g076(.A(G237), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G210), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n262), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G101), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT30), .B1(new_n258), .B2(new_n248), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n216), .A2(KEYINPUT30), .A3(new_n248), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n271), .A2(new_n272), .A3(new_n230), .ZN(new_n273));
  INV_X1    g087(.A(new_n249), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n273), .A2(new_n274), .A3(new_n269), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n271), .A2(new_n272), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n274), .B1(new_n278), .B2(new_n229), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n279), .A2(new_n280), .A3(new_n276), .A4(new_n268), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT30), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n259), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n272), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n229), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n285), .A2(new_n276), .A3(new_n249), .A4(new_n268), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT71), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n277), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(G472), .A2(G902), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n187), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n216), .A2(new_n248), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n229), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n253), .A2(KEYINPUT29), .A3(new_n293), .A4(new_n268), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(KEYINPUT72), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n279), .A2(new_n268), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n261), .A2(new_n269), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n298), .A2(KEYINPUT29), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G472), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n287), .A2(new_n281), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n285), .A2(new_n249), .A3(new_n268), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n303), .A2(KEYINPUT31), .B1(new_n269), .B2(new_n261), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n289), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n291), .A2(new_n301), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G217), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(G234), .B2(new_n295), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n312));
  XNOR2_X1  g126(.A(G125), .B(G140), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(new_n313), .B2(KEYINPUT16), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT76), .B1(new_n314), .B2(G146), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G125), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n311), .A2(G140), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT16), .ZN(new_n319));
  OR3_X1    g133(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n192), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n314), .A2(G146), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n315), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n326), .B1(new_n218), .B2(G128), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n239), .A2(G119), .ZN(new_n328));
  MUX2_X1   g142(.A(new_n326), .B(new_n327), .S(new_n328), .Z(new_n329));
  XOR2_X1   g143(.A(KEYINPUT24), .B(G110), .Z(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT23), .B1(new_n239), .B2(G119), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT74), .B1(new_n239), .B2(G119), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n334), .A2(KEYINPUT75), .A3(G110), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT75), .B1(new_n334), .B2(G110), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n325), .B(new_n331), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n324), .A2(KEYINPUT77), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n314), .A2(new_n339), .A3(G146), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n313), .A2(new_n192), .ZN(new_n342));
  OAI22_X1  g156(.A1(G110), .A2(new_n334), .B1(new_n329), .B2(new_n330), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT78), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(KEYINPUT22), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n346), .B(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT22), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n205), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n347), .A2(KEYINPUT22), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n351), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G137), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n345), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n337), .A2(new_n344), .A3(new_n356), .A4(new_n353), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n295), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n358), .A2(KEYINPUT25), .A3(new_n359), .A4(new_n295), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n310), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n358), .A2(new_n359), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n365), .A2(G902), .A3(new_n309), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT79), .B1(new_n364), .B2(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G214), .B1(G237), .B2(G902), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(G210), .B1(G237), .B2(G902), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G107), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(G107), .ZN(new_n378));
  NAND2_X1  g192(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n381));
  OR2_X1    g195(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n382));
  INV_X1    g196(.A(G107), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G104), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n381), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G101), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n379), .B1(new_n378), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G101), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n384), .A2(new_n381), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .A4(new_n377), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n386), .A2(new_n391), .A3(KEYINPUT4), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n393), .B(G101), .C1(new_n380), .C2(new_n385), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n229), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n218), .A3(G116), .ZN(new_n397));
  OAI211_X1 g211(.A(G113), .B(new_n397), .C1(new_n224), .C2(new_n396), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n376), .B2(G107), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n377), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n384), .A2(new_n399), .ZN(new_n402));
  OAI21_X1  g216(.A(G101), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n398), .A2(new_n228), .A3(new_n391), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G122), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n395), .A2(new_n404), .A3(new_n408), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(KEYINPUT6), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n191), .A2(new_n199), .A3(G125), .A4(new_n200), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n244), .A2(new_n247), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(G125), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n264), .A2(G224), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n416), .B(KEYINPUT85), .Z(new_n417));
  XNOR2_X1  g231(.A(new_n415), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n405), .A2(new_n419), .A3(new_n409), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n412), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT86), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT7), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n415), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n416), .A2(KEYINPUT7), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n408), .B(KEYINPUT8), .ZN(new_n427));
  INV_X1    g241(.A(new_n404), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n398), .A2(new_n228), .B1(new_n391), .B2(new_n403), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n415), .A2(KEYINPUT86), .A3(KEYINPUT7), .A4(new_n416), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n426), .A2(new_n430), .A3(new_n411), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n295), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n375), .B1(new_n421), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n412), .A2(new_n418), .A3(new_n420), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n435), .A2(new_n295), .A3(new_n374), .A4(new_n432), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n373), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(G234), .A2(G237), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(G952), .A3(new_n264), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT21), .B(G898), .Z(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(G902), .A3(G953), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G113), .B(G122), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n376), .ZN(new_n449));
  NOR2_X1   g263(.A1(KEYINPUT87), .A2(G143), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n450), .A2(G214), .A3(new_n263), .A4(new_n264), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT87), .B(G143), .ZN(new_n452));
  INV_X1    g266(.A(G214), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n453), .A2(G237), .A3(G953), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n451), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT18), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n455), .B1(new_n456), .B2(new_n213), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n313), .B(new_n192), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n451), .B(G131), .C1(new_n452), .C2(new_n454), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n457), .B(new_n458), .C1(new_n456), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n213), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT17), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(new_n459), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n459), .A2(new_n462), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n449), .B(new_n460), .C1(new_n465), .C2(new_n325), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT90), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n322), .B1(new_n321), .B2(new_n192), .ZN(new_n468));
  AOI211_X1 g282(.A(KEYINPUT76), .B(G146), .C1(new_n319), .C2(new_n320), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n470), .A2(new_n324), .A3(new_n464), .A4(new_n463), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n449), .A4(new_n460), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n461), .A2(new_n459), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n476), .B1(new_n313), .B2(KEYINPUT89), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT19), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT19), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n313), .B2(new_n476), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n478), .B(new_n192), .C1(new_n477), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n341), .A2(new_n475), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n449), .B1(new_n482), .B2(new_n460), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n474), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G475), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n295), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT20), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n220), .A2(G122), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT92), .B1(new_n490), .B2(KEYINPUT14), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n220), .A2(G122), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(KEYINPUT14), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT92), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT14), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n220), .A4(G122), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G107), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n194), .A2(G128), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n239), .A2(G143), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n202), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n202), .B1(new_n500), .B2(new_n501), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n499), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT91), .A3(new_n502), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n492), .A2(new_n490), .A3(new_n383), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n498), .A2(new_n505), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n492), .A2(new_n490), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G107), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n508), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT13), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n501), .B1(new_n500), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT13), .B1(new_n194), .B2(G128), .ZN(new_n515));
  OAI21_X1  g329(.A(G134), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(new_n502), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT9), .B(G234), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n519), .A2(new_n308), .A3(G953), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n509), .A2(new_n517), .A3(new_n520), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n295), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT15), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(G478), .ZN(new_n527));
  INV_X1    g341(.A(G478), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n524), .B(new_n295), .C1(KEYINPUT15), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n449), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n471), .A2(new_n460), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n467), .A2(new_n473), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G475), .B1(new_n534), .B2(G902), .ZN(new_n535));
  AOI21_X1  g349(.A(G475), .B1(new_n474), .B2(new_n484), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(KEYINPUT20), .A3(new_n295), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n489), .A2(new_n531), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(G221), .B1(new_n519), .B2(G902), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT80), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n391), .A2(KEYINPUT10), .A3(new_n403), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n242), .A2(new_n243), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n196), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n246), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n239), .B1(new_n193), .B2(KEYINPUT1), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n246), .B1(new_n546), .B2(new_n189), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n391), .A2(new_n547), .A3(new_n403), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT10), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n542), .A2(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n392), .A2(new_n201), .A3(new_n394), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n215), .ZN(new_n553));
  INV_X1    g367(.A(new_n215), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n554), .A3(new_n551), .ZN(new_n555));
  XNOR2_X1  g369(.A(G110), .B(G140), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n264), .A2(G227), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n391), .A2(new_n547), .A3(new_n403), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n391), .A2(new_n403), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n560), .B1(new_n414), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT83), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n215), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT12), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT12), .ZN(new_n566));
  INV_X1    g380(.A(new_n564), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n414), .A2(new_n561), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n560), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n565), .A2(new_n555), .A3(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(G469), .B(new_n559), .C1(new_n570), .C2(new_n558), .ZN(new_n571));
  INV_X1    g385(.A(G469), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n295), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n558), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n550), .A2(new_n554), .A3(new_n551), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n554), .B1(new_n550), .B2(new_n551), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n565), .A2(new_n555), .A3(new_n569), .A4(new_n558), .ZN(new_n580));
  AOI211_X1 g394(.A(G469), .B(G902), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n541), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n447), .A2(new_n538), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n307), .A2(new_n371), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G101), .ZN(G3));
  AOI21_X1  g399(.A(new_n582), .B1(new_n369), .B2(new_n370), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n305), .A2(new_n295), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(G472), .ZN(new_n589));
  INV_X1    g403(.A(G472), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n305), .B(new_n295), .C1(KEYINPUT93), .C2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n586), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n592), .B(KEYINPUT94), .Z(new_n593));
  NAND3_X1  g407(.A1(new_n489), .A2(new_n535), .A3(new_n537), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n595));
  INV_X1    g409(.A(new_n523), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n520), .B1(new_n509), .B2(new_n517), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n522), .A2(KEYINPUT33), .A3(new_n523), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G478), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n524), .A2(new_n528), .A3(new_n295), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n528), .A2(new_n295), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT95), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n601), .A2(new_n607), .A3(new_n602), .A4(new_n604), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n594), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n593), .A2(new_n447), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT34), .B(G104), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n489), .A2(new_n530), .A3(new_n535), .A4(new_n537), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n373), .B(new_n445), .C1(new_n434), .C2(new_n436), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n447), .A2(KEYINPUT96), .A3(new_n614), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n593), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT35), .B(G107), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  NOR2_X1   g435(.A1(new_n357), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(new_n345), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n295), .A3(new_n310), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n625), .A2(new_n364), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n583), .A2(new_n589), .A3(new_n591), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT37), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n628), .B(G110), .Z(G12));
  AOI21_X1  g443(.A(KEYINPUT20), .B1(new_n536), .B2(new_n295), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n483), .B1(new_n467), .B2(new_n473), .ZN(new_n631));
  NOR4_X1   g445(.A1(new_n631), .A2(new_n488), .A3(G475), .A4(G902), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n533), .A2(new_n532), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n474), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n486), .B1(new_n634), .B2(new_n295), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n630), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n439), .B1(new_n443), .B2(G900), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT97), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n636), .A2(new_n437), .A3(new_n530), .A4(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n615), .A2(KEYINPUT98), .A3(new_n437), .A4(new_n639), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n582), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n644), .A2(new_n307), .A3(new_n645), .A4(new_n626), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  NAND2_X1  g461(.A1(new_n434), .A2(new_n436), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT99), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT38), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n594), .A2(new_n530), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n650), .A2(new_n373), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT32), .B1(new_n305), .B2(new_n289), .ZN(new_n653));
  AOI211_X1 g467(.A(new_n187), .B(new_n290), .C1(new_n302), .C2(new_n304), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n279), .A2(new_n269), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n293), .A2(new_n249), .A3(new_n269), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n295), .ZN(new_n658));
  OAI21_X1  g472(.A(G472), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n638), .B(KEYINPUT39), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n645), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n626), .B1(new_n662), .B2(KEYINPUT40), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n652), .A2(new_n660), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  NAND4_X1  g480(.A1(new_n307), .A2(new_n437), .A3(new_n645), .A4(new_n626), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n606), .A2(new_n608), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n668), .A2(new_n636), .A3(new_n638), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n192), .ZN(G48));
  INV_X1    g486(.A(new_n371), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n655), .B2(new_n301), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n609), .A2(new_n447), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n579), .A2(new_n580), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n572), .B1(new_n676), .B2(new_n295), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n581), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n541), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n674), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NOR2_X1   g497(.A1(new_n618), .A2(new_n617), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n674), .A2(new_n684), .A3(new_n680), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NOR2_X1   g500(.A1(new_n447), .A2(new_n538), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n307), .A2(new_n687), .A3(new_n626), .A4(new_n680), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G119), .ZN(G21));
  NAND2_X1  g503(.A1(new_n587), .A2(G472), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n276), .B1(new_n279), .B2(new_n268), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n268), .B1(new_n253), .B2(new_n293), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT100), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n692), .B1(new_n303), .B2(KEYINPUT31), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT100), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n693), .A2(new_n696), .A3(new_n302), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n289), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n690), .A2(new_n367), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n680), .A2(new_n616), .A3(new_n530), .A4(new_n594), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT101), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n651), .A2(new_n447), .A3(new_n679), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n587), .A2(G472), .B1(new_n697), .B2(new_n289), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .A4(new_n367), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  INV_X1    g521(.A(new_n437), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n679), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n703), .A2(new_n626), .A3(new_n669), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n582), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n434), .A2(new_n372), .A3(new_n436), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  OAI211_X1 g529(.A(KEYINPUT102), .B(new_n541), .C1(new_n575), .C2(new_n581), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT103), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n713), .A2(new_n719), .A3(new_n715), .A4(new_n716), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n307), .A2(KEYINPUT104), .A3(new_n367), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT104), .B1(new_n307), .B2(new_n367), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n669), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n307), .A2(new_n371), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n720), .B2(new_n718), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n670), .A2(KEYINPUT42), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n724), .A2(KEYINPUT42), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  NOR2_X1   g543(.A1(new_n614), .A2(new_n638), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n721), .A2(new_n674), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT106), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  OAI21_X1  g549(.A(new_n559), .B1(new_n570), .B2(new_n558), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT45), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n737), .A2(G469), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT107), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(KEYINPUT107), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n573), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n742));
  INV_X1    g556(.A(new_n581), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n741), .B2(KEYINPUT46), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n541), .B(new_n661), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n668), .A2(new_n594), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT43), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n589), .A2(new_n591), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n626), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n746), .A2(new_n715), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT108), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n205), .ZN(G39));
  OAI21_X1  g570(.A(new_n541), .B1(new_n742), .B2(new_n744), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT47), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n307), .A2(new_n670), .A3(new_n371), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n760), .B(new_n541), .C1(new_n742), .C2(new_n744), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(new_n715), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G140), .ZN(G42));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n646), .B(new_n710), .C1(new_n670), .C2(new_n667), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n626), .A2(new_n638), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n651), .A2(new_n708), .A3(new_n582), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n660), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n764), .B1(new_n765), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n538), .A2(new_n714), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n773), .B1(new_n774), .B2(new_n639), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n538), .A2(new_n714), .A3(KEYINPUT112), .A4(new_n638), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n307), .A3(new_n645), .A4(new_n626), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n626), .A2(new_n669), .A3(new_n690), .A4(new_n698), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n721), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n733), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT113), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n733), .A2(new_n778), .A3(new_n780), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n447), .B1(new_n609), .B2(new_n614), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n591), .A3(new_n589), .A4(new_n586), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n584), .A2(new_n787), .A3(new_n627), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n584), .A2(new_n787), .A3(new_n627), .A4(KEYINPUT111), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n706), .A2(new_n681), .A3(new_n685), .A4(new_n688), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n772), .A2(new_n785), .A3(new_n728), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n770), .A2(new_n771), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT53), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n794), .A2(new_n728), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n646), .A2(new_n710), .ZN(new_n800));
  INV_X1    g614(.A(new_n671), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n800), .A2(new_n801), .A3(new_n771), .A4(new_n768), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT52), .B1(new_n765), .B2(new_n769), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n798), .A2(new_n799), .A3(new_n785), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n797), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n798), .A2(new_n785), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(KEYINPUT53), .A3(new_n804), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n799), .B1(new_n795), .B2(new_n796), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n810), .A2(KEYINPUT115), .A3(KEYINPUT53), .A4(new_n804), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n809), .B1(new_n816), .B2(KEYINPUT54), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n748), .A2(new_n440), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n818), .A2(new_n367), .A3(new_n703), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n709), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n758), .A2(new_n761), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n677), .A2(new_n581), .A3(new_n541), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n715), .B(new_n819), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n679), .A2(new_n714), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n626), .A3(new_n703), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n819), .A2(new_n373), .A3(new_n650), .A4(new_n680), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT50), .Z(new_n828));
  NAND2_X1  g642(.A1(new_n824), .A2(new_n371), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n660), .A2(new_n829), .A3(new_n439), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n636), .A3(new_n668), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n823), .A2(new_n826), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT51), .ZN(new_n833));
  INV_X1    g647(.A(new_n609), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(G952), .A3(new_n264), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n722), .A2(new_n723), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n825), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n817), .A2(new_n820), .A3(new_n833), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(G952), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n264), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT49), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n367), .B(new_n541), .C1(new_n678), .C2(new_n847), .ZN(new_n848));
  NOR4_X1   g662(.A1(new_n848), .A2(new_n373), .A3(new_n594), .A4(new_n668), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT109), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n849), .A2(new_n850), .B1(new_n847), .B2(new_n678), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  INV_X1    g666(.A(new_n650), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n852), .A2(new_n853), .A3(new_n660), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT110), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n846), .A2(new_n855), .ZN(G75));
  NOR2_X1   g670(.A1(new_n806), .A2(new_n295), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT56), .B1(new_n857), .B2(G210), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n412), .A2(new_n420), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(new_n418), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT55), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n858), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n844), .A2(G953), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT117), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n862), .A2(new_n865), .ZN(G51));
  NAND3_X1  g680(.A1(new_n797), .A2(KEYINPUT54), .A3(new_n805), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n797), .A2(KEYINPUT118), .A3(new_n805), .A4(KEYINPUT54), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n808), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n573), .B(KEYINPUT57), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT119), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n871), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n676), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n857), .A2(new_n739), .A3(new_n740), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n865), .B1(new_n877), .B2(new_n878), .ZN(G54));
  NAND2_X1  g693(.A1(new_n857), .A2(KEYINPUT58), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n880), .A2(new_n486), .A3(new_n631), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n631), .B1(new_n880), .B2(new_n486), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(KEYINPUT120), .B(new_n631), .C1(new_n880), .C2(new_n486), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n865), .B(new_n881), .C1(new_n884), .C2(new_n885), .ZN(G60));
  XNOR2_X1  g700(.A(new_n603), .B(KEYINPUT59), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n600), .B1(new_n817), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n887), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n871), .A2(new_n598), .A3(new_n599), .A4(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n888), .A2(new_n864), .A3(new_n890), .ZN(G63));
  NAND2_X1  g705(.A1(G217), .A2(G902), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT60), .Z(new_n893));
  NAND3_X1  g707(.A1(new_n797), .A2(new_n805), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n365), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n797), .A2(new_n623), .A3(new_n805), .A4(new_n893), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n864), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT61), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n897), .B(new_n899), .ZN(G66));
  INV_X1    g714(.A(G224), .ZN(new_n901));
  OAI21_X1  g715(.A(G953), .B1(new_n442), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n794), .B2(G953), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n859), .B1(G898), .B2(new_n264), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT122), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n903), .B(new_n905), .ZN(G69));
  OAI21_X1  g720(.A(new_n478), .B1(new_n477), .B2(new_n480), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n278), .B(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(G227), .B1(new_n909), .B2(KEYINPUT125), .ZN(new_n910));
  INV_X1    g724(.A(G900), .ZN(new_n911));
  OAI21_X1  g725(.A(G953), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n754), .A2(new_n762), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n651), .A2(new_n708), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n746), .A2(new_n837), .A3(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n915), .A2(new_n728), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n765), .B(KEYINPUT123), .Z(new_n917));
  AND2_X1   g731(.A1(new_n917), .A2(new_n733), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n913), .A2(new_n916), .A3(new_n264), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(G900), .A2(G953), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n919), .A2(new_n909), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n917), .A2(new_n665), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n923), .B2(KEYINPUT62), .ZN(new_n924));
  XOR2_X1   g738(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n925));
  NAND3_X1  g739(.A1(new_n917), .A2(new_n665), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n725), .B1(new_n609), .B2(new_n614), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n927), .A2(new_n645), .A3(new_n661), .A4(new_n715), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n913), .A2(new_n924), .A3(new_n926), .A4(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n909), .B1(new_n929), .B2(new_n264), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n921), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n912), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n932), .B(new_n912), .C1(new_n921), .C2(new_n930), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n933), .A2(new_n935), .ZN(G72));
  NAND2_X1  g750(.A1(G472), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT63), .Z(new_n938));
  NAND3_X1  g752(.A1(new_n913), .A2(new_n918), .A3(new_n916), .ZN(new_n939));
  INV_X1    g753(.A(new_n794), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n941), .A2(KEYINPUT127), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n279), .A2(new_n269), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n941), .B2(KEYINPUT127), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n865), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n938), .B1(new_n929), .B2(new_n940), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT126), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n948), .B(new_n938), .C1(new_n929), .C2(new_n940), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n656), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n656), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n816), .A2(new_n951), .A3(new_n938), .A4(new_n943), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n945), .A2(new_n950), .A3(new_n952), .ZN(G57));
endmodule


