//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT24), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n205), .A2(G183gat), .A3(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n212), .A2(new_n213), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT64), .B1(new_n218), .B2(KEYINPUT23), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n214), .A2(new_n220), .A3(new_n216), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n211), .B(new_n217), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n207), .B1(new_n228), .B2(G183gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n218), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(KEYINPUT23), .A3(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n229), .A2(KEYINPUT25), .A3(new_n233), .A4(new_n217), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n224), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n208), .A2(KEYINPUT27), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT27), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G183gat), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n225), .A2(new_n227), .A3(new_n236), .A4(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT28), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT67), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n239), .A2(new_n243), .A3(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n236), .A2(new_n238), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n228), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n236), .A2(new_n238), .A3(KEYINPUT68), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT28), .A4(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n242), .A2(new_n244), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT26), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n230), .A2(new_n252), .A3(new_n232), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n215), .B1(KEYINPUT26), .B2(new_n214), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n253), .A2(new_n254), .B1(G183gat), .B2(G190gat), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n251), .A2(KEYINPUT69), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT69), .B1(new_n251), .B2(new_n255), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n235), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G120gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(G113gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT70), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(new_n259), .B2(G113gat), .ZN(new_n263));
  INV_X1    g062(.A(G113gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n261), .B(new_n263), .C1(new_n264), .C2(G120gat), .ZN(new_n265));
  XOR2_X1   g064(.A(G127gat), .B(G134gat), .Z(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n264), .A2(G120gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n269), .B1(new_n270), .B2(new_n260), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n266), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT71), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n265), .A2(new_n267), .B1(new_n271), .B2(new_n266), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n258), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G227gat), .A2(G233gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n278), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n281), .B(new_n235), .C1(new_n257), .C2(new_n256), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT34), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT34), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n279), .A2(new_n282), .A3(new_n285), .A4(new_n280), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n202), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G15gat), .B(G43gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT72), .ZN(new_n290));
  XOR2_X1   g089(.A(G71gat), .B(G99gat), .Z(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n280), .B1(new_n279), .B2(new_n282), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(KEYINPUT33), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT32), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n294), .A2(new_n296), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n288), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n294), .A2(new_n296), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n296), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(new_n287), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT36), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n284), .B(new_n286), .C1(new_n297), .C2(new_n298), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n284), .A2(new_n286), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(new_n301), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G155gat), .ZN(new_n310));
  INV_X1    g109(.A(G162gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G141gat), .B(G148gat), .Z(new_n315));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G141gat), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT80), .B1(new_n319), .B2(G148gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT80), .ZN(new_n321));
  INV_X1    g120(.A(G148gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n322), .A3(G141gat), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n320), .B(new_n323), .C1(G141gat), .C2(new_n322), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n313), .B1(new_n312), .B2(KEYINPUT2), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(KEYINPUT81), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT81), .B1(new_n324), .B2(new_n325), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n318), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n275), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n324), .A2(new_n325), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n317), .B1(new_n333), .B2(new_n326), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G225gat), .A2(G233gat), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n274), .A2(new_n334), .A3(new_n277), .A4(KEYINPUT4), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n275), .B(new_n318), .C1(new_n328), .C2(new_n327), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n337), .A2(new_n338), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT5), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n273), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n340), .ZN(new_n346));
  INV_X1    g145(.A(new_n338), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n347), .B1(new_n330), .B2(new_n336), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n274), .A2(new_n334), .A3(new_n277), .A4(new_n341), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n340), .A2(KEYINPUT4), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT82), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT82), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n340), .A2(new_n354), .A3(KEYINPUT4), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n350), .A2(new_n353), .A3(new_n344), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT0), .ZN(new_n359));
  XNOR2_X1  g158(.A(G57gat), .B(G85gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(KEYINPUT6), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n349), .A2(new_n361), .A3(new_n356), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n357), .A2(new_n362), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n365), .B1(new_n364), .B2(new_n366), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n363), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n372));
  XNOR2_X1  g171(.A(G197gat), .B(G204gat), .ZN(new_n373));
  INV_X1    g172(.A(G211gat), .ZN(new_n374));
  INV_X1    g173(.A(G218gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(KEYINPUT22), .B2(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(G211gat), .B(G218gat), .Z(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n258), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n251), .A2(new_n255), .B1(new_n224), .B2(new_n234), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n385), .B1(new_n386), .B2(new_n381), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n251), .A2(new_n255), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n235), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n389), .A2(KEYINPUT75), .A3(new_n382), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n380), .B1(new_n384), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n258), .A2(new_n382), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n388), .B2(new_n235), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT76), .B1(new_n394), .B2(new_n382), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n396), .B(new_n381), .C1(new_n386), .C2(KEYINPUT29), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n393), .A2(new_n395), .A3(new_n379), .A4(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n372), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G8gat), .B(G36gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n392), .A2(new_n372), .A3(new_n398), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n400), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n405), .A3(new_n398), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n371), .A2(new_n408), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT84), .B(G22gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT31), .B(G50gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G78gat), .B(G106gat), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n379), .B1(new_n336), .B2(new_n383), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n379), .A2(new_n383), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n334), .B1(new_n420), .B2(new_n335), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n418), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n419), .A2(new_n421), .A3(new_n418), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n417), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G228gat), .A2(G233gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n419), .A2(new_n421), .ZN(new_n427));
  INV_X1    g226(.A(new_n418), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(new_n416), .A3(new_n422), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n426), .B1(new_n425), .B2(new_n430), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n415), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n433), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(new_n414), .A3(new_n431), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n304), .A2(new_n309), .B1(new_n413), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n364), .A2(new_n366), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n361), .B(KEYINPUT85), .Z(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n349), .B2(new_n356), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n363), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n410), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT37), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n392), .A2(new_n444), .A3(new_n398), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n379), .B1(new_n384), .B2(new_n391), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n393), .A2(new_n395), .A3(new_n380), .A4(new_n397), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(KEYINPUT37), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n405), .A2(KEYINPUT38), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n392), .A2(new_n372), .A3(new_n398), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n452), .A2(new_n399), .A3(new_n444), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT86), .B1(new_n453), .B2(new_n405), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n400), .A2(KEYINPUT37), .A3(new_n407), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n406), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n457), .A3(new_n445), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n451), .B1(new_n458), .B2(KEYINPUT38), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n434), .A2(new_n436), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n411), .A2(new_n408), .A3(new_n412), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n353), .A2(new_n337), .A3(new_n355), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n347), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n464), .B(KEYINPUT39), .C1(new_n347), .C2(new_n346), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n465), .B(new_n440), .C1(KEYINPUT39), .C2(new_n464), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT40), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n441), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n467), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n460), .B1(new_n462), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n438), .B1(new_n459), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n303), .A2(new_n460), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT35), .B1(new_n472), .B2(new_n413), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT35), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n460), .A2(new_n474), .A3(new_n442), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n305), .A2(new_n307), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n462), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n473), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT87), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n471), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n484));
  INV_X1    g283(.A(G36gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n486), .A2(KEYINPUT92), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(KEYINPUT92), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT91), .B(G29gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(new_n485), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT93), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n494), .B2(new_n485), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n490), .A2(new_n493), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n488), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n488), .A2(new_n500), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n501), .A2(new_n502), .A3(new_n486), .ZN(new_n503));
  OAI211_X1 g302(.A(KEYINPUT15), .B(new_n491), .C1(new_n503), .C2(new_n495), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT16), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(G1gat), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(G1gat), .B2(new_n507), .ZN(new_n510));
  INV_X1    g309(.A(G8gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n506), .A2(KEYINPUT17), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n514), .A2(new_n512), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n506), .A2(KEYINPUT17), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT18), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(KEYINPUT18), .A3(new_n518), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n505), .B(new_n512), .Z(new_n523));
  XOR2_X1   g322(.A(new_n518), .B(KEYINPUT13), .Z(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT89), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(new_n264), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(new_n319), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n529), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT12), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n526), .B(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(G71gat), .A2(G78gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(G71gat), .A2(G78gat), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(KEYINPUT9), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G57gat), .ZN(new_n538));
  INV_X1    g337(.A(G64gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G57gat), .A2(G64gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT95), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544));
  AND2_X1   g343(.A1(G57gat), .A2(G64gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(G57gat), .A2(G64gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n536), .A2(KEYINPUT9), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n544), .B(new_n547), .C1(new_n548), .C2(new_n535), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT94), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n545), .B2(new_n546), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n540), .A2(KEYINPUT94), .A3(new_n541), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT9), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n535), .A2(new_n536), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n543), .A2(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(KEYINPUT97), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n561));
  AND2_X1   g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(new_n557), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT7), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(G85gat), .A3(G92gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G85gat), .ZN(new_n570));
  INV_X1    g369(.A(G92gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(KEYINPUT8), .A2(new_n559), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n564), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n560), .A2(new_n563), .A3(new_n569), .A4(new_n572), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT10), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n556), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT99), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n573), .A2(KEYINPUT98), .A3(new_n563), .A4(new_n560), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT98), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n569), .B(new_n572), .C1(new_n564), .C2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n555), .A2(new_n580), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n555), .A2(new_n581), .A3(new_n583), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT99), .B1(new_n555), .B2(new_n576), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n579), .B1(new_n587), .B2(new_n578), .ZN(new_n588));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n587), .A2(new_n589), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n599), .B1(new_n591), .B2(new_n593), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n534), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n555), .A2(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n606), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G183gat), .B(G211gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT21), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n512), .B1(new_n612), .B2(new_n556), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n516), .A2(new_n514), .A3(new_n577), .ZN(new_n620));
  AND2_X1   g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n505), .A2(new_n576), .B1(KEYINPUT41), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n603), .A2(new_n619), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n483), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n483), .A2(KEYINPUT100), .A3(new_n633), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n371), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g440(.A(KEYINPUT101), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G8gat), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(new_n461), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n511), .B1(new_n638), .B2(new_n461), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT42), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT42), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(G1325gat));
  INV_X1    g449(.A(new_n476), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(G15gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n638), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(G15gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n304), .A2(new_n309), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n655), .B1(new_n636), .B2(new_n637), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n653), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT102), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n653), .B(new_n659), .C1(new_n654), .C2(new_n656), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(G1326gat));
  NAND2_X1  g460(.A1(new_n638), .A2(new_n437), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT43), .B(G22gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  INV_X1    g463(.A(new_n533), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n526), .B(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n480), .B2(new_n482), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n619), .A2(new_n632), .A3(new_n602), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n667), .A2(new_n639), .A3(new_n494), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT45), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n631), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n471), .A2(new_n481), .A3(new_n478), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n481), .B1(new_n471), .B2(new_n478), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n479), .A2(new_n632), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n672), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n618), .B(KEYINPUT103), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n603), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n371), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n671), .B1(new_n494), .B2(new_n684), .ZN(G1328gat));
  NAND4_X1  g484(.A1(new_n667), .A2(new_n485), .A3(new_n461), .A4(new_n669), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT46), .Z(new_n687));
  OAI21_X1  g486(.A(G36gat), .B1(new_n683), .B2(new_n462), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(G1329gat));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT47), .ZN(new_n691));
  INV_X1    g490(.A(new_n655), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n676), .A2(new_n692), .A3(new_n678), .A4(new_n682), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n668), .A2(new_n651), .A3(G43gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n693), .A2(G43gat), .B1(new_n667), .B2(new_n695), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n690), .B(new_n691), .C1(new_n696), .C2(KEYINPUT104), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n693), .A2(G43gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n667), .A2(new_n695), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT105), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT47), .B1(new_n696), .B2(new_n690), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n697), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(G1330gat));
  NAND3_X1  g504(.A1(new_n667), .A2(new_n437), .A3(new_n669), .ZN(new_n706));
  INV_X1    g505(.A(G50gat), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n706), .A2(new_n707), .B1(new_n708), .B2(KEYINPUT48), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n437), .A2(G50gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n683), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n708), .A2(KEYINPUT48), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n711), .B(new_n713), .ZN(G1331gat));
  NAND3_X1  g513(.A1(new_n666), .A2(new_n618), .A3(new_n631), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n602), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT107), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n717), .A2(new_n479), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n639), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g519(.A(new_n462), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT108), .Z(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n723), .B(new_n724), .Z(G1333gat));
  NAND2_X1  g524(.A1(new_n718), .A2(new_n692), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n651), .A2(G71gat), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n726), .A2(G71gat), .B1(new_n718), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n718), .A2(new_n437), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g530(.A1(new_n534), .A2(new_n602), .A3(new_n618), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n679), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n371), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n631), .B1(new_n471), .B2(new_n478), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n534), .A2(new_n618), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(KEYINPUT51), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n735), .A2(new_n736), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n739), .A2(new_n740), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n602), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n745), .B2(new_n744), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n639), .A2(new_n570), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n734), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  NAND3_X1  g548(.A1(new_n679), .A2(new_n461), .A3(new_n732), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G92gat), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n462), .A2(G92gat), .A3(new_n602), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n744), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n743), .A2(new_n737), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n750), .A2(G92gat), .B1(new_n756), .B2(new_n754), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n753), .A2(new_n755), .B1(new_n757), .B2(new_n752), .ZN(G1337gat));
  OR2_X1    g557(.A1(new_n651), .A2(G99gat), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n733), .B2(new_n655), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G99gat), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n733), .A2(new_n760), .A3(new_n655), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n747), .A2(new_n759), .B1(new_n762), .B2(new_n763), .ZN(G1338gat));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n460), .A2(G106gat), .A3(new_n602), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n744), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n765), .B1(new_n744), .B2(new_n766), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n676), .A2(new_n437), .A3(new_n678), .A4(new_n732), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT113), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G106gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n771), .A2(KEYINPUT113), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n771), .A2(G106gat), .B1(new_n756), .B2(new_n766), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n769), .A2(new_n775), .B1(new_n770), .B2(new_n776), .ZN(G1339gat));
  NAND2_X1  g576(.A1(new_n526), .A2(new_n533), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n517), .A2(new_n518), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n523), .A2(new_n524), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n532), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n601), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n598), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n597), .B1(new_n591), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n587), .A2(new_n578), .ZN(new_n787));
  INV_X1    g586(.A(new_n579), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n784), .B1(new_n789), .B2(new_n589), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n588), .A2(KEYINPUT114), .A3(new_n590), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(new_n590), .A3(new_n788), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n790), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n790), .A2(new_n794), .A3(KEYINPUT115), .A4(new_n791), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n786), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n783), .B1(new_n799), .B2(KEYINPUT55), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT54), .B1(new_n588), .B2(new_n590), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT114), .B1(new_n588), .B2(new_n590), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT115), .B1(new_n803), .B2(new_n791), .ZN(new_n804));
  INV_X1    g603(.A(new_n798), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n785), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n800), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n782), .B1(new_n809), .B2(new_n666), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n631), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n778), .A2(new_n781), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n809), .A2(new_n631), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n680), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n715), .A2(new_n601), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n461), .A2(new_n371), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n472), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(G113gat), .B1(new_n823), .B2(new_n534), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n437), .B1(new_n815), .B2(new_n817), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n820), .A2(new_n651), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n666), .A2(new_n264), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(G1340gat));
  AOI21_X1  g628(.A(G120gat), .B1(new_n823), .B2(new_n601), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n602), .A2(new_n259), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n827), .B2(new_n831), .ZN(G1341gat));
  INV_X1    g631(.A(new_n827), .ZN(new_n833));
  OAI21_X1  g632(.A(G127gat), .B1(new_n833), .B2(new_n680), .ZN(new_n834));
  INV_X1    g633(.A(G127gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n823), .A2(new_n835), .A3(new_n618), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(G1342gat));
  OR2_X1    g636(.A1(new_n631), .A2(G134gat), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n822), .A2(new_n838), .B1(new_n839), .B2(KEYINPUT56), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n840), .B(new_n841), .Z(new_n842));
  OAI21_X1  g641(.A(G134gat), .B1(new_n833), .B2(new_n631), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(G1343gat));
  NOR2_X1   g646(.A1(new_n692), .A2(new_n460), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n819), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n815), .B2(new_n817), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n534), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n319), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n655), .A2(new_n819), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n460), .B1(new_n815), .B2(new_n817), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(KEYINPUT55), .B(new_n785), .C1(new_n804), .C2(new_n805), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n598), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n799), .A2(KEYINPUT55), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT118), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n800), .A2(new_n861), .A3(new_n808), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n534), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n632), .B1(new_n863), .B2(new_n782), .ZN(new_n864));
  INV_X1    g663(.A(new_n813), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n619), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n460), .B1(new_n866), .B2(new_n817), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n856), .B1(new_n855), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n534), .A2(G141gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n852), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT119), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT58), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n870), .A2(KEYINPUT119), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1344gat));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n876), .B(G148gat), .C1(new_n868), .C2(new_n602), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n681), .B1(new_n811), .B2(new_n813), .ZN(new_n878));
  OAI211_X1 g677(.A(KEYINPUT57), .B(new_n437), .C1(new_n878), .C2(new_n816), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n867), .B2(KEYINPUT57), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n655), .A2(new_n601), .A3(new_n819), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n322), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n877), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n850), .A2(new_n322), .A3(new_n601), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1345gat));
  OAI21_X1  g685(.A(G155gat), .B1(new_n868), .B2(new_n680), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n850), .A2(new_n310), .A3(new_n618), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(KEYINPUT120), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1346gat));
  OAI21_X1  g692(.A(G162gat), .B1(new_n868), .B2(new_n631), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n850), .A2(new_n311), .A3(new_n632), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n462), .A2(new_n639), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT122), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n898), .A2(new_n476), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n825), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(new_n212), .A3(new_n666), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n818), .A2(new_n897), .ZN(new_n902));
  INV_X1    g701(.A(new_n472), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n534), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n901), .B1(new_n907), .B2(new_n212), .ZN(G1348gat));
  OAI21_X1  g707(.A(G176gat), .B1(new_n900), .B2(new_n602), .ZN(new_n909));
  INV_X1    g708(.A(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n601), .A2(new_n213), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(G1349gat));
  INV_X1    g711(.A(new_n904), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n913), .A2(new_n247), .A3(new_n249), .A4(new_n618), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(new_n900), .B2(new_n680), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n825), .A2(KEYINPUT123), .A3(new_n681), .A4(new_n899), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(G183gat), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT60), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n914), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1350gat));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n248), .A3(new_n632), .ZN(new_n924));
  OAI21_X1  g723(.A(G190gat), .B1(new_n900), .B2(new_n631), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(KEYINPUT61), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(KEYINPUT61), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G1351gat));
  AND2_X1   g727(.A1(new_n902), .A2(new_n848), .ZN(new_n929));
  AOI21_X1  g728(.A(G197gat), .B1(new_n929), .B2(new_n534), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n898), .A2(new_n655), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT125), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n880), .A2(KEYINPUT124), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n935), .B(new_n879), .C1(new_n867), .C2(KEYINPUT57), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n534), .A2(G197gat), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n930), .B1(new_n937), .B2(new_n938), .ZN(G1352gat));
  INV_X1    g738(.A(new_n782), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n666), .B1(new_n809), .B2(KEYINPUT118), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n862), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n813), .B1(new_n942), .B2(new_n632), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n816), .B1(new_n943), .B2(new_n619), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n855), .B1(new_n944), .B2(new_n460), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n935), .B1(new_n945), .B2(new_n879), .ZN(new_n946));
  INV_X1    g745(.A(new_n936), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n932), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(G204gat), .B1(new_n948), .B2(new_n602), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n602), .A2(G204gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n902), .A2(new_n848), .A3(new_n950), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT62), .Z(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(new_n952), .ZN(G1353gat));
  NOR2_X1   g752(.A1(new_n931), .A2(new_n619), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n374), .B1(new_n880), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT63), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n929), .A2(new_n374), .A3(new_n618), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1354gat));
  NAND4_X1  g757(.A1(new_n818), .A2(new_n632), .A3(new_n848), .A4(new_n897), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(new_n375), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT126), .Z(new_n961));
  NAND2_X1  g760(.A1(new_n632), .A2(G218gat), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n937), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n948), .A2(KEYINPUT127), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(G1355gat));
endmodule


