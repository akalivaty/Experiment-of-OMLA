

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(G1384), .A2(n772), .ZN(n614) );
  OR2_X1 U553 ( .A1(n646), .A2(n933), .ZN(n645) );
  NOR2_X1 U554 ( .A1(n615), .A2(n745), .ZN(n617) );
  NAND2_X1 U555 ( .A1(n614), .A2(n613), .ZN(n615) );
  BUF_X1 U556 ( .A(n772), .Z(G164) );
  INV_X1 U557 ( .A(KEYINPUT64), .ZN(n633) );
  INV_X1 U558 ( .A(n688), .ZN(n672) );
  AND2_X1 U559 ( .A1(n699), .A2(n698), .ZN(n701) );
  XNOR2_X1 U560 ( .A(n537), .B(KEYINPUT17), .ZN(n598) );
  INV_X1 U561 ( .A(G2104), .ZN(n536) );
  BUF_X1 U562 ( .A(n598), .Z(n905) );
  NOR2_X2 U563 ( .A1(n564), .A2(n525), .ZN(n621) );
  OR2_X1 U564 ( .A1(n724), .A2(n723), .ZN(n520) );
  INV_X1 U565 ( .A(KEYINPUT26), .ZN(n616) );
  INV_X1 U566 ( .A(KEYINPUT93), .ZN(n651) );
  XNOR2_X1 U567 ( .A(n651), .B(KEYINPUT27), .ZN(n652) );
  XNOR2_X1 U568 ( .A(n653), .B(n652), .ZN(n656) );
  INV_X1 U569 ( .A(KEYINPUT95), .ZN(n649) );
  XNOR2_X1 U570 ( .A(n678), .B(KEYINPUT30), .ZN(n679) );
  INV_X1 U571 ( .A(KEYINPUT96), .ZN(n680) );
  INV_X1 U572 ( .A(KEYINPUT29), .ZN(n669) );
  INV_X1 U573 ( .A(KEYINPUT97), .ZN(n700) );
  INV_X1 U574 ( .A(KEYINPUT99), .ZN(n707) );
  BUF_X1 U575 ( .A(n615), .Z(n688) );
  NAND2_X1 U576 ( .A1(G8), .A2(n688), .ZN(n724) );
  AND2_X1 U577 ( .A1(n725), .A2(n520), .ZN(n726) );
  INV_X1 U578 ( .A(KEYINPUT100), .ZN(n728) );
  INV_X1 U579 ( .A(G2105), .ZN(n535) );
  XNOR2_X1 U580 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U581 ( .A(KEYINPUT13), .B(KEYINPUT68), .ZN(n626) );
  NOR2_X2 U582 ( .A1(G651), .A2(G543), .ZN(n794) );
  XNOR2_X1 U583 ( .A(n627), .B(n626), .ZN(n628) );
  BUF_X1 U584 ( .A(n599), .Z(n906) );
  AND2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n909) );
  NOR2_X1 U586 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U587 ( .A1(n631), .A2(n630), .ZN(n946) );
  AND2_X1 U588 ( .A1(n543), .A2(n542), .ZN(G160) );
  NAND2_X1 U589 ( .A1(n794), .A2(G89), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n521), .B(KEYINPUT4), .ZN(n523) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n564) );
  INV_X1 U592 ( .A(G651), .ZN(n525) );
  NAND2_X1 U593 ( .A1(G76), .A2(n621), .ZN(n522) );
  NAND2_X1 U594 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U595 ( .A(n524), .B(KEYINPUT5), .ZN(n531) );
  NOR2_X1 U596 ( .A1(G543), .A2(n525), .ZN(n526) );
  XOR2_X2 U597 ( .A(KEYINPUT1), .B(n526), .Z(n793) );
  NAND2_X1 U598 ( .A1(G63), .A2(n793), .ZN(n528) );
  NOR2_X2 U599 ( .A1(G651), .A2(n564), .ZN(n791) );
  NAND2_X1 U600 ( .A1(G51), .A2(n791), .ZN(n527) );
  NAND2_X1 U601 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U602 ( .A(KEYINPUT6), .B(n529), .Z(n530) );
  NAND2_X1 U603 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U604 ( .A(n532), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U605 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U606 ( .A1(n535), .A2(G2104), .ZN(n533) );
  XNOR2_X2 U607 ( .A(n533), .B(KEYINPUT65), .ZN(n599) );
  NAND2_X1 U608 ( .A1(G101), .A2(n599), .ZN(n534) );
  XOR2_X1 U609 ( .A(n534), .B(KEYINPUT23), .Z(n543) );
  NAND2_X1 U610 ( .A1(n536), .A2(n535), .ZN(n537) );
  AND2_X1 U611 ( .A1(n598), .A2(G137), .ZN(n541) );
  NAND2_X1 U612 ( .A1(G113), .A2(n909), .ZN(n539) );
  NOR2_X1 U613 ( .A1(G2104), .A2(n535), .ZN(n600) );
  NAND2_X1 U614 ( .A1(G125), .A2(n600), .ZN(n538) );
  NAND2_X1 U615 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U616 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U617 ( .A1(G72), .A2(n621), .ZN(n545) );
  NAND2_X1 U618 ( .A1(G85), .A2(n794), .ZN(n544) );
  NAND2_X1 U619 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U620 ( .A1(G60), .A2(n793), .ZN(n547) );
  NAND2_X1 U621 ( .A1(G47), .A2(n791), .ZN(n546) );
  NAND2_X1 U622 ( .A1(n547), .A2(n546), .ZN(n548) );
  OR2_X1 U623 ( .A1(n549), .A2(n548), .ZN(G290) );
  NAND2_X1 U624 ( .A1(G64), .A2(n793), .ZN(n551) );
  NAND2_X1 U625 ( .A1(G52), .A2(n791), .ZN(n550) );
  NAND2_X1 U626 ( .A1(n551), .A2(n550), .ZN(n556) );
  NAND2_X1 U627 ( .A1(G77), .A2(n621), .ZN(n553) );
  NAND2_X1 U628 ( .A1(G90), .A2(n794), .ZN(n552) );
  NAND2_X1 U629 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U630 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U631 ( .A1(n556), .A2(n555), .ZN(G171) );
  INV_X1 U632 ( .A(G171), .ZN(G301) );
  NAND2_X1 U633 ( .A1(G88), .A2(n794), .ZN(n558) );
  NAND2_X1 U634 ( .A1(G50), .A2(n791), .ZN(n557) );
  NAND2_X1 U635 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U636 ( .A1(G62), .A2(n793), .ZN(n560) );
  NAND2_X1 U637 ( .A1(G75), .A2(n621), .ZN(n559) );
  NAND2_X1 U638 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U639 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U640 ( .A(n563), .B(KEYINPUT80), .ZN(G166) );
  INV_X1 U641 ( .A(G166), .ZN(G303) );
  NAND2_X1 U642 ( .A1(n564), .A2(G87), .ZN(n565) );
  XNOR2_X1 U643 ( .A(KEYINPUT78), .B(n565), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n791), .A2(G49), .ZN(n566) );
  XNOR2_X1 U645 ( .A(n566), .B(KEYINPUT76), .ZN(n568) );
  NAND2_X1 U646 ( .A1(G74), .A2(G651), .ZN(n567) );
  NAND2_X1 U647 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U648 ( .A1(n793), .A2(n569), .ZN(n570) );
  XOR2_X1 U649 ( .A(KEYINPUT77), .B(n570), .Z(n571) );
  NAND2_X1 U650 ( .A1(n572), .A2(n571), .ZN(G288) );
  NAND2_X1 U651 ( .A1(G73), .A2(n621), .ZN(n573) );
  XNOR2_X1 U652 ( .A(n573), .B(KEYINPUT2), .ZN(n580) );
  NAND2_X1 U653 ( .A1(G61), .A2(n793), .ZN(n575) );
  NAND2_X1 U654 ( .A1(G48), .A2(n791), .ZN(n574) );
  NAND2_X1 U655 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U656 ( .A1(G86), .A2(n794), .ZN(n576) );
  XNOR2_X1 U657 ( .A(KEYINPUT79), .B(n576), .ZN(n577) );
  NOR2_X1 U658 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U659 ( .A1(n580), .A2(n579), .ZN(G305) );
  NAND2_X1 U660 ( .A1(G131), .A2(n905), .ZN(n582) );
  NAND2_X1 U661 ( .A1(G95), .A2(n906), .ZN(n581) );
  NAND2_X1 U662 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U663 ( .A(KEYINPUT90), .B(n583), .ZN(n587) );
  NAND2_X1 U664 ( .A1(G107), .A2(n909), .ZN(n585) );
  BUF_X1 U665 ( .A(n600), .Z(n910) );
  NAND2_X1 U666 ( .A1(G119), .A2(n910), .ZN(n584) );
  NAND2_X1 U667 ( .A1(n585), .A2(n584), .ZN(n586) );
  OR2_X1 U668 ( .A1(n587), .A2(n586), .ZN(n888) );
  AND2_X1 U669 ( .A1(n888), .A2(G1991), .ZN(n597) );
  INV_X1 U670 ( .A(G1996), .ZN(n745) );
  NAND2_X1 U671 ( .A1(n905), .A2(G141), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G117), .A2(n909), .ZN(n589) );
  NAND2_X1 U673 ( .A1(G129), .A2(n910), .ZN(n588) );
  NAND2_X1 U674 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U675 ( .A1(n906), .A2(G105), .ZN(n590) );
  XOR2_X1 U676 ( .A(KEYINPUT38), .B(n590), .Z(n591) );
  NOR2_X1 U677 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U679 ( .A(KEYINPUT91), .B(n595), .ZN(n916) );
  NOR2_X1 U680 ( .A1(n745), .A2(n916), .ZN(n596) );
  NOR2_X1 U681 ( .A1(n597), .A2(n596), .ZN(n1010) );
  AND2_X1 U682 ( .A1(G138), .A2(n598), .ZN(n606) );
  NAND2_X1 U683 ( .A1(G102), .A2(n599), .ZN(n604) );
  NAND2_X1 U684 ( .A1(G114), .A2(n909), .ZN(n602) );
  NAND2_X1 U685 ( .A1(G126), .A2(n600), .ZN(n601) );
  AND2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U688 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U689 ( .A(n607), .B(KEYINPUT86), .ZN(n772) );
  NAND2_X1 U690 ( .A1(G160), .A2(G40), .ZN(n612) );
  NOR2_X1 U691 ( .A1(n614), .A2(n612), .ZN(n759) );
  INV_X1 U692 ( .A(n759), .ZN(n608) );
  NOR2_X1 U693 ( .A1(n1010), .A2(n608), .ZN(n749) );
  INV_X1 U694 ( .A(n749), .ZN(n611) );
  XNOR2_X1 U695 ( .A(G1986), .B(G290), .ZN(n935) );
  NAND2_X1 U696 ( .A1(n935), .A2(n759), .ZN(n609) );
  XOR2_X1 U697 ( .A(KEYINPUT87), .B(n609), .Z(n610) );
  NAND2_X1 U698 ( .A1(n611), .A2(n610), .ZN(n731) );
  INV_X1 U699 ( .A(n612), .ZN(n613) );
  XNOR2_X1 U700 ( .A(n617), .B(n616), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n688), .A2(G1341), .ZN(n618) );
  NAND2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n632) );
  NAND2_X1 U703 ( .A1(n793), .A2(G56), .ZN(n620) );
  XOR2_X1 U704 ( .A(KEYINPUT14), .B(n620), .Z(n629) );
  NAND2_X1 U705 ( .A1(n621), .A2(G68), .ZN(n622) );
  XNOR2_X1 U706 ( .A(KEYINPUT67), .B(n622), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n794), .A2(G81), .ZN(n623) );
  XOR2_X1 U708 ( .A(n623), .B(KEYINPUT12), .Z(n624) );
  NOR2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n791), .A2(G43), .ZN(n630) );
  NOR2_X1 U711 ( .A1(n632), .A2(n946), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n634), .B(n633), .ZN(n646) );
  NAND2_X1 U713 ( .A1(G66), .A2(n793), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G79), .A2(n621), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G92), .A2(n794), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G54), .A2(n791), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U719 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U720 ( .A(KEYINPUT15), .B(n641), .Z(n851) );
  INV_X1 U721 ( .A(n851), .ZN(n933) );
  NOR2_X1 U722 ( .A1(n672), .A2(G1348), .ZN(n643) );
  NOR2_X1 U723 ( .A1(G2067), .A2(n688), .ZN(n642) );
  NOR2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n646), .A2(n933), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U728 ( .A(n650), .B(n649), .ZN(n664) );
  NAND2_X1 U729 ( .A1(G2072), .A2(n672), .ZN(n653) );
  NAND2_X1 U730 ( .A1(G1956), .A2(n688), .ZN(n654) );
  XOR2_X1 U731 ( .A(KEYINPUT94), .B(n654), .Z(n655) );
  NOR2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n665) );
  NAND2_X1 U733 ( .A1(G65), .A2(n793), .ZN(n658) );
  NAND2_X1 U734 ( .A1(G53), .A2(n791), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U736 ( .A1(G78), .A2(n621), .ZN(n660) );
  NAND2_X1 U737 ( .A1(G91), .A2(n794), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U739 ( .A1(n662), .A2(n661), .ZN(n936) );
  NAND2_X1 U740 ( .A1(n665), .A2(n936), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n664), .A2(n663), .ZN(n668) );
  NOR2_X1 U742 ( .A1(n665), .A2(n936), .ZN(n666) );
  XOR2_X1 U743 ( .A(n666), .B(KEYINPUT28), .Z(n667) );
  NAND2_X1 U744 ( .A1(n668), .A2(n667), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n670), .B(n669), .ZN(n676) );
  XOR2_X1 U746 ( .A(KEYINPUT25), .B(G2078), .Z(n990) );
  NOR2_X1 U747 ( .A1(n990), .A2(n688), .ZN(n671) );
  XNOR2_X1 U748 ( .A(n671), .B(KEYINPUT92), .ZN(n674) );
  NOR2_X1 U749 ( .A1(n672), .A2(G1961), .ZN(n673) );
  NOR2_X1 U750 ( .A1(n674), .A2(n673), .ZN(n682) );
  OR2_X1 U751 ( .A1(n682), .A2(G301), .ZN(n675) );
  NAND2_X1 U752 ( .A1(n676), .A2(n675), .ZN(n687) );
  NOR2_X1 U753 ( .A1(G2084), .A2(n688), .ZN(n702) );
  NOR2_X1 U754 ( .A1(G1966), .A2(n724), .ZN(n697) );
  NOR2_X1 U755 ( .A1(n702), .A2(n697), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n677), .A2(G8), .ZN(n678) );
  NOR2_X1 U757 ( .A1(G168), .A2(n679), .ZN(n681) );
  XNOR2_X1 U758 ( .A(n681), .B(n680), .ZN(n684) );
  NAND2_X1 U759 ( .A1(n682), .A2(G301), .ZN(n683) );
  NAND2_X1 U760 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U761 ( .A(KEYINPUT31), .B(n685), .ZN(n686) );
  NAND2_X1 U762 ( .A1(n687), .A2(n686), .ZN(n699) );
  NAND2_X1 U763 ( .A1(n699), .A2(G286), .ZN(n694) );
  NOR2_X1 U764 ( .A1(G2090), .A2(n688), .ZN(n689) );
  XNOR2_X1 U765 ( .A(n689), .B(KEYINPUT98), .ZN(n691) );
  NOR2_X1 U766 ( .A1(n724), .A2(G1971), .ZN(n690) );
  NOR2_X1 U767 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U768 ( .A1(G303), .A2(n692), .ZN(n693) );
  NAND2_X1 U769 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U770 ( .A1(n695), .A2(G8), .ZN(n696) );
  XNOR2_X1 U771 ( .A(n696), .B(KEYINPUT32), .ZN(n706) );
  INV_X1 U772 ( .A(n697), .ZN(n698) );
  XNOR2_X1 U773 ( .A(n701), .B(n700), .ZN(n704) );
  NAND2_X1 U774 ( .A1(G8), .A2(n702), .ZN(n703) );
  NAND2_X1 U775 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U777 ( .A(n708), .B(n707), .ZN(n718) );
  NOR2_X1 U778 ( .A1(G1976), .A2(G288), .ZN(n713) );
  NOR2_X1 U779 ( .A1(G303), .A2(G1971), .ZN(n709) );
  NOR2_X1 U780 ( .A1(n713), .A2(n709), .ZN(n940) );
  NAND2_X1 U781 ( .A1(n718), .A2(n940), .ZN(n710) );
  NAND2_X1 U782 ( .A1(G1976), .A2(G288), .ZN(n939) );
  NAND2_X1 U783 ( .A1(n710), .A2(n939), .ZN(n711) );
  NOR2_X1 U784 ( .A1(n724), .A2(n711), .ZN(n712) );
  NOR2_X1 U785 ( .A1(KEYINPUT33), .A2(n712), .ZN(n716) );
  NAND2_X1 U786 ( .A1(n713), .A2(KEYINPUT33), .ZN(n714) );
  NOR2_X1 U787 ( .A1(n714), .A2(n724), .ZN(n715) );
  NOR2_X1 U788 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U789 ( .A(G1981), .B(G305), .Z(n931) );
  NAND2_X1 U790 ( .A1(n717), .A2(n931), .ZN(n727) );
  NOR2_X1 U791 ( .A1(G2090), .A2(G303), .ZN(n719) );
  NAND2_X1 U792 ( .A1(G8), .A2(n719), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n718), .A2(n720), .ZN(n721) );
  NAND2_X1 U794 ( .A1(n721), .A2(n724), .ZN(n725) );
  NOR2_X1 U795 ( .A1(G1981), .A2(G305), .ZN(n722) );
  XOR2_X1 U796 ( .A(n722), .B(KEYINPUT24), .Z(n723) );
  NAND2_X1 U797 ( .A1(n727), .A2(n726), .ZN(n729) );
  NOR2_X1 U798 ( .A1(n731), .A2(n730), .ZN(n744) );
  XNOR2_X1 U799 ( .A(G2067), .B(KEYINPUT37), .ZN(n757) );
  XNOR2_X1 U800 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n742) );
  NAND2_X1 U801 ( .A1(G116), .A2(n909), .ZN(n733) );
  NAND2_X1 U802 ( .A1(G128), .A2(n910), .ZN(n732) );
  NAND2_X1 U803 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U804 ( .A(KEYINPUT35), .B(n734), .ZN(n740) );
  NAND2_X1 U805 ( .A1(n906), .A2(G104), .ZN(n735) );
  XNOR2_X1 U806 ( .A(n735), .B(KEYINPUT88), .ZN(n737) );
  NAND2_X1 U807 ( .A1(G140), .A2(n905), .ZN(n736) );
  NAND2_X1 U808 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U809 ( .A(KEYINPUT34), .B(n738), .Z(n739) );
  NAND2_X1 U810 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U811 ( .A(n742), .B(n741), .ZN(n919) );
  NOR2_X1 U812 ( .A1(n757), .A2(n919), .ZN(n754) );
  NAND2_X1 U813 ( .A1(n754), .A2(n759), .ZN(n743) );
  NAND2_X1 U814 ( .A1(n744), .A2(n743), .ZN(n762) );
  XOR2_X1 U815 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n753) );
  AND2_X1 U816 ( .A1(n745), .A2(n916), .ZN(n1007) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n747) );
  NOR2_X1 U818 ( .A1(G1991), .A2(n888), .ZN(n746) );
  XOR2_X1 U819 ( .A(KEYINPUT101), .B(n746), .Z(n1015) );
  NOR2_X1 U820 ( .A1(n747), .A2(n1015), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U822 ( .A(n750), .B(KEYINPUT102), .ZN(n751) );
  NOR2_X1 U823 ( .A1(n1007), .A2(n751), .ZN(n752) );
  XNOR2_X1 U824 ( .A(n753), .B(n752), .ZN(n755) );
  INV_X1 U825 ( .A(n754), .ZN(n1017) );
  NAND2_X1 U826 ( .A1(n755), .A2(n1017), .ZN(n756) );
  XNOR2_X1 U827 ( .A(n756), .B(KEYINPUT104), .ZN(n758) );
  NAND2_X1 U828 ( .A1(n757), .A2(n919), .ZN(n1019) );
  NAND2_X1 U829 ( .A1(n758), .A2(n1019), .ZN(n760) );
  NAND2_X1 U830 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U831 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U832 ( .A(n763), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U834 ( .A1(G111), .A2(n909), .ZN(n765) );
  NAND2_X1 U835 ( .A1(G135), .A2(n905), .ZN(n764) );
  NAND2_X1 U836 ( .A1(n765), .A2(n764), .ZN(n768) );
  NAND2_X1 U837 ( .A1(n910), .A2(G123), .ZN(n766) );
  XOR2_X1 U838 ( .A(KEYINPUT18), .B(n766), .Z(n767) );
  NOR2_X1 U839 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U840 ( .A1(n906), .A2(G99), .ZN(n769) );
  NAND2_X1 U841 ( .A1(n770), .A2(n769), .ZN(n1012) );
  XNOR2_X1 U842 ( .A(G2096), .B(n1012), .ZN(n771) );
  OR2_X1 U843 ( .A1(G2100), .A2(n771), .ZN(G156) );
  INV_X1 U844 ( .A(n936), .ZN(G299) );
  INV_X1 U845 ( .A(G57), .ZN(G237) );
  NAND2_X1 U846 ( .A1(G7), .A2(G661), .ZN(n774) );
  XNOR2_X1 U847 ( .A(n774), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U848 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n776) );
  INV_X1 U849 ( .A(G223), .ZN(n833) );
  NAND2_X1 U850 ( .A1(G567), .A2(n833), .ZN(n775) );
  XNOR2_X1 U851 ( .A(n776), .B(n775), .ZN(G234) );
  INV_X1 U852 ( .A(G860), .ZN(n783) );
  OR2_X1 U853 ( .A1(n946), .A2(n783), .ZN(G153) );
  NOR2_X1 U854 ( .A1(n851), .A2(G868), .ZN(n777) );
  XNOR2_X1 U855 ( .A(n777), .B(KEYINPUT69), .ZN(n779) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n778) );
  NAND2_X1 U857 ( .A1(n779), .A2(n778), .ZN(G284) );
  INV_X1 U858 ( .A(G868), .ZN(n815) );
  XNOR2_X1 U859 ( .A(KEYINPUT70), .B(n815), .ZN(n780) );
  NOR2_X1 U860 ( .A1(G286), .A2(n780), .ZN(n782) );
  NOR2_X1 U861 ( .A1(G868), .A2(G299), .ZN(n781) );
  NOR2_X1 U862 ( .A1(n782), .A2(n781), .ZN(G297) );
  NAND2_X1 U863 ( .A1(n783), .A2(G559), .ZN(n784) );
  NAND2_X1 U864 ( .A1(n784), .A2(n851), .ZN(n785) );
  XNOR2_X1 U865 ( .A(n785), .B(KEYINPUT16), .ZN(n786) );
  XOR2_X1 U866 ( .A(KEYINPUT71), .B(n786), .Z(G148) );
  NAND2_X1 U867 ( .A1(n851), .A2(G868), .ZN(n787) );
  NOR2_X1 U868 ( .A1(G559), .A2(n787), .ZN(n788) );
  XNOR2_X1 U869 ( .A(n788), .B(KEYINPUT72), .ZN(n790) );
  NOR2_X1 U870 ( .A1(n946), .A2(G868), .ZN(n789) );
  NOR2_X1 U871 ( .A1(n790), .A2(n789), .ZN(G282) );
  NAND2_X1 U872 ( .A1(G55), .A2(n791), .ZN(n792) );
  XNOR2_X1 U873 ( .A(n792), .B(KEYINPUT74), .ZN(n801) );
  NAND2_X1 U874 ( .A1(G67), .A2(n793), .ZN(n796) );
  NAND2_X1 U875 ( .A1(G93), .A2(n794), .ZN(n795) );
  NAND2_X1 U876 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U877 ( .A1(G80), .A2(n621), .ZN(n797) );
  XNOR2_X1 U878 ( .A(KEYINPUT73), .B(n797), .ZN(n798) );
  NOR2_X1 U879 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U880 ( .A1(n801), .A2(n800), .ZN(n814) );
  NAND2_X1 U881 ( .A1(G559), .A2(n851), .ZN(n802) );
  XNOR2_X1 U882 ( .A(n802), .B(n946), .ZN(n811) );
  NOR2_X1 U883 ( .A1(n811), .A2(G860), .ZN(n803) );
  XNOR2_X1 U884 ( .A(n803), .B(KEYINPUT75), .ZN(n804) );
  XNOR2_X1 U885 ( .A(n814), .B(n804), .ZN(G145) );
  XNOR2_X1 U886 ( .A(G303), .B(G288), .ZN(n805) );
  XNOR2_X1 U887 ( .A(n805), .B(n814), .ZN(n806) );
  XNOR2_X1 U888 ( .A(KEYINPUT81), .B(n806), .ZN(n808) );
  XNOR2_X1 U889 ( .A(G290), .B(KEYINPUT19), .ZN(n807) );
  XNOR2_X1 U890 ( .A(n808), .B(n807), .ZN(n809) );
  XNOR2_X1 U891 ( .A(n809), .B(G299), .ZN(n810) );
  XNOR2_X1 U892 ( .A(n810), .B(G305), .ZN(n854) );
  XNOR2_X1 U893 ( .A(n854), .B(n811), .ZN(n812) );
  NAND2_X1 U894 ( .A1(n812), .A2(G868), .ZN(n813) );
  XNOR2_X1 U895 ( .A(n813), .B(KEYINPUT82), .ZN(n817) );
  NAND2_X1 U896 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U897 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U898 ( .A1(G2084), .A2(G2078), .ZN(n820) );
  XNOR2_X1 U899 ( .A(KEYINPUT83), .B(KEYINPUT20), .ZN(n818) );
  XNOR2_X1 U900 ( .A(n818), .B(KEYINPUT84), .ZN(n819) );
  XNOR2_X1 U901 ( .A(n820), .B(n819), .ZN(n821) );
  NAND2_X1 U902 ( .A1(n821), .A2(G2090), .ZN(n822) );
  XNOR2_X1 U903 ( .A(KEYINPUT21), .B(n822), .ZN(n823) );
  NAND2_X1 U904 ( .A1(n823), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U905 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U906 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n825) );
  NAND2_X1 U907 ( .A1(G132), .A2(G82), .ZN(n824) );
  XNOR2_X1 U908 ( .A(n825), .B(n824), .ZN(n826) );
  NOR2_X1 U909 ( .A1(n826), .A2(G218), .ZN(n827) );
  NAND2_X1 U910 ( .A1(G96), .A2(n827), .ZN(n839) );
  NAND2_X1 U911 ( .A1(n839), .A2(G2106), .ZN(n831) );
  NAND2_X1 U912 ( .A1(G69), .A2(G120), .ZN(n828) );
  NOR2_X1 U913 ( .A1(G237), .A2(n828), .ZN(n829) );
  NAND2_X1 U914 ( .A1(G108), .A2(n829), .ZN(n840) );
  NAND2_X1 U915 ( .A1(n840), .A2(G567), .ZN(n830) );
  NAND2_X1 U916 ( .A1(n831), .A2(n830), .ZN(n928) );
  NAND2_X1 U917 ( .A1(G661), .A2(G483), .ZN(n832) );
  NOR2_X1 U918 ( .A1(n928), .A2(n832), .ZN(n838) );
  NAND2_X1 U919 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n833), .ZN(G217) );
  INV_X1 U921 ( .A(G661), .ZN(n835) );
  NAND2_X1 U922 ( .A1(G2), .A2(G15), .ZN(n834) );
  NOR2_X1 U923 ( .A1(n835), .A2(n834), .ZN(n836) );
  XOR2_X1 U924 ( .A(KEYINPUT106), .B(n836), .Z(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U926 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U928 ( .A(G132), .ZN(G219) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G82), .ZN(G220) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U935 ( .A(G1348), .B(G2454), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n841), .B(G2430), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n842), .B(G1341), .ZN(n848) );
  XOR2_X1 U938 ( .A(G2443), .B(G2427), .Z(n844) );
  XNOR2_X1 U939 ( .A(G2438), .B(G2446), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(n846) );
  XOR2_X1 U941 ( .A(G2451), .B(G2435), .Z(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n848), .B(n847), .ZN(n849) );
  NAND2_X1 U944 ( .A1(n849), .A2(G14), .ZN(n850) );
  XNOR2_X1 U945 ( .A(KEYINPUT105), .B(n850), .ZN(G401) );
  XOR2_X1 U946 ( .A(KEYINPUT115), .B(G286), .Z(n853) );
  XNOR2_X1 U947 ( .A(G171), .B(n851), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n853), .B(n852), .ZN(n856) );
  XOR2_X1 U949 ( .A(n946), .B(n854), .Z(n855) );
  XNOR2_X1 U950 ( .A(n856), .B(n855), .ZN(n857) );
  NOR2_X1 U951 ( .A1(G37), .A2(n857), .ZN(G397) );
  XNOR2_X1 U952 ( .A(G1996), .B(KEYINPUT110), .ZN(n867) );
  XOR2_X1 U953 ( .A(G1981), .B(G1956), .Z(n859) );
  XNOR2_X1 U954 ( .A(G1991), .B(G1966), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U956 ( .A(G1976), .B(G1971), .Z(n861) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1961), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U959 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U960 ( .A(G2474), .B(KEYINPUT41), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U962 ( .A(n867), .B(n866), .ZN(G229) );
  XNOR2_X1 U963 ( .A(G2090), .B(G2084), .ZN(n868) );
  XNOR2_X1 U964 ( .A(n868), .B(KEYINPUT108), .ZN(n878) );
  XOR2_X1 U965 ( .A(KEYINPUT109), .B(G2678), .Z(n870) );
  XNOR2_X1 U966 ( .A(KEYINPUT42), .B(G2096), .ZN(n869) );
  XNOR2_X1 U967 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U968 ( .A(G2100), .B(G2072), .Z(n872) );
  XNOR2_X1 U969 ( .A(G2067), .B(G2078), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U971 ( .A(n874), .B(n873), .Z(n876) );
  XNOR2_X1 U972 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n875) );
  XNOR2_X1 U973 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U974 ( .A(n878), .B(n877), .ZN(G227) );
  NAND2_X1 U975 ( .A1(G124), .A2(n910), .ZN(n879) );
  XNOR2_X1 U976 ( .A(n879), .B(KEYINPUT44), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n909), .A2(G112), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n885) );
  NAND2_X1 U979 ( .A1(G136), .A2(n905), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G100), .A2(n906), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n884) );
  NOR2_X1 U982 ( .A1(n885), .A2(n884), .ZN(G162) );
  XOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n886) );
  XNOR2_X1 U984 ( .A(n1012), .B(n886), .ZN(n887) );
  XOR2_X1 U985 ( .A(n887), .B(KEYINPUT113), .Z(n890) );
  XOR2_X1 U986 ( .A(n888), .B(KEYINPUT46), .Z(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n901) );
  NAND2_X1 U988 ( .A1(G118), .A2(n909), .ZN(n892) );
  NAND2_X1 U989 ( .A1(G130), .A2(n910), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n899) );
  XNOR2_X1 U991 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n897) );
  NAND2_X1 U992 ( .A1(n906), .A2(G106), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n905), .A2(G142), .ZN(n893) );
  XOR2_X1 U994 ( .A(KEYINPUT111), .B(n893), .Z(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U996 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U999 ( .A(G164), .B(G160), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1001 ( .A(n904), .B(G162), .Z(n918) );
  NAND2_X1 U1002 ( .A1(G139), .A2(n905), .ZN(n908) );
  NAND2_X1 U1003 ( .A1(G103), .A2(n906), .ZN(n907) );
  NAND2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n915) );
  NAND2_X1 U1005 ( .A1(G115), .A2(n909), .ZN(n912) );
  NAND2_X1 U1006 ( .A1(G127), .A2(n910), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1008 ( .A(KEYINPUT47), .B(n913), .Z(n914) );
  NOR2_X1 U1009 ( .A1(n915), .A2(n914), .ZN(n1002) );
  XNOR2_X1 U1010 ( .A(n916), .B(n1002), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(n918), .B(n917), .ZN(n920) );
  XOR2_X1 U1012 ( .A(n920), .B(n919), .Z(n921) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n921), .ZN(G395) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n928), .ZN(n925) );
  NOR2_X1 U1015 ( .A1(G229), .A2(G227), .ZN(n922) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1017 ( .A1(G397), .A2(n923), .ZN(n924) );
  NAND2_X1 U1018 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1019 ( .A1(n926), .A2(G395), .ZN(n927) );
  XNOR2_X1 U1020 ( .A(n927), .B(KEYINPUT116), .ZN(G308) );
  INV_X1 U1021 ( .A(G308), .ZN(G225) );
  INV_X1 U1022 ( .A(n928), .ZN(G319) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1024 ( .A(KEYINPUT56), .B(G16), .ZN(n956) );
  XOR2_X1 U1025 ( .A(G1966), .B(G168), .Z(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT123), .B(n929), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(KEYINPUT57), .B(n932), .ZN(n954) );
  XNOR2_X1 U1029 ( .A(G171), .B(G1961), .ZN(n951) );
  XNOR2_X1 U1030 ( .A(G1348), .B(n933), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n945) );
  XNOR2_X1 U1032 ( .A(G1956), .B(n936), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(G1971), .A2(G303), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(n943), .B(KEYINPUT124), .ZN(n944) );
  NAND2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n949) );
  XOR2_X1 U1039 ( .A(G1341), .B(n946), .Z(n947) );
  XNOR2_X1 U1040 ( .A(KEYINPUT125), .B(n947), .ZN(n948) );
  NOR2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1042 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1043 ( .A(KEYINPUT126), .B(n952), .Z(n953) );
  NAND2_X1 U1044 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1045 ( .A1(n956), .A2(n955), .ZN(n1032) );
  XNOR2_X1 U1046 ( .A(G1966), .B(G21), .ZN(n958) );
  XNOR2_X1 U1047 ( .A(G1961), .B(G5), .ZN(n957) );
  NOR2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n968) );
  XOR2_X1 U1049 ( .A(G1348), .B(KEYINPUT59), .Z(n959) );
  XNOR2_X1 U1050 ( .A(G4), .B(n959), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G20), .B(G1956), .ZN(n960) );
  NOR2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n965) );
  XNOR2_X1 U1053 ( .A(G1341), .B(G19), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G6), .B(G1981), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1057 ( .A(KEYINPUT60), .B(n966), .Z(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n975) );
  XNOR2_X1 U1059 ( .A(G1986), .B(G24), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(G1971), .B(G22), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n972) );
  XOR2_X1 U1062 ( .A(G1976), .B(G23), .Z(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(KEYINPUT58), .B(n973), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(n976), .B(KEYINPUT61), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(G16), .B(KEYINPUT127), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(G11), .A2(n979), .ZN(n1030) );
  XNOR2_X1 U1070 ( .A(G2084), .B(G34), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(n980), .B(KEYINPUT54), .ZN(n998) );
  XOR2_X1 U1072 ( .A(G2090), .B(G35), .Z(n981) );
  XNOR2_X1 U1073 ( .A(KEYINPUT119), .B(n981), .ZN(n995) );
  XNOR2_X1 U1074 ( .A(G1996), .B(G32), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(G33), .B(G2072), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n989) );
  XOR2_X1 U1077 ( .A(G25), .B(G1991), .Z(n984) );
  NAND2_X1 U1078 ( .A1(n984), .A2(G28), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(KEYINPUT120), .B(G2067), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(G26), .B(n985), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(G27), .B(n990), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(n993), .B(KEYINPUT53), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n996), .B(KEYINPUT121), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(KEYINPUT122), .B(n999), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(G29), .A2(n1000), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(n1001), .B(KEYINPUT55), .ZN(n1028) );
  XOR2_X1 U1092 ( .A(G2072), .B(n1002), .Z(n1004) );
  XOR2_X1 U1093 ( .A(G164), .B(G2078), .Z(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT50), .B(n1005), .ZN(n1024) );
  XOR2_X1 U1096 ( .A(G2090), .B(G162), .Z(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1098 ( .A(KEYINPUT51), .B(n1008), .Z(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT118), .B(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1022) );
  XNOR2_X1 U1101 ( .A(G160), .B(G2084), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(n1018), .B(KEYINPUT117), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(KEYINPUT52), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(G29), .A2(n1026), .ZN(n1027) );
  NAND2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1112 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1113 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

