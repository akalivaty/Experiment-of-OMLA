//key=1010101010101010101010101010101010101010101010101010101010101010


module locked_locked_c3540 ( G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, 
        G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, 
        G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, 
        G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, 
        G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, 
        G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, 
        G409, G405, G402, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, 
        KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, 
        KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, 
        KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, 
        KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, 
        KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, 
        KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, 
        KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, 
        KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, 
        KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, 
        KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, 
        KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, 
        KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, 
        KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, 
        KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, 
        KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, 
        KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, 
        KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92, 
        KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, 
        KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80, 
        KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, 
        KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, 
        KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
         G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
         G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
         G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330,
         G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60,
         KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55,
         KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50,
         KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45,
         KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40,
         KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35,
         KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30,
         KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25,
         KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20,
         KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15,
         KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9,
         KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3,
         KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126,
         KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121,
         KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116,
         KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111,
         KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106,
         KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101,
         KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96,
         KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91,
         KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86,
         KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81,
         KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76,
         KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71,
         KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66,
         KEYINPUT65, KEYINPUT64;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
         G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire   n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046;

  XOR2_X1 U1018 ( .A(KEYINPUT29), .B(n1679), .Z(n1752) );
  INV_X1 U1019 ( .A(n1587), .ZN(n1307) );
  INV_X1 U1020 ( .A(G20), .ZN(n1155) );
  NOR2_X2 U1021 ( .A1(n1730), .A2(n1729), .ZN(n1748) );
  INV_X2 U1022 ( .A(n1138), .ZN(n1121) );
  XNOR2_X2 U1023 ( .A(n1115), .B(KEYINPUT2), .ZN(n1138) );
  AND2_X1 U1024 ( .A1(n1311), .A2(n1310), .ZN(n1111) );
  INV_X1 U1025 ( .A(n1886), .ZN(n1881) );
  INV_X1 U1026 ( .A(n1313), .ZN(n1614) );
  INV_X1 U1027 ( .A(n1424), .ZN(n1623) );
  AND2_X1 U1028 ( .A1(n1143), .A2(n1148), .ZN(n1332) );
  INV_X1 U1029 ( .A(G33), .ZN(n1246) );
  NAND2_X1 U1030 ( .A1(n1727), .A2(n1011), .ZN(G381) );
  NOR2_X1 U1031 ( .A1(n1819), .A2(n1746), .ZN(n1747) );
  XNOR2_X1 U1032 ( .A(n1745), .B(n1744), .ZN(n1819) );
  AND2_X1 U1033 ( .A1(n1877), .A2(n1876), .ZN(n1043) );
  NOR2_X1 U1034 ( .A1(n1327), .A2(n1320), .ZN(n1321) );
  XNOR2_X1 U1035 ( .A(n1095), .B(KEYINPUT0), .ZN(n1327) );
  NAND2_X1 U1036 ( .A1(n1096), .A2(n1074), .ZN(n1095) );
  NOR2_X1 U1037 ( .A1(n1332), .A2(n1034), .ZN(n1033) );
  BUF_X1 U1038 ( .A(n1304), .Z(n1633) );
  XNOR2_X1 U1039 ( .A(n1140), .B(n1139), .ZN(n1304) );
  NOR2_X2 U1040 ( .A1(n1075), .A2(n1120), .ZN(n1611) );
  OR2_X1 U1041 ( .A1(n1415), .A2(n1123), .ZN(n1117) );
  NOR2_X2 U1042 ( .A1(n1199), .A2(G1), .ZN(n1363) );
  OR2_X1 U1043 ( .A1(n2017), .A2(n1134), .ZN(n1136) );
  NAND2_X1 U1044 ( .A1(G13), .A2(G1), .ZN(n1115) );
  AND2_X1 U1045 ( .A1(n1101), .A2(n1003), .ZN(n1100) );
  NAND2_X1 U1046 ( .A1(n1317), .A2(n1111), .ZN(n1378) );
  XNOR2_X1 U1047 ( .A(n1065), .B(KEYINPUT71), .ZN(n1123) );
  AND2_X1 U1048 ( .A1(n1023), .A2(n1303), .ZN(n1325) );
  NOR2_X1 U1049 ( .A1(n1306), .A2(n1001), .ZN(n1023) );
  NOR2_X1 U1050 ( .A1(n1045), .A2(n1880), .ZN(n1044) );
  AND2_X1 U1051 ( .A1(n1380), .A2(n1126), .ZN(n1127) );
  XNOR2_X1 U1052 ( .A(n1685), .B(n1053), .ZN(n1817) );
  INV_X1 U1053 ( .A(KEYINPUT38), .ZN(n1053) );
  OR2_X1 U1054 ( .A1(n1323), .A2(n1547), .ZN(n1040) );
  XNOR2_X1 U1055 ( .A(n1026), .B(n1025), .ZN(n1966) );
  XNOR2_X1 U1056 ( .A(n1960), .B(n1027), .ZN(n1026) );
  XNOR2_X1 U1057 ( .A(G381), .B(G387), .ZN(n1025) );
  XNOR2_X1 U1058 ( .A(n1958), .B(n1028), .ZN(n1027) );
  XNOR2_X1 U1059 ( .A(n1071), .B(n1389), .ZN(n1070) );
  NAND2_X1 U1060 ( .A1(n1073), .A2(n1072), .ZN(n1071) );
  INV_X1 U1061 ( .A(n1322), .ZN(n1072) );
  NAND2_X1 U1062 ( .A1(n1611), .A2(G257), .ZN(n1009) );
  NOR2_X1 U1063 ( .A1(n1377), .A2(n1375), .ZN(n1031) );
  AND2_X1 U1064 ( .A1(n1765), .A2(G33), .ZN(n1103) );
  NAND2_X1 U1065 ( .A1(n1121), .A2(n1087), .ZN(n1313) );
  AND2_X1 U1066 ( .A1(n1246), .A2(n1120), .ZN(n1087) );
  NAND2_X1 U1067 ( .A1(n1121), .A2(n1246), .ZN(n1075) );
  NOR2_X1 U1068 ( .A1(n1075), .A2(G20), .ZN(n1622) );
  NAND2_X1 U1069 ( .A1(n1032), .A2(n1881), .ZN(n1392) );
  XNOR2_X1 U1070 ( .A(n1386), .B(KEYINPUT85), .ZN(n1032) );
  NAND2_X1 U1071 ( .A1(n2005), .A2(n1886), .ZN(n1082) );
  NAND2_X1 U1072 ( .A1(n1109), .A2(n1105), .ZN(n1606) );
  NAND2_X1 U1073 ( .A1(n1022), .A2(n1018), .ZN(n1096) );
  NOR2_X1 U1074 ( .A1(n1325), .A2(n999), .ZN(n1022) );
  XNOR2_X1 U1075 ( .A(n1020), .B(n1019), .ZN(n1018) );
  INV_X1 U1076 ( .A(KEYINPUT70), .ZN(n1116) );
  NOR2_X1 U1077 ( .A1(n1054), .A2(n1055), .ZN(n1037) );
  INV_X1 U1078 ( .A(KEYINPUT77), .ZN(n1056) );
  NOR2_X1 U1079 ( .A1(n1671), .A2(n1670), .ZN(n1732) );
  NOR2_X1 U1080 ( .A1(n1881), .A2(n1728), .ZN(n1729) );
  NOR2_X1 U1081 ( .A1(n1752), .A2(n1881), .ZN(n1088) );
  INV_X1 U1082 ( .A(G330), .ZN(n1061) );
  OR2_X1 U1083 ( .A1(n1368), .A2(n1086), .ZN(n1085) );
  NAND2_X1 U1084 ( .A1(n1353), .A2(n1352), .ZN(n1372) );
  NAND2_X1 U1085 ( .A1(n1439), .A2(n1437), .ZN(n1667) );
  NAND2_X1 U1086 ( .A1(n1281), .A2(n1283), .ZN(n1341) );
  AND2_X1 U1087 ( .A1(n1372), .A2(n1085), .ZN(n1387) );
  XNOR2_X1 U1088 ( .A(n1338), .B(KEYINPUT52), .ZN(n1875) );
  XNOR2_X1 U1089 ( .A(n1013), .B(n1817), .ZN(n1012) );
  XNOR2_X1 U1090 ( .A(n1746), .B(KEYINPUT46), .ZN(n1013) );
  INV_X1 U1091 ( .A(KEYINPUT41), .ZN(n1076) );
  XNOR2_X1 U1092 ( .A(n1052), .B(n1819), .ZN(n1051) );
  XOR2_X1 U1093 ( .A(KEYINPUT1), .B(n1113), .Z(n1820) );
  NOR2_X1 U1094 ( .A1(n1151), .A2(n1150), .ZN(n1152) );
  NOR2_X1 U1095 ( .A1(G41), .A2(n1979), .ZN(n2014) );
  XNOR2_X1 U1096 ( .A(n1963), .B(KEYINPUT63), .ZN(n1964) );
  AND2_X1 U1097 ( .A1(n1308), .A2(G294), .ZN(n1048) );
  NAND2_X1 U1098 ( .A1(n1047), .A2(KEYINPUT14), .ZN(n1049) );
  NAND2_X1 U1099 ( .A1(n1307), .A2(G294), .ZN(n1047) );
  AND2_X1 U1100 ( .A1(n1103), .A2(KEYINPUT65), .ZN(n1102) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1316), .ZN(n1317) );
  NAND2_X1 U1102 ( .A1(n1009), .A2(n1315), .ZN(n1010) );
  OR2_X1 U1103 ( .A1(n1623), .A2(n1420), .ZN(n1297) );
  NAND2_X1 U1104 ( .A1(n1030), .A2(n1029), .ZN(n1385) );
  NOR2_X1 U1105 ( .A1(n1376), .A2(n1144), .ZN(n1029) );
  XNOR2_X1 U1106 ( .A(n1031), .B(KEYINPUT18), .ZN(n1030) );
  OR2_X1 U1107 ( .A1(n1129), .A2(G20), .ZN(n1017) );
  NOR2_X1 U1108 ( .A1(n1584), .A2(n1583), .ZN(n1586) );
  XNOR2_X1 U1109 ( .A(n1015), .B(n1014), .ZN(n1301) );
  INV_X1 U1110 ( .A(KEYINPUT16), .ZN(n1014) );
  NOR2_X1 U1111 ( .A1(n1017), .A2(n1016), .ZN(n1015) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1317), .ZN(n1020) );
  AND2_X1 U1113 ( .A1(n1111), .A2(n1126), .ZN(n1021) );
  INV_X1 U1114 ( .A(KEYINPUT15), .ZN(n1019) );
  XNOR2_X1 U1115 ( .A(n1118), .B(n1119), .ZN(n1054) );
  OR2_X1 U1116 ( .A1(n1108), .A2(n1125), .ZN(n1055) );
  INV_X1 U1117 ( .A(KEYINPUT4), .ZN(n1139) );
  INV_X1 U1118 ( .A(n1666), .ZN(n1045) );
  XNOR2_X1 U1119 ( .A(n1360), .B(n1359), .ZN(n1361) );
  XNOR2_X1 U1120 ( .A(n1358), .B(KEYINPUT8), .ZN(n1359) );
  INV_X1 U1121 ( .A(KEYINPUT69), .ZN(n1358) );
  NOR2_X1 U1122 ( .A1(n1346), .A2(n1345), .ZN(n1347) );
  INV_X1 U1123 ( .A(n1017), .ZN(n1626) );
  NAND2_X1 U1124 ( .A1(n1082), .A2(n1392), .ZN(n1756) );
  NOR2_X1 U1125 ( .A1(n1678), .A2(n1677), .ZN(n1679) );
  NOR2_X1 U1126 ( .A1(n2006), .A2(n1756), .ZN(n2020) );
  AND2_X1 U1127 ( .A1(n1392), .A2(G330), .ZN(n1081) );
  INV_X1 U1128 ( .A(n1096), .ZN(n1324) );
  AND2_X1 U1129 ( .A1(n1609), .A2(n1106), .ZN(n1659) );
  NOR2_X1 U1130 ( .A1(n1621), .A2(n1620), .ZN(n1640) );
  AND2_X1 U1131 ( .A1(n1318), .A2(n1319), .ZN(n1094) );
  NOR2_X1 U1132 ( .A1(n1261), .A2(n1260), .ZN(n1262) );
  INV_X1 U1133 ( .A(G393), .ZN(n1028) );
  XNOR2_X1 U1134 ( .A(G396), .B(n1957), .ZN(n1958) );
  INV_X1 U1135 ( .A(G45), .ZN(n1199) );
  NAND2_X1 U1136 ( .A1(n1059), .A2(n1057), .ZN(n1551) );
  AND2_X1 U1137 ( .A1(n1062), .A2(n1060), .ZN(n1059) );
  NAND2_X1 U1138 ( .A1(G343), .A2(n1761), .ZN(n1886) );
  AND2_X1 U1139 ( .A1(n1342), .A2(n1097), .ZN(n1373) );
  NOR2_X1 U1140 ( .A1(n1387), .A2(n1098), .ZN(n1097) );
  NOR2_X1 U1141 ( .A1(n1372), .A2(n1371), .ZN(n1880) );
  XNOR2_X1 U1142 ( .A(n1033), .B(KEYINPUT11), .ZN(n1388) );
  AND2_X1 U1143 ( .A1(n1035), .A2(n1145), .ZN(n1034) );
  NAND2_X1 U1144 ( .A1(n1084), .A2(n1083), .ZN(n1951) );
  INV_X1 U1145 ( .A(n1387), .ZN(n1084) );
  INV_X1 U1146 ( .A(n1880), .ZN(n1083) );
  NOR2_X1 U1147 ( .A1(n1004), .A2(n1214), .ZN(n1038) );
  XNOR2_X1 U1148 ( .A(n1040), .B(KEYINPUT62), .ZN(n1039) );
  AND2_X1 U1149 ( .A1(n1024), .A2(G330), .ZN(n1064) );
  NOR2_X1 U1150 ( .A1(n1739), .A2(n1656), .ZN(n1681) );
  NAND2_X1 U1151 ( .A1(n1012), .A2(n2014), .ZN(n1011) );
  XNOR2_X1 U1152 ( .A(n1093), .B(n1771), .ZN(n1091) );
  NAND2_X1 U1153 ( .A1(n1871), .A2(n1870), .ZN(G378) );
  NOR2_X1 U1154 ( .A1(n1869), .A2(n1110), .ZN(n1870) );
  NAND2_X1 U1155 ( .A1(n1051), .A2(n2014), .ZN(n1871) );
  INV_X1 U1156 ( .A(KEYINPUT55), .ZN(n1068) );
  NAND2_X1 U1157 ( .A1(n1041), .A2(n1000), .ZN(n1069) );
  AND2_X1 U1158 ( .A1(n1378), .A2(n1605), .ZN(n999) );
  INV_X1 U1159 ( .A(G1), .ZN(n2017) );
  OR2_X1 U1160 ( .A1(n1956), .A2(n1955), .ZN(n1000) );
  AND2_X1 U1161 ( .A1(G87), .A2(n1622), .ZN(n1001) );
  XNOR2_X1 U1162 ( .A(n1069), .B(n1068), .ZN(G387) );
  XNOR2_X1 U1163 ( .A(n1152), .B(KEYINPUT79), .ZN(n1323) );
  AND2_X1 U1164 ( .A1(G190), .A2(n1380), .ZN(n1002) );
  OR2_X1 U1165 ( .A1(n1103), .A2(KEYINPUT65), .ZN(n1003) );
  AND2_X1 U1166 ( .A1(n1183), .A2(n1182), .ZN(n1004) );
  AND2_X1 U1167 ( .A1(n1039), .A2(n1038), .ZN(n1005) );
  OR2_X1 U1168 ( .A1(n1138), .A2(n1067), .ZN(n1066) );
  OR2_X1 U1169 ( .A1(n1121), .A2(KEYINPUT65), .ZN(n1006) );
  AND2_X1 U1170 ( .A1(n1037), .A2(n1036), .ZN(n1380) );
  AND2_X1 U1171 ( .A1(n1815), .A2(n1820), .ZN(n1007) );
  NAND2_X1 U1172 ( .A1(n1282), .A2(n1341), .ZN(n1389) );
  AND2_X1 U1173 ( .A1(n1077), .A2(n1007), .ZN(n1008) );
  INV_X1 U1174 ( .A(G116), .ZN(n1016) );
  OR2_X1 U1175 ( .A1(n1339), .A2(n1881), .ZN(n1073) );
  NOR2_X2 U1176 ( .A1(n1126), .A2(n1177), .ZN(n1934) );
  NOR2_X2 U1177 ( .A1(n1126), .A2(n1171), .ZN(n1931) );
  NOR2_X2 U1178 ( .A1(n1126), .A2(n1156), .ZN(n1927) );
  NOR2_X2 U1179 ( .A1(G179), .A2(n1171), .ZN(n1933) );
  XNOR2_X2 U1180 ( .A(n1168), .B(KEYINPUT87), .ZN(n1926) );
  INV_X1 U1181 ( .A(n1328), .ZN(n1329) );
  NOR2_X1 U1182 ( .A1(n1328), .A2(n1389), .ZN(n1390) );
  XNOR2_X1 U1183 ( .A(n1328), .B(n1336), .ZN(n1337) );
  NOR2_X1 U1184 ( .A1(n1024), .A2(n1547), .ZN(n1548) );
  NAND2_X1 U1185 ( .A1(n1330), .A2(n1331), .ZN(n1024) );
  NOR2_X1 U1186 ( .A1(n1002), .A2(n1148), .ZN(n1035) );
  NOR2_X1 U1187 ( .A1(n1380), .A2(G169), .ZN(n1128) );
  XNOR2_X1 U1188 ( .A(n1122), .B(n1056), .ZN(n1036) );
  NAND2_X1 U1189 ( .A1(n1043), .A2(n1042), .ZN(n1041) );
  XNOR2_X1 U1190 ( .A(n1893), .B(n1892), .ZN(n1042) );
  NOR2_X1 U1191 ( .A1(n1373), .A2(n1880), .ZN(n1657) );
  NAND2_X1 U1192 ( .A1(n1046), .A2(n1044), .ZN(n1668) );
  INV_X1 U1193 ( .A(n1373), .ZN(n1046) );
  NAND2_X1 U1194 ( .A1(n1307), .A2(n1048), .ZN(n1050) );
  NAND2_X1 U1195 ( .A1(n1050), .A2(n1049), .ZN(n1311) );
  AND2_X1 U1196 ( .A1(n1817), .A2(n1816), .ZN(n1052) );
  NAND2_X1 U1197 ( .A1(n1323), .A2(n1058), .ZN(n1057) );
  NOR2_X1 U1198 ( .A1(n1337), .A2(n1061), .ZN(n1058) );
  NAND2_X1 U1199 ( .A1(n1337), .A2(n1061), .ZN(n1060) );
  NAND2_X1 U1200 ( .A1(n1063), .A2(n1337), .ZN(n1062) );
  INV_X1 U1201 ( .A(n1323), .ZN(n1063) );
  NAND2_X1 U1202 ( .A1(n1323), .A2(n1064), .ZN(n2007) );
  NAND2_X1 U1203 ( .A1(n1363), .A2(n1765), .ZN(n1065) );
  INV_X1 U1204 ( .A(n1066), .ZN(n1415) );
  NOR2_X1 U1205 ( .A1(n1765), .A2(n1246), .ZN(n1067) );
  XNOR2_X2 U1206 ( .A(n2007), .B(n1070), .ZN(n1401) );
  NAND2_X1 U1207 ( .A1(n1094), .A2(n1325), .ZN(n1074) );
  INV_X1 U1208 ( .A(n1817), .ZN(n1078) );
  XNOR2_X1 U1209 ( .A(n1747), .B(n1076), .ZN(n1080) );
  NAND2_X1 U1210 ( .A1(n1079), .A2(n1008), .ZN(n1092) );
  NAND2_X1 U1211 ( .A1(n1078), .A2(n2014), .ZN(n1077) );
  NAND2_X1 U1212 ( .A1(n1080), .A2(n2014), .ZN(n1079) );
  NAND2_X1 U1213 ( .A1(n1082), .A2(n1081), .ZN(n1671) );
  INV_X1 U1214 ( .A(n1085), .ZN(n1888) );
  INV_X1 U1215 ( .A(n1372), .ZN(n1885) );
  NOR2_X1 U1216 ( .A1(n1381), .A2(n1605), .ZN(n1086) );
  NAND2_X1 U1217 ( .A1(n1669), .A2(n1886), .ZN(n1089) );
  AND2_X1 U1218 ( .A1(n1669), .A2(n1088), .ZN(n1730) );
  NAND2_X1 U1219 ( .A1(n1089), .A2(n1672), .ZN(n1680) );
  NAND2_X1 U1220 ( .A1(n2018), .A2(n1757), .ZN(n1093) );
  AND2_X2 U1221 ( .A1(n1092), .A2(n1090), .ZN(G375) );
  NAND2_X1 U1222 ( .A1(n1091), .A2(n1815), .ZN(n1090) );
  NAND2_X1 U1223 ( .A1(n1342), .A2(n1341), .ZN(n1099) );
  INV_X1 U1224 ( .A(n1341), .ZN(n1098) );
  XNOR2_X1 U1225 ( .A(n1099), .B(n1878), .ZN(n1879) );
  NAND2_X1 U1226 ( .A1(n1006), .A2(n1100), .ZN(n1587) );
  NAND2_X1 U1227 ( .A1(n1121), .A2(n1102), .ZN(n1101) );
  NAND2_X1 U1228 ( .A1(n1121), .A2(G33), .ZN(n1129) );
  NOR2_X1 U1229 ( .A1(n1951), .A2(n1388), .ZN(n1391) );
  NOR2_X1 U1230 ( .A1(n1298), .A2(n1522), .ZN(n1104) );
  OR2_X1 U1231 ( .A1(n1587), .A2(n1687), .ZN(n1105) );
  AND2_X1 U1232 ( .A1(n1608), .A2(n1607), .ZN(n1106) );
  XOR2_X1 U1233 ( .A(KEYINPUT36), .B(n1615), .Z(n1107) );
  AND2_X1 U1234 ( .A1(n1611), .A2(G264), .ZN(n1108) );
  AND2_X1 U1235 ( .A1(n1586), .A2(n1585), .ZN(n1109) );
  AND2_X1 U1236 ( .A1(n1868), .A2(n1867), .ZN(n1110) );
  INV_X1 U1237 ( .A(KEYINPUT64), .ZN(n1312) );
  INV_X1 U1238 ( .A(n1951), .ZN(n1878) );
  XNOR2_X1 U1239 ( .A(n1313), .B(n1312), .ZN(n1314) );
  XNOR2_X1 U1240 ( .A(n1743), .B(KEYINPUT68), .ZN(n1744) );
  NAND2_X1 U1241 ( .A1(n1610), .A2(n1728), .ZN(n1676) );
  INV_X1 U1242 ( .A(G384), .ZN(n1959) );
  XNOR2_X1 U1243 ( .A(G390), .B(n1959), .ZN(n1960) );
  NOR2_X1 U1244 ( .A1(G13), .A2(G33), .ZN(n1821) );
  INV_X1 U1245 ( .A(G87), .ZN(n1508) );
  NOR2_X1 U1246 ( .A1(G97), .A2(G107), .ZN(n1509) );
  OR2_X1 U1247 ( .A1(n1508), .A2(n1509), .ZN(G355) );
  NAND2_X1 U1248 ( .A1(n1155), .A2(G13), .ZN(n1146) );
  NOR2_X1 U1249 ( .A1(n1199), .A2(n1146), .ZN(n1112) );
  NOR2_X1 U1250 ( .A1(n2017), .A2(n1112), .ZN(n1113) );
  NOR2_X1 U1251 ( .A1(n2017), .A2(n1155), .ZN(n2002) );
  INV_X1 U1252 ( .A(G13), .ZN(n1114) );
  NAND2_X1 U1253 ( .A1(n2002), .A2(n1114), .ZN(n1979) );
  INV_X1 U1254 ( .A(n2014), .ZN(n1818) );
  NAND2_X1 U1255 ( .A1(n1820), .A2(n1818), .ZN(n1876) );
  INV_X1 U1256 ( .A(n1876), .ZN(n1902) );
  XNOR2_X1 U1257 ( .A(G330), .B(KEYINPUT95), .ZN(n1153) );
  XOR2_X1 U1258 ( .A(KEYINPUT10), .B(KEYINPUT76), .Z(n1119) );
  INV_X1 U1259 ( .A(G41), .ZN(n1765) );
  XNOR2_X2 U1260 ( .A(n1117), .B(n1116), .ZN(n1309) );
  NAND2_X1 U1261 ( .A1(G270), .A2(n1309), .ZN(n1118) );
  INV_X1 U1262 ( .A(G1698), .ZN(n1120) );
  NAND2_X1 U1263 ( .A1(G303), .A2(n1307), .ZN(n1122) );
  NAND2_X1 U1264 ( .A1(G274), .A2(n1123), .ZN(n1315) );
  NAND2_X1 U1265 ( .A1(n1614), .A2(G257), .ZN(n1124) );
  NAND2_X1 U1266 ( .A1(n1315), .A2(n1124), .ZN(n1125) );
  INV_X1 U1267 ( .A(G179), .ZN(n1126) );
  NOR2_X1 U1268 ( .A1(n1128), .A2(n1127), .ZN(n1143) );
  NAND2_X1 U1269 ( .A1(G283), .A2(n1626), .ZN(n1131) );
  NAND2_X1 U1270 ( .A1(n1622), .A2(G97), .ZN(n1130) );
  NAND2_X1 U1271 ( .A1(n1131), .A2(n1130), .ZN(n1133) );
  NOR2_X1 U1272 ( .A1(n1155), .A2(G1), .ZN(n1421) );
  NAND2_X1 U1273 ( .A1(G13), .A2(n1421), .ZN(n1424) );
  NOR2_X1 U1274 ( .A1(G116), .A2(n1424), .ZN(n1132) );
  NOR2_X1 U1275 ( .A1(n1133), .A2(n1132), .ZN(n1142) );
  NOR2_X1 U1276 ( .A1(G1), .A2(n1246), .ZN(n1298) );
  NAND2_X1 U1277 ( .A1(G20), .A2(G33), .ZN(n1134) );
  XOR2_X1 U1278 ( .A(KEYINPUT3), .B(KEYINPUT72), .Z(n1135) );
  XNOR2_X1 U1279 ( .A(n1136), .B(n1135), .ZN(n1137) );
  NAND2_X1 U1280 ( .A1(n1138), .A2(n1137), .ZN(n1420) );
  NOR2_X1 U1281 ( .A1(n1298), .A2(n1297), .ZN(n1265) );
  NAND2_X1 U1282 ( .A1(n1420), .A2(G20), .ZN(n1140) );
  NOR2_X1 U1283 ( .A1(n1265), .A2(n1633), .ZN(n1346) );
  OR2_X1 U1284 ( .A1(n1016), .A2(n1346), .ZN(n1141) );
  NAND2_X1 U1285 ( .A1(n1142), .A2(n1141), .ZN(n1148) );
  INV_X1 U1286 ( .A(n1380), .ZN(n1144) );
  NAND2_X1 U1287 ( .A1(G200), .A2(n1144), .ZN(n1145) );
  INV_X1 U1288 ( .A(G213), .ZN(n1976) );
  OR2_X1 U1289 ( .A1(n1976), .A2(n1146), .ZN(n1147) );
  NOR2_X1 U1290 ( .A1(G1), .A2(n1147), .ZN(n1761) );
  AND2_X1 U1291 ( .A1(n1148), .A2(n1881), .ZN(n1149) );
  NOR2_X1 U1292 ( .A1(n1388), .A2(n1149), .ZN(n1151) );
  INV_X1 U1293 ( .A(n1332), .ZN(n1320) );
  NOR2_X1 U1294 ( .A1(n1320), .A2(n1886), .ZN(n1150) );
  XNOR2_X1 U1295 ( .A(n1153), .B(n1323), .ZN(n1154) );
  NOR2_X1 U1296 ( .A1(n1902), .A2(n1154), .ZN(n1216) );
  NAND2_X1 U1297 ( .A1(n1821), .A2(n1155), .ZN(n1547) );
  NOR2_X1 U1298 ( .A1(G190), .A2(n1155), .ZN(n1159) );
  NAND2_X1 U1299 ( .A1(G200), .A2(n1159), .ZN(n1156) );
  NAND2_X1 U1300 ( .A1(G317), .A2(n1927), .ZN(n1158) );
  NOR2_X1 U1301 ( .A1(G179), .A2(n1156), .ZN(n1844) );
  NAND2_X1 U1302 ( .A1(n1844), .A2(G283), .ZN(n1157) );
  NAND2_X1 U1303 ( .A1(n1158), .A2(n1157), .ZN(n1165) );
  INV_X1 U1304 ( .A(G200), .ZN(n1639) );
  NAND2_X1 U1305 ( .A1(n1159), .A2(n1639), .ZN(n1171) );
  NAND2_X1 U1306 ( .A1(n1933), .A2(G329), .ZN(n1162) );
  INV_X1 U1307 ( .A(G190), .ZN(n1432) );
  NOR2_X1 U1308 ( .A1(G200), .A2(n1432), .ZN(n1176) );
  NAND2_X1 U1309 ( .A1(n1176), .A2(n1126), .ZN(n1160) );
  NAND2_X1 U1310 ( .A1(G20), .A2(n1160), .ZN(n1909) );
  NAND2_X1 U1311 ( .A1(G294), .A2(n1909), .ZN(n1161) );
  NAND2_X1 U1312 ( .A1(n1162), .A2(n1161), .ZN(n1163) );
  XOR2_X1 U1313 ( .A(KEYINPUT93), .B(n1163), .Z(n1164) );
  NOR2_X1 U1314 ( .A1(n1165), .A2(n1164), .ZN(n1166) );
  XNOR2_X1 U1315 ( .A(n1166), .B(KEYINPUT94), .ZN(n1170) );
  NOR2_X1 U1316 ( .A1(n1432), .A2(n1639), .ZN(n1167) );
  AND2_X1 U1317 ( .A1(G20), .A2(n1167), .ZN(n1178) );
  NAND2_X1 U1318 ( .A1(n1178), .A2(G179), .ZN(n1168) );
  NAND2_X1 U1319 ( .A1(G326), .A2(n1926), .ZN(n1169) );
  NAND2_X1 U1320 ( .A1(n1170), .A2(n1169), .ZN(n1174) );
  NAND2_X1 U1321 ( .A1(n1931), .A2(G311), .ZN(n1172) );
  XOR2_X1 U1322 ( .A(KEYINPUT92), .B(n1172), .Z(n1173) );
  NOR2_X1 U1323 ( .A1(n1174), .A2(n1173), .ZN(n1183) );
  INV_X1 U1324 ( .A(G169), .ZN(n1605) );
  NAND2_X1 U1325 ( .A1(G20), .A2(n1605), .ZN(n1175) );
  NAND2_X1 U1326 ( .A1(n1121), .A2(n1175), .ZN(n1197) );
  INV_X1 U1327 ( .A(n1197), .ZN(n1766) );
  NAND2_X1 U1328 ( .A1(G33), .A2(n1766), .ZN(n1829) );
  NAND2_X1 U1329 ( .A1(G20), .A2(n1176), .ZN(n1177) );
  NAND2_X1 U1330 ( .A1(G322), .A2(n1934), .ZN(n1180) );
  NAND2_X1 U1331 ( .A1(n1126), .A2(n1178), .ZN(n1924) );
  INV_X1 U1332 ( .A(n1924), .ZN(n1912) );
  NAND2_X1 U1333 ( .A1(n1912), .A2(G303), .ZN(n1179) );
  NAND2_X1 U1334 ( .A1(n1180), .A2(n1179), .ZN(n1181) );
  NOR2_X1 U1335 ( .A1(n1829), .A2(n1181), .ZN(n1182) );
  NAND2_X1 U1336 ( .A1(n1926), .A2(G50), .ZN(n1196) );
  NOR2_X1 U1337 ( .A1(G33), .A2(n1197), .ZN(n1946) );
  NAND2_X1 U1338 ( .A1(G107), .A2(n1844), .ZN(n1224) );
  NAND2_X1 U1339 ( .A1(n1946), .A2(n1224), .ZN(n1194) );
  NAND2_X1 U1340 ( .A1(n1927), .A2(G68), .ZN(n1188) );
  INV_X1 U1341 ( .A(n1909), .ZN(n1709) );
  INV_X1 U1342 ( .A(G97), .ZN(n1687) );
  NOR2_X1 U1343 ( .A1(n1709), .A2(n1687), .ZN(n1475) );
  NAND2_X1 U1344 ( .A1(n1933), .A2(G159), .ZN(n1185) );
  NAND2_X1 U1345 ( .A1(n1931), .A2(G77), .ZN(n1184) );
  NAND2_X1 U1346 ( .A1(n1185), .A2(n1184), .ZN(n1186) );
  NOR2_X1 U1347 ( .A1(n1475), .A2(n1186), .ZN(n1187) );
  NAND2_X1 U1348 ( .A1(n1188), .A2(n1187), .ZN(n1189) );
  XNOR2_X1 U1349 ( .A(n1189), .B(KEYINPUT61), .ZN(n1192) );
  NOR2_X1 U1350 ( .A1(n1508), .A2(n1924), .ZN(n1825) );
  AND2_X1 U1351 ( .A1(n1934), .A2(G58), .ZN(n1190) );
  NOR2_X1 U1352 ( .A1(n1825), .A2(n1190), .ZN(n1191) );
  NAND2_X1 U1353 ( .A1(n1192), .A2(n1191), .ZN(n1193) );
  NOR2_X1 U1354 ( .A1(n1194), .A2(n1193), .ZN(n1195) );
  NAND2_X1 U1355 ( .A1(n1196), .A2(n1195), .ZN(n1213) );
  NAND2_X1 U1356 ( .A1(n1197), .A2(n1547), .ZN(n1899) );
  XNOR2_X1 U1357 ( .A(G50), .B(G77), .ZN(n1198) );
  XNOR2_X1 U1358 ( .A(G68), .B(G58), .ZN(n1562) );
  XNOR2_X1 U1359 ( .A(n1198), .B(n1562), .ZN(n2043) );
  NAND2_X1 U1360 ( .A1(G45), .A2(n2043), .ZN(n1201) );
  NOR2_X1 U1361 ( .A1(G68), .A2(G58), .ZN(n1632) );
  INV_X1 U1362 ( .A(G50), .ZN(n1767) );
  NOR2_X1 U1363 ( .A1(n1632), .A2(n1767), .ZN(n2013) );
  NAND2_X1 U1364 ( .A1(n2013), .A2(n1199), .ZN(n1200) );
  NAND2_X1 U1365 ( .A1(n1201), .A2(n1200), .ZN(n1202) );
  XOR2_X1 U1366 ( .A(KEYINPUT90), .B(n1202), .Z(n1204) );
  NOR2_X1 U1367 ( .A1(n1979), .A2(n1246), .ZN(n1203) );
  XNOR2_X1 U1368 ( .A(n1203), .B(KEYINPUT24), .ZN(n1896) );
  NAND2_X1 U1369 ( .A1(n1204), .A2(n1896), .ZN(n1206) );
  NAND2_X1 U1370 ( .A1(n1821), .A2(G355), .ZN(n1205) );
  NAND2_X1 U1371 ( .A1(n1206), .A2(n1205), .ZN(n1209) );
  NAND2_X1 U1372 ( .A1(n1016), .A2(n1979), .ZN(n1207) );
  XOR2_X1 U1373 ( .A(KEYINPUT60), .B(n1207), .Z(n1208) );
  NOR2_X1 U1374 ( .A1(n1209), .A2(n1208), .ZN(n1210) );
  NOR2_X1 U1375 ( .A1(n1899), .A2(n1210), .ZN(n1211) );
  XNOR2_X1 U1376 ( .A(n1211), .B(KEYINPUT91), .ZN(n1212) );
  NAND2_X1 U1377 ( .A1(n1213), .A2(n1212), .ZN(n1214) );
  NOR2_X1 U1378 ( .A1(n1876), .A2(n1005), .ZN(n1215) );
  NOR2_X1 U1379 ( .A1(n1216), .A2(n1215), .ZN(G396) );
  NAND2_X1 U1380 ( .A1(n1934), .A2(G311), .ZN(n1217) );
  NAND2_X1 U1381 ( .A1(G33), .A2(n1217), .ZN(n1227) );
  NAND2_X1 U1382 ( .A1(G322), .A2(n1933), .ZN(n1219) );
  NAND2_X1 U1383 ( .A1(n1931), .A2(G294), .ZN(n1218) );
  NAND2_X1 U1384 ( .A1(n1219), .A2(n1218), .ZN(n1223) );
  NAND2_X1 U1385 ( .A1(G303), .A2(n1927), .ZN(n1221) );
  NAND2_X1 U1386 ( .A1(G116), .A2(n1909), .ZN(n1220) );
  NAND2_X1 U1387 ( .A1(n1221), .A2(n1220), .ZN(n1222) );
  NOR2_X1 U1388 ( .A1(n1223), .A2(n1222), .ZN(n1225) );
  NAND2_X1 U1389 ( .A1(n1225), .A2(n1224), .ZN(n1226) );
  NOR2_X1 U1390 ( .A1(n1227), .A2(n1226), .ZN(n1228) );
  XNOR2_X1 U1391 ( .A(n1228), .B(KEYINPUT58), .ZN(n1234) );
  XNOR2_X1 U1392 ( .A(KEYINPUT88), .B(KEYINPUT59), .ZN(n1232) );
  NAND2_X1 U1393 ( .A1(G317), .A2(n1926), .ZN(n1230) );
  NAND2_X1 U1394 ( .A1(n1912), .A2(G283), .ZN(n1229) );
  NAND2_X1 U1395 ( .A1(n1230), .A2(n1229), .ZN(n1231) );
  XNOR2_X1 U1396 ( .A(n1232), .B(n1231), .ZN(n1233) );
  NAND2_X1 U1397 ( .A1(n1234), .A2(n1233), .ZN(n1253) );
  NAND2_X1 U1398 ( .A1(n1931), .A2(G58), .ZN(n1236) );
  NAND2_X1 U1399 ( .A1(n1927), .A2(G50), .ZN(n1235) );
  NAND2_X1 U1400 ( .A1(n1236), .A2(n1235), .ZN(n1242) );
  NAND2_X1 U1401 ( .A1(G150), .A2(n1926), .ZN(n1237) );
  XNOR2_X1 U1402 ( .A(n1237), .B(KEYINPUT56), .ZN(n1239) );
  NAND2_X1 U1403 ( .A1(n1912), .A2(G68), .ZN(n1238) );
  NAND2_X1 U1404 ( .A1(n1239), .A2(n1238), .ZN(n1240) );
  XOR2_X1 U1405 ( .A(KEYINPUT57), .B(n1240), .Z(n1241) );
  NOR2_X1 U1406 ( .A1(n1242), .A2(n1241), .ZN(n1251) );
  INV_X1 U1407 ( .A(G77), .ZN(n2030) );
  NOR2_X1 U1408 ( .A1(n1709), .A2(n2030), .ZN(n1826) );
  NAND2_X1 U1409 ( .A1(G143), .A2(n1933), .ZN(n1244) );
  NAND2_X1 U1410 ( .A1(n1934), .A2(G159), .ZN(n1243) );
  NAND2_X1 U1411 ( .A1(n1244), .A2(n1243), .ZN(n1245) );
  NOR2_X1 U1412 ( .A1(n1826), .A2(n1245), .ZN(n1247) );
  NAND2_X1 U1413 ( .A1(n1247), .A2(n1246), .ZN(n1249) );
  NAND2_X1 U1414 ( .A1(n1844), .A2(G87), .ZN(n1248) );
  XOR2_X1 U1415 ( .A(KEYINPUT22), .B(n1248), .Z(n1479) );
  NOR2_X1 U1416 ( .A1(n1249), .A2(n1479), .ZN(n1250) );
  NAND2_X1 U1417 ( .A1(n1251), .A2(n1250), .ZN(n1252) );
  NAND2_X1 U1418 ( .A1(n1253), .A2(n1252), .ZN(n1254) );
  NAND2_X1 U1419 ( .A1(n1766), .A2(n1254), .ZN(n1255) );
  XNOR2_X1 U1420 ( .A(KEYINPUT89), .B(n1255), .ZN(n1256) );
  NOR2_X1 U1421 ( .A1(n1876), .A2(n1256), .ZN(n1288) );
  INV_X1 U1422 ( .A(n1547), .ZN(n1952) );
  NAND2_X1 U1423 ( .A1(G244), .A2(n1614), .ZN(n1258) );
  NAND2_X1 U1424 ( .A1(G250), .A2(n1611), .ZN(n1257) );
  NAND2_X1 U1425 ( .A1(n1258), .A2(n1257), .ZN(n1261) );
  NAND2_X1 U1426 ( .A1(n1307), .A2(G283), .ZN(n1259) );
  NAND2_X1 U1427 ( .A1(n1315), .A2(n1259), .ZN(n1260) );
  XNOR2_X1 U1428 ( .A(n1262), .B(KEYINPUT12), .ZN(n1264) );
  NAND2_X1 U1429 ( .A1(G257), .A2(n1309), .ZN(n1263) );
  NAND2_X1 U1430 ( .A1(n1264), .A2(n1263), .ZN(n1377) );
  NAND2_X1 U1431 ( .A1(n1377), .A2(G200), .ZN(n1278) );
  NOR2_X1 U1432 ( .A1(n1432), .A2(n1377), .ZN(n1276) );
  NAND2_X1 U1433 ( .A1(G77), .A2(n1622), .ZN(n1267) );
  NAND2_X1 U1434 ( .A1(n1265), .A2(G97), .ZN(n1266) );
  NAND2_X1 U1435 ( .A1(n1267), .A2(n1266), .ZN(n1270) );
  INV_X1 U1436 ( .A(n1304), .ZN(n1343) );
  XOR2_X1 U1437 ( .A(G97), .B(G107), .Z(n1268) );
  XNOR2_X1 U1438 ( .A(KEYINPUT80), .B(n1268), .ZN(n2038) );
  NOR2_X1 U1439 ( .A1(n1343), .A2(n2038), .ZN(n1269) );
  NOR2_X1 U1440 ( .A1(n1270), .A2(n1269), .ZN(n1275) );
  INV_X1 U1441 ( .A(G107), .ZN(n1522) );
  XNOR2_X1 U1442 ( .A(n1626), .B(KEYINPUT81), .ZN(n1423) );
  NOR2_X1 U1443 ( .A1(n1522), .A2(n1423), .ZN(n1272) );
  NOR2_X1 U1444 ( .A1(G97), .A2(n1424), .ZN(n1271) );
  NOR2_X1 U1445 ( .A1(n1272), .A2(n1271), .ZN(n1273) );
  XOR2_X1 U1446 ( .A(KEYINPUT13), .B(n1273), .Z(n1274) );
  NAND2_X1 U1447 ( .A1(n1275), .A2(n1274), .ZN(n1283) );
  NOR2_X1 U1448 ( .A1(n1276), .A2(n1283), .ZN(n1277) );
  NAND2_X1 U1449 ( .A1(n1278), .A2(n1277), .ZN(n1282) );
  NOR2_X1 U1450 ( .A1(G179), .A2(n1377), .ZN(n1280) );
  AND2_X1 U1451 ( .A1(n1605), .A2(n1377), .ZN(n1279) );
  NOR2_X1 U1452 ( .A1(n1280), .A2(n1279), .ZN(n1281) );
  NAND2_X1 U1453 ( .A1(n1283), .A2(n1881), .ZN(n1284) );
  XOR2_X1 U1454 ( .A(KEYINPUT82), .B(n1284), .Z(n1322) );
  NOR2_X1 U1455 ( .A1(n1389), .A2(n1322), .ZN(n1286) );
  NOR2_X1 U1456 ( .A1(n1341), .A2(n1886), .ZN(n1285) );
  NOR2_X1 U1457 ( .A1(n1286), .A2(n1285), .ZN(n1891) );
  NAND2_X1 U1458 ( .A1(n1952), .A2(n1891), .ZN(n1287) );
  NAND2_X1 U1459 ( .A1(n1288), .A2(n1287), .ZN(n1296) );
  NAND2_X1 U1460 ( .A1(G97), .A2(n1979), .ZN(n1289) );
  XNOR2_X1 U1461 ( .A(n1289), .B(KEYINPUT86), .ZN(n1293) );
  XNOR2_X1 U1462 ( .A(n2038), .B(KEYINPUT51), .ZN(n1291) );
  XNOR2_X1 U1463 ( .A(G87), .B(G116), .ZN(n1290) );
  XNOR2_X1 U1464 ( .A(n1291), .B(n1290), .ZN(n2044) );
  NAND2_X1 U1465 ( .A1(n2044), .A2(n1896), .ZN(n1292) );
  NAND2_X1 U1466 ( .A1(n1293), .A2(n1292), .ZN(n1294) );
  NOR2_X1 U1467 ( .A1(n1899), .A2(n1294), .ZN(n1295) );
  NOR2_X1 U1468 ( .A1(n1296), .A2(n1295), .ZN(n1399) );
  XNOR2_X1 U1469 ( .A(n1297), .B(KEYINPUT73), .ZN(n1299) );
  NAND2_X1 U1470 ( .A1(n1299), .A2(n1104), .ZN(n1300) );
  NAND2_X1 U1471 ( .A1(n1301), .A2(n1300), .ZN(n1302) );
  XNOR2_X1 U1472 ( .A(n1302), .B(KEYINPUT17), .ZN(n1303) );
  NOR2_X1 U1473 ( .A1(n1304), .A2(n1623), .ZN(n1594) );
  NOR2_X1 U1474 ( .A1(n1594), .A2(G107), .ZN(n1305) );
  XNOR2_X1 U1475 ( .A(n1305), .B(KEYINPUT74), .ZN(n1306) );
  INV_X1 U1476 ( .A(KEYINPUT14), .ZN(n1308) );
  NAND2_X1 U1477 ( .A1(n1309), .A2(G264), .ZN(n1310) );
  AND2_X1 U1478 ( .A1(n1314), .A2(G250), .ZN(n1316) );
  NAND2_X1 U1479 ( .A1(G200), .A2(n1378), .ZN(n1319) );
  INV_X1 U1480 ( .A(n1378), .ZN(n1374) );
  NAND2_X1 U1481 ( .A1(G190), .A2(n1374), .ZN(n1318) );
  NOR2_X1 U1482 ( .A1(n1321), .A2(n1324), .ZN(n1339) );
  NAND2_X1 U1483 ( .A1(n1881), .A2(n1324), .ZN(n1331) );
  NOR2_X1 U1484 ( .A1(n1886), .A2(n1325), .ZN(n1326) );
  XNOR2_X1 U1485 ( .A(n1326), .B(KEYINPUT75), .ZN(n1333) );
  BUF_X1 U1486 ( .A(n1327), .Z(n1328) );
  NAND2_X1 U1487 ( .A1(n1333), .A2(n1329), .ZN(n1330) );
  NAND2_X1 U1488 ( .A1(n1886), .A2(n1332), .ZN(n1334) );
  NAND2_X1 U1489 ( .A1(n1334), .A2(n1333), .ZN(n1335) );
  XNOR2_X1 U1490 ( .A(n1335), .B(KEYINPUT78), .ZN(n1336) );
  NAND2_X1 U1491 ( .A1(n1401), .A2(n1551), .ZN(n1338) );
  INV_X1 U1492 ( .A(n1401), .ZN(n1395) );
  NOR2_X1 U1493 ( .A1(n1339), .A2(n1389), .ZN(n1340) );
  XNOR2_X1 U1494 ( .A(n1340), .B(KEYINPUT83), .ZN(n1342) );
  NOR2_X1 U1495 ( .A1(G87), .A2(n1424), .ZN(n1351) );
  NOR2_X1 U1496 ( .A1(n1343), .A2(n1509), .ZN(n1344) );
  NOR2_X1 U1497 ( .A1(G87), .A2(n1344), .ZN(n1345) );
  XNOR2_X1 U1498 ( .A(n1347), .B(KEYINPUT9), .ZN(n1349) );
  NAND2_X1 U1499 ( .A1(n1622), .A2(G68), .ZN(n1348) );
  NAND2_X1 U1500 ( .A1(n1349), .A2(n1348), .ZN(n1350) );
  NOR2_X1 U1501 ( .A1(n1351), .A2(n1350), .ZN(n1353) );
  NAND2_X1 U1502 ( .A1(G97), .A2(n1626), .ZN(n1352) );
  NAND2_X1 U1503 ( .A1(n1363), .A2(G274), .ZN(n1355) );
  NAND2_X1 U1504 ( .A1(G116), .A2(n1307), .ZN(n1354) );
  NAND2_X1 U1505 ( .A1(n1355), .A2(n1354), .ZN(n1362) );
  NAND2_X1 U1506 ( .A1(G244), .A2(n1611), .ZN(n1357) );
  NAND2_X1 U1507 ( .A1(n1614), .A2(G238), .ZN(n1356) );
  NAND2_X1 U1508 ( .A1(n1357), .A2(n1356), .ZN(n1360) );
  NOR2_X1 U1509 ( .A1(n1362), .A2(n1361), .ZN(n1367) );
  NAND2_X1 U1510 ( .A1(G250), .A2(n1066), .ZN(n1364) );
  NOR2_X1 U1511 ( .A1(n1364), .A2(n1363), .ZN(n1365) );
  XOR2_X1 U1512 ( .A(KEYINPUT84), .B(n1365), .Z(n1366) );
  NAND2_X1 U1513 ( .A1(n1367), .A2(n1366), .ZN(n1375) );
  INV_X1 U1514 ( .A(n1375), .ZN(n1381) );
  NOR2_X1 U1515 ( .A1(n1126), .A2(n1375), .ZN(n1368) );
  NAND2_X1 U1516 ( .A1(G200), .A2(n1375), .ZN(n1370) );
  NAND2_X1 U1517 ( .A1(G190), .A2(n1381), .ZN(n1369) );
  NAND2_X1 U1518 ( .A1(n1370), .A2(n1369), .ZN(n1371) );
  NAND2_X1 U1519 ( .A1(n1657), .A2(n1886), .ZN(n1393) );
  NAND2_X1 U1520 ( .A1(G179), .A2(n1374), .ZN(n1376) );
  NAND2_X1 U1521 ( .A1(n1378), .A2(n1377), .ZN(n1379) );
  NOR2_X1 U1522 ( .A1(n1380), .A2(n1379), .ZN(n1383) );
  NOR2_X1 U1523 ( .A1(n1381), .A2(G179), .ZN(n1382) );
  NAND2_X1 U1524 ( .A1(n1383), .A2(n1382), .ZN(n1384) );
  NAND2_X1 U1525 ( .A1(n1385), .A2(n1384), .ZN(n1386) );
  NAND2_X1 U1526 ( .A1(n1391), .A2(n1390), .ZN(n2005) );
  NAND2_X1 U1527 ( .A1(n1393), .A2(n1671), .ZN(n1873) );
  INV_X1 U1528 ( .A(n1873), .ZN(n2008) );
  NAND2_X1 U1529 ( .A1(n2008), .A2(n1551), .ZN(n1394) );
  NAND2_X1 U1530 ( .A1(n1395), .A2(n1394), .ZN(n1396) );
  NAND2_X1 U1531 ( .A1(n1875), .A2(n1396), .ZN(n1397) );
  NOR2_X1 U1532 ( .A1(n1397), .A2(n1818), .ZN(n1398) );
  NOR2_X1 U1533 ( .A1(n1399), .A2(n1398), .ZN(n1404) );
  NAND2_X1 U1534 ( .A1(n2014), .A2(n1873), .ZN(n1400) );
  NAND2_X1 U1535 ( .A1(n1820), .A2(n1400), .ZN(n1402) );
  NAND2_X1 U1536 ( .A1(n1402), .A2(n1401), .ZN(n1403) );
  NAND2_X1 U1537 ( .A1(n1404), .A2(n1403), .ZN(G390) );
  NAND2_X1 U1538 ( .A1(n1307), .A2(G107), .ZN(n1406) );
  NAND2_X1 U1539 ( .A1(G232), .A2(n1614), .ZN(n1405) );
  NAND2_X1 U1540 ( .A1(n1406), .A2(n1405), .ZN(n1409) );
  NAND2_X1 U1541 ( .A1(G238), .A2(n1611), .ZN(n1407) );
  XOR2_X1 U1542 ( .A(KEYINPUT6), .B(n1407), .Z(n1408) );
  NOR2_X1 U1543 ( .A1(n1409), .A2(n1408), .ZN(n1412) );
  NOR2_X1 U1544 ( .A1(G41), .A2(G45), .ZN(n1410) );
  XNOR2_X1 U1545 ( .A(n1410), .B(KEYINPUT96), .ZN(n1411) );
  NOR2_X1 U1546 ( .A1(G1), .A2(n1411), .ZN(n1414) );
  NAND2_X1 U1547 ( .A1(n1414), .A2(G274), .ZN(n1613) );
  NAND2_X1 U1548 ( .A1(n1412), .A2(n1613), .ZN(n1413) );
  XNOR2_X1 U1549 ( .A(n1413), .B(KEYINPUT7), .ZN(n1417) );
  NOR2_X1 U1550 ( .A1(n1415), .A2(n1414), .ZN(n1617) );
  NAND2_X1 U1551 ( .A1(G244), .A2(n1617), .ZN(n1416) );
  NAND2_X1 U1552 ( .A1(n1417), .A2(n1416), .ZN(n1434) );
  NAND2_X1 U1553 ( .A1(G169), .A2(n1434), .ZN(n1419) );
  OR2_X1 U1554 ( .A1(n1126), .A2(n1434), .ZN(n1418) );
  NAND2_X1 U1555 ( .A1(n1419), .A2(n1418), .ZN(n1439) );
  NOR2_X1 U1556 ( .A1(n1421), .A2(n1420), .ZN(n1627) );
  NOR2_X1 U1557 ( .A1(n1627), .A2(n1633), .ZN(n1422) );
  NOR2_X1 U1558 ( .A1(n2030), .A2(n1422), .ZN(n1429) );
  NOR2_X1 U1559 ( .A1(n1508), .A2(n1423), .ZN(n1426) );
  NOR2_X1 U1560 ( .A1(G77), .A2(n1424), .ZN(n1425) );
  NOR2_X1 U1561 ( .A1(n1426), .A2(n1425), .ZN(n1427) );
  XNOR2_X1 U1562 ( .A(n1427), .B(KEYINPUT97), .ZN(n1428) );
  NOR2_X1 U1563 ( .A1(n1429), .A2(n1428), .ZN(n1431) );
  NAND2_X1 U1564 ( .A1(n1622), .A2(G58), .ZN(n1430) );
  NAND2_X1 U1565 ( .A1(n1431), .A2(n1430), .ZN(n1437) );
  NOR2_X1 U1566 ( .A1(n1432), .A2(n1434), .ZN(n1433) );
  NOR2_X1 U1567 ( .A1(n1433), .A2(n1437), .ZN(n1436) );
  NAND2_X1 U1568 ( .A1(G200), .A2(n1434), .ZN(n1435) );
  NAND2_X1 U1569 ( .A1(n1436), .A2(n1435), .ZN(n1666) );
  NAND2_X1 U1570 ( .A1(n1667), .A2(n1666), .ZN(n1653) );
  NAND2_X1 U1571 ( .A1(n1881), .A2(n1437), .ZN(n1438) );
  XOR2_X1 U1572 ( .A(KEYINPUT5), .B(n1438), .Z(n1440) );
  AND2_X1 U1573 ( .A1(n1653), .A2(n1440), .ZN(n1442) );
  NOR2_X1 U1574 ( .A1(n1440), .A2(n1439), .ZN(n1441) );
  NOR2_X1 U1575 ( .A1(n1442), .A2(n1441), .ZN(n1754) );
  INV_X1 U1576 ( .A(n1754), .ZN(n1670) );
  XNOR2_X1 U1577 ( .A(n1873), .B(n1670), .ZN(n1443) );
  NAND2_X1 U1578 ( .A1(n1443), .A2(n1876), .ZN(n1488) );
  NAND2_X1 U1579 ( .A1(G143), .A2(n1934), .ZN(n1444) );
  XOR2_X1 U1580 ( .A(KEYINPUT123), .B(n1444), .Z(n1445) );
  NAND2_X1 U1581 ( .A1(n1946), .A2(n1445), .ZN(n1455) );
  NAND2_X1 U1582 ( .A1(G137), .A2(n1926), .ZN(n1447) );
  NAND2_X1 U1583 ( .A1(n1931), .A2(G159), .ZN(n1446) );
  NAND2_X1 U1584 ( .A1(n1447), .A2(n1446), .ZN(n1448) );
  XNOR2_X1 U1585 ( .A(n1448), .B(KEYINPUT124), .ZN(n1450) );
  NOR2_X1 U1586 ( .A1(n1767), .A2(n1924), .ZN(n1449) );
  NOR2_X1 U1587 ( .A1(n1450), .A2(n1449), .ZN(n1452) );
  NAND2_X1 U1588 ( .A1(G58), .A2(n1909), .ZN(n1451) );
  NAND2_X1 U1589 ( .A1(n1452), .A2(n1451), .ZN(n1453) );
  XNOR2_X1 U1590 ( .A(KEYINPUT20), .B(n1453), .ZN(n1454) );
  NOR2_X1 U1591 ( .A1(n1455), .A2(n1454), .ZN(n1461) );
  NAND2_X1 U1592 ( .A1(G68), .A2(n1844), .ZN(n1823) );
  NAND2_X1 U1593 ( .A1(G150), .A2(n1927), .ZN(n1456) );
  NAND2_X1 U1594 ( .A1(n1823), .A2(n1456), .ZN(n1459) );
  NAND2_X1 U1595 ( .A1(n1933), .A2(G132), .ZN(n1457) );
  XNOR2_X1 U1596 ( .A(KEYINPUT19), .B(n1457), .ZN(n1458) );
  NOR2_X1 U1597 ( .A1(n1459), .A2(n1458), .ZN(n1460) );
  NAND2_X1 U1598 ( .A1(n1461), .A2(n1460), .ZN(n1463) );
  NOR2_X1 U1599 ( .A1(n1766), .A2(n1821), .ZN(n1861) );
  NAND2_X1 U1600 ( .A1(n1861), .A2(n2030), .ZN(n1462) );
  NAND2_X1 U1601 ( .A1(n1463), .A2(n1462), .ZN(n1464) );
  NOR2_X1 U1602 ( .A1(n1876), .A2(n1464), .ZN(n1483) );
  INV_X1 U1603 ( .A(n1829), .ZN(n1914) );
  NAND2_X1 U1604 ( .A1(G283), .A2(n1927), .ZN(n1465) );
  NAND2_X1 U1605 ( .A1(n1914), .A2(n1465), .ZN(n1472) );
  NAND2_X1 U1606 ( .A1(n1926), .A2(G303), .ZN(n1467) );
  NAND2_X1 U1607 ( .A1(n1934), .A2(G294), .ZN(n1466) );
  NAND2_X1 U1608 ( .A1(n1467), .A2(n1466), .ZN(n1469) );
  NOR2_X1 U1609 ( .A1(n1522), .A2(n1924), .ZN(n1468) );
  NOR2_X1 U1610 ( .A1(n1469), .A2(n1468), .ZN(n1470) );
  XOR2_X1 U1611 ( .A(KEYINPUT122), .B(n1470), .Z(n1471) );
  NOR2_X1 U1612 ( .A1(n1472), .A2(n1471), .ZN(n1481) );
  NAND2_X1 U1613 ( .A1(G116), .A2(n1931), .ZN(n1473) );
  XNOR2_X1 U1614 ( .A(KEYINPUT21), .B(n1473), .ZN(n1474) );
  NOR2_X1 U1615 ( .A1(n1475), .A2(n1474), .ZN(n1477) );
  NAND2_X1 U1616 ( .A1(n1933), .A2(G311), .ZN(n1476) );
  NAND2_X1 U1617 ( .A1(n1477), .A2(n1476), .ZN(n1478) );
  NOR2_X1 U1618 ( .A1(n1479), .A2(n1478), .ZN(n1480) );
  NAND2_X1 U1619 ( .A1(n1481), .A2(n1480), .ZN(n1482) );
  NAND2_X1 U1620 ( .A1(n1483), .A2(n1482), .ZN(n1484) );
  XNOR2_X1 U1621 ( .A(n1484), .B(KEYINPUT125), .ZN(n1486) );
  NAND2_X1 U1622 ( .A1(n1821), .A2(n1670), .ZN(n1485) );
  NAND2_X1 U1623 ( .A1(n1486), .A2(n1485), .ZN(n1487) );
  NAND2_X1 U1624 ( .A1(n1488), .A2(n1487), .ZN(G384) );
  NAND2_X1 U1625 ( .A1(G322), .A2(n1926), .ZN(n1490) );
  NAND2_X1 U1626 ( .A1(n1912), .A2(G294), .ZN(n1489) );
  NAND2_X1 U1627 ( .A1(n1490), .A2(n1489), .ZN(n1491) );
  XOR2_X1 U1628 ( .A(KEYINPUT26), .B(n1491), .Z(n1494) );
  NAND2_X1 U1629 ( .A1(n1844), .A2(G116), .ZN(n1492) );
  XOR2_X1 U1630 ( .A(KEYINPUT25), .B(n1492), .Z(n1493) );
  NAND2_X1 U1631 ( .A1(n1494), .A2(n1493), .ZN(n1506) );
  NAND2_X1 U1632 ( .A1(G317), .A2(n1934), .ZN(n1495) );
  XOR2_X1 U1633 ( .A(KEYINPUT116), .B(n1495), .Z(n1496) );
  NOR2_X1 U1634 ( .A1(n1829), .A2(n1496), .ZN(n1504) );
  NAND2_X1 U1635 ( .A1(n1927), .A2(G311), .ZN(n1498) );
  NAND2_X1 U1636 ( .A1(G283), .A2(n1909), .ZN(n1497) );
  NAND2_X1 U1637 ( .A1(n1498), .A2(n1497), .ZN(n1502) );
  NAND2_X1 U1638 ( .A1(G326), .A2(n1933), .ZN(n1500) );
  NAND2_X1 U1639 ( .A1(n1931), .A2(G303), .ZN(n1499) );
  NAND2_X1 U1640 ( .A1(n1500), .A2(n1499), .ZN(n1501) );
  NOR2_X1 U1641 ( .A1(n1502), .A2(n1501), .ZN(n1503) );
  NAND2_X1 U1642 ( .A1(n1504), .A2(n1503), .ZN(n1505) );
  NOR2_X1 U1643 ( .A1(n1506), .A2(n1505), .ZN(n1507) );
  NOR2_X1 U1644 ( .A1(n1876), .A2(n1507), .ZN(n1546) );
  NAND2_X1 U1645 ( .A1(n1509), .A2(n1508), .ZN(n1510) );
  NOR2_X1 U1646 ( .A1(G116), .A2(n1510), .ZN(n2009) );
  AND2_X1 U1647 ( .A1(G58), .A2(n2009), .ZN(n1512) );
  NAND2_X1 U1648 ( .A1(G68), .A2(G77), .ZN(n1511) );
  NAND2_X1 U1649 ( .A1(n1512), .A2(n1511), .ZN(n1513) );
  NOR2_X1 U1650 ( .A1(G50), .A2(n1513), .ZN(n1514) );
  NOR2_X1 U1651 ( .A1(G45), .A2(n1514), .ZN(n1516) );
  XOR2_X1 U1652 ( .A(KEYINPUT23), .B(KEYINPUT117), .Z(n1515) );
  XNOR2_X1 U1653 ( .A(n1516), .B(n1515), .ZN(n1520) );
  XOR2_X1 U1654 ( .A(G244), .B(G226), .Z(n1518) );
  XNOR2_X1 U1655 ( .A(G238), .B(G232), .ZN(n1517) );
  XNOR2_X1 U1656 ( .A(n1518), .B(n1517), .ZN(n2046) );
  NAND2_X1 U1657 ( .A1(G45), .A2(n2046), .ZN(n1519) );
  NAND2_X1 U1658 ( .A1(n1520), .A2(n1519), .ZN(n1521) );
  NAND2_X1 U1659 ( .A1(n1521), .A2(n1896), .ZN(n1524) );
  NAND2_X1 U1660 ( .A1(n1979), .A2(n1522), .ZN(n1523) );
  NAND2_X1 U1661 ( .A1(n1524), .A2(n1523), .ZN(n1526) );
  INV_X1 U1662 ( .A(n1821), .ZN(n1770) );
  NOR2_X1 U1663 ( .A1(n2009), .A2(n1770), .ZN(n1525) );
  NOR2_X1 U1664 ( .A1(n1526), .A2(n1525), .ZN(n1527) );
  NOR2_X1 U1665 ( .A1(n1899), .A2(n1527), .ZN(n1544) );
  NAND2_X1 U1666 ( .A1(G97), .A2(n1844), .ZN(n1905) );
  NAND2_X1 U1667 ( .A1(n1946), .A2(n1905), .ZN(n1541) );
  NOR2_X1 U1668 ( .A1(n2030), .A2(n1924), .ZN(n1794) );
  NAND2_X1 U1669 ( .A1(n1926), .A2(G159), .ZN(n1529) );
  NAND2_X1 U1670 ( .A1(n1934), .A2(G50), .ZN(n1528) );
  NAND2_X1 U1671 ( .A1(n1529), .A2(n1528), .ZN(n1530) );
  NOR2_X1 U1672 ( .A1(n1794), .A2(n1530), .ZN(n1539) );
  NAND2_X1 U1673 ( .A1(n1931), .A2(G68), .ZN(n1531) );
  NAND2_X1 U1674 ( .A1(G87), .A2(n1909), .ZN(n1692) );
  NAND2_X1 U1675 ( .A1(n1531), .A2(n1692), .ZN(n1532) );
  XNOR2_X1 U1676 ( .A(n1532), .B(KEYINPUT114), .ZN(n1537) );
  NAND2_X1 U1677 ( .A1(n1933), .A2(G150), .ZN(n1534) );
  NAND2_X1 U1678 ( .A1(n1927), .A2(G58), .ZN(n1533) );
  NAND2_X1 U1679 ( .A1(n1534), .A2(n1533), .ZN(n1535) );
  XOR2_X1 U1680 ( .A(KEYINPUT113), .B(n1535), .Z(n1536) );
  NOR2_X1 U1681 ( .A1(n1537), .A2(n1536), .ZN(n1538) );
  NAND2_X1 U1682 ( .A1(n1539), .A2(n1538), .ZN(n1540) );
  NOR2_X1 U1683 ( .A1(n1541), .A2(n1540), .ZN(n1542) );
  XOR2_X1 U1684 ( .A(KEYINPUT115), .B(n1542), .Z(n1543) );
  NOR2_X1 U1685 ( .A1(n1544), .A2(n1543), .ZN(n1545) );
  NAND2_X1 U1686 ( .A1(n1546), .A2(n1545), .ZN(n1549) );
  NOR2_X1 U1687 ( .A1(n1549), .A2(n1548), .ZN(n1555) );
  XNOR2_X1 U1688 ( .A(n1551), .B(n1873), .ZN(n1550) );
  NAND2_X1 U1689 ( .A1(n1550), .A2(n2014), .ZN(n1553) );
  INV_X1 U1690 ( .A(n1820), .ZN(n1872) );
  NAND2_X1 U1691 ( .A1(n1551), .A2(n1872), .ZN(n1552) );
  NAND2_X1 U1692 ( .A1(n1553), .A2(n1552), .ZN(n1554) );
  OR2_X1 U1693 ( .A1(n1555), .A2(n1554), .ZN(G393) );
  NAND2_X1 U1694 ( .A1(n1622), .A2(G159), .ZN(n1557) );
  INV_X1 U1695 ( .A(G58), .ZN(n1925) );
  NAND2_X1 U1696 ( .A1(n1623), .A2(n1925), .ZN(n1556) );
  NAND2_X1 U1697 ( .A1(n1557), .A2(n1556), .ZN(n1561) );
  NAND2_X1 U1698 ( .A1(G58), .A2(n1627), .ZN(n1559) );
  NAND2_X1 U1699 ( .A1(n1626), .A2(G68), .ZN(n1558) );
  NAND2_X1 U1700 ( .A1(n1559), .A2(n1558), .ZN(n1560) );
  NOR2_X1 U1701 ( .A1(n1561), .A2(n1560), .ZN(n1564) );
  NAND2_X1 U1702 ( .A1(n1633), .A2(n1562), .ZN(n1563) );
  NAND2_X1 U1703 ( .A1(n1564), .A2(n1563), .ZN(n1565) );
  XOR2_X1 U1704 ( .A(KEYINPUT30), .B(n1565), .Z(n1737) );
  XNOR2_X1 U1705 ( .A(KEYINPUT103), .B(n1737), .ZN(n1651) );
  XOR2_X1 U1706 ( .A(KEYINPUT104), .B(KEYINPUT31), .Z(n1567) );
  NAND2_X1 U1707 ( .A1(G87), .A2(n1307), .ZN(n1566) );
  XNOR2_X1 U1708 ( .A(n1567), .B(n1566), .ZN(n1569) );
  NAND2_X1 U1709 ( .A1(n1617), .A2(G232), .ZN(n1568) );
  NAND2_X1 U1710 ( .A1(n1569), .A2(n1568), .ZN(n1575) );
  NAND2_X1 U1711 ( .A1(n1611), .A2(G226), .ZN(n1570) );
  XNOR2_X1 U1712 ( .A(n1570), .B(KEYINPUT32), .ZN(n1572) );
  NAND2_X1 U1713 ( .A1(G223), .A2(n1614), .ZN(n1571) );
  NAND2_X1 U1714 ( .A1(n1572), .A2(n1571), .ZN(n1573) );
  XOR2_X1 U1715 ( .A(KEYINPUT33), .B(n1573), .Z(n1574) );
  NOR2_X1 U1716 ( .A1(n1575), .A2(n1574), .ZN(n1576) );
  NAND2_X1 U1717 ( .A1(n1576), .A2(n1613), .ZN(n1648) );
  INV_X1 U1718 ( .A(n1648), .ZN(n1578) );
  NOR2_X1 U1719 ( .A1(n1578), .A2(n1639), .ZN(n1577) );
  XNOR2_X1 U1720 ( .A(n1577), .B(KEYINPUT35), .ZN(n1580) );
  NAND2_X1 U1721 ( .A1(n1578), .A2(G190), .ZN(n1579) );
  NAND2_X1 U1722 ( .A1(n1580), .A2(n1579), .ZN(n1581) );
  NOR2_X1 U1723 ( .A1(n1651), .A2(n1581), .ZN(n1739) );
  XOR2_X1 U1724 ( .A(KEYINPUT101), .B(KEYINPUT28), .Z(n1590) );
  NAND2_X1 U1725 ( .A1(n1614), .A2(G226), .ZN(n1582) );
  NAND2_X1 U1726 ( .A1(n1613), .A2(n1582), .ZN(n1584) );
  AND2_X1 U1727 ( .A1(n1611), .A2(G232), .ZN(n1583) );
  NAND2_X1 U1728 ( .A1(G238), .A2(n1617), .ZN(n1585) );
  INV_X1 U1729 ( .A(n1606), .ZN(n1588) );
  NAND2_X1 U1730 ( .A1(G190), .A2(n1588), .ZN(n1589) );
  XNOR2_X1 U1731 ( .A(n1590), .B(n1589), .ZN(n1602) );
  NAND2_X1 U1732 ( .A1(n1627), .A2(G68), .ZN(n1591) );
  XNOR2_X1 U1733 ( .A(n1591), .B(KEYINPUT98), .ZN(n1598) );
  NAND2_X1 U1734 ( .A1(G77), .A2(n1626), .ZN(n1593) );
  NAND2_X1 U1735 ( .A1(G50), .A2(n1622), .ZN(n1592) );
  NAND2_X1 U1736 ( .A1(n1593), .A2(n1592), .ZN(n1596) );
  NOR2_X1 U1737 ( .A1(G68), .A2(n1594), .ZN(n1595) );
  NOR2_X1 U1738 ( .A1(n1596), .A2(n1595), .ZN(n1597) );
  NAND2_X1 U1739 ( .A1(n1598), .A2(n1597), .ZN(n1607) );
  NAND2_X1 U1740 ( .A1(G200), .A2(n1606), .ZN(n1599) );
  XNOR2_X1 U1741 ( .A(KEYINPUT27), .B(n1599), .ZN(n1600) );
  NOR2_X1 U1742 ( .A1(n1607), .A2(n1600), .ZN(n1601) );
  NAND2_X1 U1743 ( .A1(n1602), .A2(n1601), .ZN(n1603) );
  XNOR2_X1 U1744 ( .A(n1603), .B(KEYINPUT102), .ZN(n1610) );
  NOR2_X1 U1745 ( .A1(n1606), .A2(G179), .ZN(n1604) );
  XOR2_X1 U1746 ( .A(n1604), .B(KEYINPUT100), .Z(n1609) );
  NAND2_X1 U1747 ( .A1(n1606), .A2(n1605), .ZN(n1608) );
  INV_X1 U1748 ( .A(n1607), .ZN(n1673) );
  INV_X1 U1749 ( .A(n1659), .ZN(n1728) );
  INV_X1 U1750 ( .A(n1676), .ZN(n1655) );
  NAND2_X1 U1751 ( .A1(n1611), .A2(G223), .ZN(n1612) );
  NAND2_X1 U1752 ( .A1(n1613), .A2(n1612), .ZN(n1616) );
  NAND2_X1 U1753 ( .A1(n1614), .A2(G222), .ZN(n1615) );
  NOR2_X1 U1754 ( .A1(n1616), .A2(n1107), .ZN(n1619) );
  NAND2_X1 U1755 ( .A1(n1617), .A2(G226), .ZN(n1618) );
  NAND2_X1 U1756 ( .A1(n1619), .A2(n1618), .ZN(n1621) );
  NOR2_X1 U1757 ( .A1(n1587), .A2(n2030), .ZN(n1620) );
  NAND2_X1 U1758 ( .A1(n1640), .A2(n1126), .ZN(n1636) );
  NAND2_X1 U1759 ( .A1(n1622), .A2(G150), .ZN(n1625) );
  NAND2_X1 U1760 ( .A1(n1623), .A2(n1767), .ZN(n1624) );
  NAND2_X1 U1761 ( .A1(n1625), .A2(n1624), .ZN(n1631) );
  NAND2_X1 U1762 ( .A1(G58), .A2(n1626), .ZN(n1629) );
  NAND2_X1 U1763 ( .A1(n1627), .A2(G50), .ZN(n1628) );
  NAND2_X1 U1764 ( .A1(n1629), .A2(n1628), .ZN(n1630) );
  NOR2_X1 U1765 ( .A1(n1631), .A2(n1630), .ZN(n1635) );
  NAND2_X1 U1766 ( .A1(n1632), .A2(n1767), .ZN(n2042) );
  NAND2_X1 U1767 ( .A1(n1633), .A2(n2042), .ZN(n1634) );
  NAND2_X1 U1768 ( .A1(n1635), .A2(n1634), .ZN(n1758) );
  NAND2_X1 U1769 ( .A1(n1636), .A2(n1758), .ZN(n1638) );
  NOR2_X1 U1770 ( .A1(G169), .A2(n1640), .ZN(n1637) );
  NOR2_X1 U1771 ( .A1(n1638), .A2(n1637), .ZN(n1762) );
  OR2_X1 U1772 ( .A1(n1639), .A2(n1640), .ZN(n1642) );
  NAND2_X1 U1773 ( .A1(G190), .A2(n1640), .ZN(n1641) );
  NAND2_X1 U1774 ( .A1(n1642), .A2(n1641), .ZN(n1643) );
  NOR2_X1 U1775 ( .A1(n1758), .A2(n1643), .ZN(n1644) );
  NOR2_X1 U1776 ( .A1(n1762), .A2(n1644), .ZN(n1645) );
  XNOR2_X1 U1777 ( .A(KEYINPUT37), .B(n1645), .ZN(n1663) );
  INV_X1 U1778 ( .A(n1663), .ZN(n1759) );
  NOR2_X1 U1779 ( .A1(n1648), .A2(n1126), .ZN(n1647) );
  XNOR2_X1 U1780 ( .A(KEYINPUT34), .B(KEYINPUT105), .ZN(n1646) );
  XNOR2_X1 U1781 ( .A(n1647), .B(n1646), .ZN(n1650) );
  NAND2_X1 U1782 ( .A1(n1648), .A2(G169), .ZN(n1649) );
  NAND2_X1 U1783 ( .A1(n1650), .A2(n1649), .ZN(n1735) );
  NAND2_X1 U1784 ( .A1(n1651), .A2(n1735), .ZN(n1749) );
  NAND2_X1 U1785 ( .A1(n1759), .A2(n1749), .ZN(n1652) );
  NOR2_X1 U1786 ( .A1(n1653), .A2(n1652), .ZN(n1654) );
  NAND2_X1 U1787 ( .A1(n1655), .A2(n1654), .ZN(n1656) );
  NAND2_X1 U1788 ( .A1(n1681), .A2(n1657), .ZN(n1665) );
  INV_X1 U1789 ( .A(n1749), .ZN(n1740) );
  NOR2_X1 U1790 ( .A1(n1667), .A2(n1676), .ZN(n1658) );
  NOR2_X1 U1791 ( .A1(n1659), .A2(n1658), .ZN(n1660) );
  NOR2_X1 U1792 ( .A1(n1739), .A2(n1660), .ZN(n1661) );
  NOR2_X1 U1793 ( .A1(n1740), .A2(n1661), .ZN(n1662) );
  NOR2_X1 U1794 ( .A1(n1663), .A2(n1662), .ZN(n1664) );
  NOR2_X1 U1795 ( .A1(n1762), .A2(n1664), .ZN(n1682) );
  NAND2_X1 U1796 ( .A1(n1665), .A2(n1682), .ZN(G369) );
  NAND2_X1 U1797 ( .A1(n1668), .A2(n1667), .ZN(n1669) );
  INV_X1 U1798 ( .A(n1732), .ZN(n1672) );
  NOR2_X1 U1799 ( .A1(n1673), .A2(n1886), .ZN(n1674) );
  XOR2_X1 U1800 ( .A(KEYINPUT99), .B(n1674), .Z(n1675) );
  NOR2_X1 U1801 ( .A1(n1676), .A2(n1675), .ZN(n1678) );
  NOR2_X1 U1802 ( .A1(n1886), .A2(n1728), .ZN(n1677) );
  INV_X1 U1803 ( .A(n1752), .ZN(n1731) );
  XNOR2_X1 U1804 ( .A(n1680), .B(n1752), .ZN(n1816) );
  INV_X1 U1805 ( .A(n1816), .ZN(n1746) );
  INV_X1 U1806 ( .A(n1681), .ZN(n2006) );
  NAND2_X1 U1807 ( .A1(G330), .A2(n2020), .ZN(n1684) );
  NAND2_X1 U1808 ( .A1(n1881), .A2(n1682), .ZN(n1683) );
  NAND2_X1 U1809 ( .A1(G369), .A2(n1683), .ZN(n2025) );
  NAND2_X1 U1810 ( .A1(n1684), .A2(n2025), .ZN(n1685) );
  NAND2_X1 U1811 ( .A1(G107), .A2(n1931), .ZN(n1686) );
  NAND2_X1 U1812 ( .A1(G77), .A2(n1844), .ZN(n1937) );
  NAND2_X1 U1813 ( .A1(n1686), .A2(n1937), .ZN(n1698) );
  NOR2_X1 U1814 ( .A1(n1687), .A2(n1924), .ZN(n1688) );
  NOR2_X1 U1815 ( .A1(n1829), .A2(n1688), .ZN(n1696) );
  NAND2_X1 U1816 ( .A1(n1934), .A2(G283), .ZN(n1690) );
  NAND2_X1 U1817 ( .A1(n1927), .A2(G116), .ZN(n1689) );
  NAND2_X1 U1818 ( .A1(n1690), .A2(n1689), .ZN(n1694) );
  NAND2_X1 U1819 ( .A1(G303), .A2(n1933), .ZN(n1691) );
  NAND2_X1 U1820 ( .A1(n1692), .A2(n1691), .ZN(n1693) );
  NOR2_X1 U1821 ( .A1(n1694), .A2(n1693), .ZN(n1695) );
  NAND2_X1 U1822 ( .A1(n1696), .A2(n1695), .ZN(n1697) );
  NOR2_X1 U1823 ( .A1(n1698), .A2(n1697), .ZN(n1700) );
  NAND2_X1 U1824 ( .A1(G294), .A2(n1926), .ZN(n1699) );
  NAND2_X1 U1825 ( .A1(n1700), .A2(n1699), .ZN(n1703) );
  INV_X1 U1826 ( .A(G68), .ZN(n1701) );
  NAND2_X1 U1827 ( .A1(n1861), .A2(n1701), .ZN(n1702) );
  NAND2_X1 U1828 ( .A1(n1703), .A2(n1702), .ZN(n1720) );
  NAND2_X1 U1829 ( .A1(G143), .A2(n1927), .ZN(n1705) );
  NAND2_X1 U1830 ( .A1(G128), .A2(n1933), .ZN(n1704) );
  NAND2_X1 U1831 ( .A1(n1705), .A2(n1704), .ZN(n1718) );
  NAND2_X1 U1832 ( .A1(G150), .A2(n1931), .ZN(n1706) );
  NAND2_X1 U1833 ( .A1(n1946), .A2(n1706), .ZN(n1714) );
  NAND2_X1 U1834 ( .A1(G137), .A2(n1934), .ZN(n1708) );
  NAND2_X1 U1835 ( .A1(n1912), .A2(G159), .ZN(n1707) );
  NAND2_X1 U1836 ( .A1(n1708), .A2(n1707), .ZN(n1711) );
  NOR2_X1 U1837 ( .A1(n1709), .A2(n1767), .ZN(n1710) );
  NOR2_X1 U1838 ( .A1(n1711), .A2(n1710), .ZN(n1712) );
  NAND2_X1 U1839 ( .A1(G58), .A2(n1844), .ZN(n1800) );
  NAND2_X1 U1840 ( .A1(n1712), .A2(n1800), .ZN(n1713) );
  NOR2_X1 U1841 ( .A1(n1714), .A2(n1713), .ZN(n1716) );
  NAND2_X1 U1842 ( .A1(n1926), .A2(G132), .ZN(n1715) );
  NAND2_X1 U1843 ( .A1(n1716), .A2(n1715), .ZN(n1717) );
  NOR2_X1 U1844 ( .A1(n1718), .A2(n1717), .ZN(n1719) );
  NOR2_X1 U1845 ( .A1(n1720), .A2(n1719), .ZN(n1721) );
  NAND2_X1 U1846 ( .A1(n1902), .A2(n1721), .ZN(n1722) );
  XOR2_X1 U1847 ( .A(KEYINPUT45), .B(n1722), .Z(n1724) );
  NOR2_X1 U1848 ( .A1(n1731), .A2(n1770), .ZN(n1723) );
  NOR2_X1 U1849 ( .A1(n1724), .A2(n1723), .ZN(n1726) );
  NOR2_X1 U1850 ( .A1(n1820), .A2(n1746), .ZN(n1725) );
  NOR2_X1 U1851 ( .A1(n1726), .A2(n1725), .ZN(n1727) );
  NAND2_X1 U1852 ( .A1(n1732), .A2(n1731), .ZN(n1733) );
  XOR2_X1 U1853 ( .A(KEYINPUT39), .B(n1733), .Z(n1734) );
  NAND2_X1 U1854 ( .A1(n1748), .A2(n1734), .ZN(n1745) );
  NOR2_X1 U1855 ( .A1(n1735), .A2(n1761), .ZN(n1736) );
  NOR2_X1 U1856 ( .A1(n1737), .A2(n1736), .ZN(n1738) );
  NOR2_X1 U1857 ( .A1(n1739), .A2(n1738), .ZN(n1742) );
  AND2_X1 U1858 ( .A1(n1740), .A2(n1761), .ZN(n1741) );
  NOR2_X1 U1859 ( .A1(n1742), .A2(n1741), .ZN(n1822) );
  XOR2_X1 U1860 ( .A(KEYINPUT40), .B(n1822), .Z(n1743) );
  NOR2_X1 U1861 ( .A1(n1748), .A2(n1822), .ZN(n1751) );
  NOR2_X1 U1862 ( .A1(n1761), .A2(n1749), .ZN(n1750) );
  NOR2_X1 U1863 ( .A1(n1751), .A2(n1750), .ZN(n2018) );
  NOR2_X1 U1864 ( .A1(n1752), .A2(n1822), .ZN(n1753) );
  NAND2_X1 U1865 ( .A1(n1754), .A2(n1753), .ZN(n1755) );
  NOR2_X1 U1866 ( .A1(n1756), .A2(n1755), .ZN(n2019) );
  NAND2_X1 U1867 ( .A1(G330), .A2(n2019), .ZN(n1757) );
  NAND2_X1 U1868 ( .A1(n1758), .A2(n1761), .ZN(n1760) );
  NAND2_X1 U1869 ( .A1(n1760), .A2(n1759), .ZN(n1764) );
  NAND2_X1 U1870 ( .A1(n1762), .A2(n1761), .ZN(n1763) );
  NAND2_X1 U1871 ( .A1(n1764), .A2(n1763), .ZN(n1771) );
  NAND2_X1 U1872 ( .A1(n1766), .A2(n1765), .ZN(n1768) );
  NAND2_X1 U1873 ( .A1(n1768), .A2(n1767), .ZN(n1769) );
  NAND2_X1 U1874 ( .A1(n1770), .A2(n1769), .ZN(n1773) );
  NAND2_X1 U1875 ( .A1(n1821), .A2(n1771), .ZN(n1772) );
  NAND2_X1 U1876 ( .A1(n1773), .A2(n1772), .ZN(n1814) );
  NAND2_X1 U1877 ( .A1(n1844), .A2(G159), .ZN(n1775) );
  NAND2_X1 U1878 ( .A1(n1927), .A2(G132), .ZN(n1774) );
  NAND2_X1 U1879 ( .A1(n1775), .A2(n1774), .ZN(n1776) );
  XNOR2_X1 U1880 ( .A(n1776), .B(KEYINPUT44), .ZN(n1791) );
  NAND2_X1 U1881 ( .A1(G128), .A2(n1934), .ZN(n1777) );
  XOR2_X1 U1882 ( .A(KEYINPUT106), .B(n1777), .Z(n1781) );
  NAND2_X1 U1883 ( .A1(G150), .A2(n1909), .ZN(n1779) );
  NAND2_X1 U1884 ( .A1(n1912), .A2(G143), .ZN(n1778) );
  NAND2_X1 U1885 ( .A1(n1779), .A2(n1778), .ZN(n1780) );
  NOR2_X1 U1886 ( .A1(n1781), .A2(n1780), .ZN(n1789) );
  NAND2_X1 U1887 ( .A1(n1933), .A2(G124), .ZN(n1782) );
  NAND2_X1 U1888 ( .A1(n1946), .A2(n1782), .ZN(n1787) );
  NAND2_X1 U1889 ( .A1(n1926), .A2(G125), .ZN(n1785) );
  NAND2_X1 U1890 ( .A1(G137), .A2(n1931), .ZN(n1783) );
  XOR2_X1 U1891 ( .A(KEYINPUT43), .B(n1783), .Z(n1784) );
  NAND2_X1 U1892 ( .A1(n1785), .A2(n1784), .ZN(n1786) );
  NOR2_X1 U1893 ( .A1(n1787), .A2(n1786), .ZN(n1788) );
  NAND2_X1 U1894 ( .A1(n1789), .A2(n1788), .ZN(n1790) );
  NOR2_X1 U1895 ( .A1(n1791), .A2(n1790), .ZN(n1810) );
  NAND2_X1 U1896 ( .A1(n1926), .A2(G116), .ZN(n1796) );
  NAND2_X1 U1897 ( .A1(G283), .A2(n1933), .ZN(n1792) );
  XNOR2_X1 U1898 ( .A(KEYINPUT107), .B(n1792), .ZN(n1793) );
  NOR2_X1 U1899 ( .A1(n1794), .A2(n1793), .ZN(n1795) );
  NAND2_X1 U1900 ( .A1(n1796), .A2(n1795), .ZN(n1797) );
  XNOR2_X1 U1901 ( .A(n1797), .B(KEYINPUT108), .ZN(n1808) );
  NAND2_X1 U1902 ( .A1(G107), .A2(n1934), .ZN(n1798) );
  XOR2_X1 U1903 ( .A(KEYINPUT42), .B(n1798), .Z(n1799) );
  NOR2_X1 U1904 ( .A1(n1829), .A2(n1799), .ZN(n1806) );
  NAND2_X1 U1905 ( .A1(G68), .A2(n1909), .ZN(n1938) );
  NAND2_X1 U1906 ( .A1(n1938), .A2(n1800), .ZN(n1804) );
  NAND2_X1 U1907 ( .A1(n1931), .A2(G87), .ZN(n1802) );
  NAND2_X1 U1908 ( .A1(n1927), .A2(G97), .ZN(n1801) );
  NAND2_X1 U1909 ( .A1(n1802), .A2(n1801), .ZN(n1803) );
  NOR2_X1 U1910 ( .A1(n1804), .A2(n1803), .ZN(n1805) );
  NAND2_X1 U1911 ( .A1(n1806), .A2(n1805), .ZN(n1807) );
  NOR2_X1 U1912 ( .A1(n1808), .A2(n1807), .ZN(n1809) );
  NOR2_X1 U1913 ( .A1(n1810), .A2(n1809), .ZN(n1811) );
  NOR2_X1 U1914 ( .A1(G41), .A2(n1811), .ZN(n1812) );
  NOR2_X1 U1915 ( .A1(n1812), .A2(n1876), .ZN(n1813) );
  NAND2_X1 U1916 ( .A1(n1814), .A2(n1813), .ZN(n1815) );
  NOR2_X1 U1917 ( .A1(n1820), .A2(n1819), .ZN(n1869) );
  NAND2_X1 U1918 ( .A1(n1822), .A2(n1821), .ZN(n1868) );
  NAND2_X1 U1919 ( .A1(G107), .A2(n1927), .ZN(n1824) );
  NAND2_X1 U1920 ( .A1(n1824), .A2(n1823), .ZN(n1833) );
  NOR2_X1 U1921 ( .A1(n1826), .A2(n1825), .ZN(n1831) );
  NAND2_X1 U1922 ( .A1(n1934), .A2(G116), .ZN(n1827) );
  XNOR2_X1 U1923 ( .A(KEYINPUT47), .B(n1827), .ZN(n1828) );
  NOR2_X1 U1924 ( .A1(n1829), .A2(n1828), .ZN(n1830) );
  NAND2_X1 U1925 ( .A1(n1831), .A2(n1830), .ZN(n1832) );
  NOR2_X1 U1926 ( .A1(n1833), .A2(n1832), .ZN(n1835) );
  NAND2_X1 U1927 ( .A1(G283), .A2(n1926), .ZN(n1834) );
  NAND2_X1 U1928 ( .A1(n1835), .A2(n1834), .ZN(n1836) );
  XNOR2_X1 U1929 ( .A(KEYINPUT110), .B(n1836), .ZN(n1843) );
  NAND2_X1 U1930 ( .A1(G294), .A2(n1933), .ZN(n1837) );
  XNOR2_X1 U1931 ( .A(KEYINPUT111), .B(n1837), .ZN(n1840) );
  NAND2_X1 U1932 ( .A1(G97), .A2(n1931), .ZN(n1838) );
  XOR2_X1 U1933 ( .A(KEYINPUT112), .B(n1838), .Z(n1839) );
  NOR2_X1 U1934 ( .A1(n1840), .A2(n1839), .ZN(n1841) );
  XOR2_X1 U1935 ( .A(KEYINPUT48), .B(n1841), .Z(n1842) );
  NOR2_X1 U1936 ( .A1(n1843), .A2(n1842), .ZN(n1866) );
  NAND2_X1 U1937 ( .A1(G143), .A2(n1931), .ZN(n1846) );
  NAND2_X1 U1938 ( .A1(n1844), .A2(G50), .ZN(n1845) );
  NAND2_X1 U1939 ( .A1(n1846), .A2(n1845), .ZN(n1859) );
  NAND2_X1 U1940 ( .A1(G159), .A2(n1909), .ZN(n1847) );
  NAND2_X1 U1941 ( .A1(n1946), .A2(n1847), .ZN(n1855) );
  NAND2_X1 U1942 ( .A1(G132), .A2(n1934), .ZN(n1849) );
  NAND2_X1 U1943 ( .A1(G137), .A2(n1927), .ZN(n1848) );
  NAND2_X1 U1944 ( .A1(n1849), .A2(n1848), .ZN(n1851) );
  AND2_X1 U1945 ( .A1(G150), .A2(n1912), .ZN(n1850) );
  NOR2_X1 U1946 ( .A1(n1851), .A2(n1850), .ZN(n1853) );
  NAND2_X1 U1947 ( .A1(n1933), .A2(G125), .ZN(n1852) );
  NAND2_X1 U1948 ( .A1(n1853), .A2(n1852), .ZN(n1854) );
  NOR2_X1 U1949 ( .A1(n1855), .A2(n1854), .ZN(n1857) );
  NAND2_X1 U1950 ( .A1(n1926), .A2(G128), .ZN(n1856) );
  NAND2_X1 U1951 ( .A1(n1857), .A2(n1856), .ZN(n1858) );
  NOR2_X1 U1952 ( .A1(n1859), .A2(n1858), .ZN(n1860) );
  NOR2_X1 U1953 ( .A1(n1876), .A2(n1860), .ZN(n1863) );
  NAND2_X1 U1954 ( .A1(n1861), .A2(n1925), .ZN(n1862) );
  NAND2_X1 U1955 ( .A1(n1863), .A2(n1862), .ZN(n1864) );
  XOR2_X1 U1956 ( .A(KEYINPUT109), .B(n1864), .Z(n1865) );
  NOR2_X1 U1957 ( .A1(n1866), .A2(n1865), .ZN(n1867) );
  NOR2_X1 U1958 ( .A1(n1873), .A2(n1872), .ZN(n1874) );
  NAND2_X1 U1959 ( .A1(n1875), .A2(n1874), .ZN(n1877) );
  NAND2_X1 U1960 ( .A1(n1879), .A2(n1886), .ZN(n1883) );
  NAND2_X1 U1961 ( .A1(n1881), .A2(n1880), .ZN(n1882) );
  NAND2_X1 U1962 ( .A1(n1883), .A2(n1882), .ZN(n1884) );
  XNOR2_X1 U1963 ( .A(n1884), .B(KEYINPUT53), .ZN(n1890) );
  NOR2_X1 U1964 ( .A1(n1886), .A2(n1885), .ZN(n1887) );
  NAND2_X1 U1965 ( .A1(n1888), .A2(n1887), .ZN(n1889) );
  NAND2_X1 U1966 ( .A1(n1890), .A2(n1889), .ZN(n1893) );
  NOR2_X1 U1967 ( .A1(n1891), .A2(n2007), .ZN(n1892) );
  NAND2_X1 U1968 ( .A1(n1979), .A2(G87), .ZN(n1901) );
  XNOR2_X1 U1969 ( .A(G264), .B(G257), .ZN(n1894) );
  XNOR2_X1 U1970 ( .A(n1894), .B(G270), .ZN(n1895) );
  XNOR2_X1 U1971 ( .A(G250), .B(n1895), .ZN(n2045) );
  NAND2_X1 U1972 ( .A1(n1896), .A2(n2045), .ZN(n1897) );
  XOR2_X1 U1973 ( .A(KEYINPUT118), .B(n1897), .Z(n1898) );
  NOR2_X1 U1974 ( .A1(n1899), .A2(n1898), .ZN(n1900) );
  NAND2_X1 U1975 ( .A1(n1901), .A2(n1900), .ZN(n1903) );
  NAND2_X1 U1976 ( .A1(n1903), .A2(n1902), .ZN(n1956) );
  NAND2_X1 U1977 ( .A1(G283), .A2(n1931), .ZN(n1904) );
  NAND2_X1 U1978 ( .A1(n1905), .A2(n1904), .ZN(n1923) );
  NAND2_X1 U1979 ( .A1(G317), .A2(n1933), .ZN(n1907) );
  NAND2_X1 U1980 ( .A1(n1934), .A2(G303), .ZN(n1906) );
  NAND2_X1 U1981 ( .A1(n1907), .A2(n1906), .ZN(n1920) );
  NAND2_X1 U1982 ( .A1(G311), .A2(n1926), .ZN(n1908) );
  XNOR2_X1 U1983 ( .A(n1908), .B(KEYINPUT54), .ZN(n1918) );
  NAND2_X1 U1984 ( .A1(G294), .A2(n1927), .ZN(n1911) );
  NAND2_X1 U1985 ( .A1(G107), .A2(n1909), .ZN(n1910) );
  NAND2_X1 U1986 ( .A1(n1911), .A2(n1910), .ZN(n1916) );
  NAND2_X1 U1987 ( .A1(G116), .A2(n1912), .ZN(n1913) );
  NAND2_X1 U1988 ( .A1(n1914), .A2(n1913), .ZN(n1915) );
  NOR2_X1 U1989 ( .A1(n1916), .A2(n1915), .ZN(n1917) );
  NAND2_X1 U1990 ( .A1(n1918), .A2(n1917), .ZN(n1919) );
  NOR2_X1 U1991 ( .A1(n1920), .A2(n1919), .ZN(n1921) );
  XNOR2_X1 U1992 ( .A(n1921), .B(KEYINPUT121), .ZN(n1922) );
  NOR2_X1 U1993 ( .A1(n1923), .A2(n1922), .ZN(n1950) );
  NOR2_X1 U1994 ( .A1(n1925), .A2(n1924), .ZN(n1948) );
  NAND2_X1 U1995 ( .A1(n1926), .A2(G143), .ZN(n1930) );
  NAND2_X1 U1996 ( .A1(n1927), .A2(G159), .ZN(n1928) );
  XOR2_X1 U1997 ( .A(KEYINPUT119), .B(n1928), .Z(n1929) );
  NAND2_X1 U1998 ( .A1(n1930), .A2(n1929), .ZN(n1944) );
  NAND2_X1 U1999 ( .A1(n1931), .A2(G50), .ZN(n1932) );
  XNOR2_X1 U2000 ( .A(n1932), .B(KEYINPUT120), .ZN(n1942) );
  NAND2_X1 U2001 ( .A1(G137), .A2(n1933), .ZN(n1936) );
  NAND2_X1 U2002 ( .A1(n1934), .A2(G150), .ZN(n1935) );
  NAND2_X1 U2003 ( .A1(n1936), .A2(n1935), .ZN(n1940) );
  NAND2_X1 U2004 ( .A1(n1938), .A2(n1937), .ZN(n1939) );
  NOR2_X1 U2005 ( .A1(n1940), .A2(n1939), .ZN(n1941) );
  NAND2_X1 U2006 ( .A1(n1942), .A2(n1941), .ZN(n1943) );
  NOR2_X1 U2007 ( .A1(n1944), .A2(n1943), .ZN(n1945) );
  NAND2_X1 U2008 ( .A1(n1946), .A2(n1945), .ZN(n1947) );
  NOR2_X1 U2009 ( .A1(n1948), .A2(n1947), .ZN(n1949) );
  NOR2_X1 U2010 ( .A1(n1950), .A2(n1949), .ZN(n1954) );
  NAND2_X1 U2011 ( .A1(n1952), .A2(n1951), .ZN(n1953) );
  NAND2_X1 U2012 ( .A1(n1954), .A2(n1953), .ZN(n1955) );
  XOR2_X1 U2013 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n1957) );
  XNOR2_X1 U2014 ( .A(G375), .B(G378), .ZN(n1961) );
  XNOR2_X1 U2015 ( .A(n1966), .B(n1961), .ZN(G402) );
  NOR2_X1 U2016 ( .A1(G343), .A2(n1976), .ZN(n1962) );
  NOR2_X1 U2017 ( .A1(n1961), .A2(n1962), .ZN(n1965) );
  NAND2_X1 U2018 ( .A1(n1962), .A2(G2897), .ZN(n1963) );
  NOR2_X2 U2019 ( .A1(n1965), .A2(n1964), .ZN(n1967) );
  XNOR2_X1 U2020 ( .A(n1967), .B(n1966), .ZN(G405) );
  NOR2_X1 U2021 ( .A1(G393), .A2(G381), .ZN(n1973) );
  OR2_X1 U2022 ( .A1(G375), .A2(G378), .ZN(n1974) );
  NOR2_X1 U2023 ( .A1(G384), .A2(G390), .ZN(n1970) );
  NOR2_X1 U2024 ( .A1(G396), .A2(G387), .ZN(n1969) );
  NAND2_X1 U2025 ( .A1(n1970), .A2(n1969), .ZN(n1971) );
  NOR2_X1 U2026 ( .A1(n1974), .A2(n1971), .ZN(n1972) );
  NAND2_X1 U2027 ( .A1(n1973), .A2(n1972), .ZN(G407) );
  NOR2_X1 U2028 ( .A1(G343), .A2(n1974), .ZN(n1975) );
  NOR2_X1 U2029 ( .A1(n1976), .A2(n1975), .ZN(n1977) );
  NAND2_X1 U2030 ( .A1(n1977), .A2(G407), .ZN(G409) );
  NAND2_X1 U2031 ( .A1(G20), .A2(n1121), .ZN(n2037) );
  INV_X1 U2032 ( .A(n2037), .ZN(n1978) );
  NAND2_X1 U2033 ( .A1(n2013), .A2(n1978), .ZN(n1983) );
  NOR2_X1 U2034 ( .A1(G264), .A2(G257), .ZN(n1980) );
  NOR2_X1 U2035 ( .A1(n1980), .A2(n1979), .ZN(n1981) );
  NAND2_X1 U2036 ( .A1(G250), .A2(n1981), .ZN(n1982) );
  NAND2_X1 U2037 ( .A1(n1983), .A2(n1982), .ZN(n2004) );
  NAND2_X1 U2038 ( .A1(G257), .A2(G97), .ZN(n1984) );
  XNOR2_X1 U2039 ( .A(n1984), .B(KEYINPUT126), .ZN(n1991) );
  NAND2_X1 U2040 ( .A1(G270), .A2(G116), .ZN(n1986) );
  NAND2_X1 U2041 ( .A1(G250), .A2(G87), .ZN(n1985) );
  NAND2_X1 U2042 ( .A1(n1986), .A2(n1985), .ZN(n1989) );
  NAND2_X1 U2043 ( .A1(G107), .A2(G264), .ZN(n1987) );
  XOR2_X1 U2044 ( .A(KEYINPUT50), .B(n1987), .Z(n1988) );
  NOR2_X1 U2045 ( .A1(n1989), .A2(n1988), .ZN(n1990) );
  NAND2_X1 U2046 ( .A1(n1991), .A2(n1990), .ZN(n2000) );
  NAND2_X1 U2047 ( .A1(G58), .A2(G232), .ZN(n1993) );
  NAND2_X1 U2048 ( .A1(G68), .A2(G238), .ZN(n1992) );
  NAND2_X1 U2049 ( .A1(n1993), .A2(n1992), .ZN(n1997) );
  NAND2_X1 U2050 ( .A1(G244), .A2(G77), .ZN(n1995) );
  NAND2_X1 U2051 ( .A1(G50), .A2(G226), .ZN(n1994) );
  NAND2_X1 U2052 ( .A1(n1995), .A2(n1994), .ZN(n1996) );
  NOR2_X1 U2053 ( .A1(n1997), .A2(n1996), .ZN(n1998) );
  XNOR2_X1 U2054 ( .A(KEYINPUT49), .B(n1998), .ZN(n1999) );
  NOR2_X1 U2055 ( .A1(n2000), .A2(n1999), .ZN(n2001) );
  NOR2_X1 U2056 ( .A1(n2002), .A2(n2001), .ZN(n2003) );
  NOR2_X1 U2057 ( .A1(n2004), .A2(n2003), .ZN(G361) );
  NOR2_X1 U2058 ( .A1(n2006), .A2(n2005), .ZN(G372) );
  NAND2_X1 U2059 ( .A1(n1073), .A2(n2007), .ZN(G399) );
  NOR2_X1 U2060 ( .A1(G1), .A2(n2008), .ZN(n2012) );
  NAND2_X1 U2061 ( .A1(G1), .A2(n2009), .ZN(n2010) );
  NOR2_X1 U2062 ( .A1(n2014), .A2(n2010), .ZN(n2011) );
  NOR2_X1 U2063 ( .A1(n2012), .A2(n2011), .ZN(n2016) );
  NAND2_X1 U2064 ( .A1(n2014), .A2(n2013), .ZN(n2015) );
  NAND2_X1 U2065 ( .A1(n2016), .A2(n2015), .ZN(G364) );
  NOR2_X1 U2066 ( .A1(G13), .A2(n2017), .ZN(n2034) );
  INV_X1 U2067 ( .A(n2034), .ZN(n2028) );
  XOR2_X1 U2068 ( .A(KEYINPUT127), .B(n2018), .Z(n2023) );
  XOR2_X1 U2069 ( .A(n2020), .B(n2019), .Z(n2021) );
  NAND2_X1 U2070 ( .A1(n2021), .A2(G330), .ZN(n2022) );
  XNOR2_X1 U2071 ( .A(n2023), .B(n2022), .ZN(n2024) );
  XOR2_X1 U2072 ( .A(n2025), .B(n2024), .Z(n2026) );
  NAND2_X1 U2073 ( .A1(n2026), .A2(n2037), .ZN(n2027) );
  NAND2_X1 U2074 ( .A1(n2028), .A2(n2027), .ZN(n2036) );
  NAND2_X1 U2075 ( .A1(G58), .A2(G50), .ZN(n2029) );
  XNOR2_X1 U2076 ( .A(n2029), .B(G68), .ZN(n2032) );
  NAND2_X1 U2077 ( .A1(n2030), .A2(G50), .ZN(n2031) );
  NAND2_X1 U2078 ( .A1(n2032), .A2(n2031), .ZN(n2033) );
  NAND2_X1 U2079 ( .A1(n2034), .A2(n2033), .ZN(n2035) );
  NAND2_X1 U2080 ( .A1(n2036), .A2(n2035), .ZN(n2041) );
  NOR2_X1 U2081 ( .A1(n1016), .A2(n2037), .ZN(n2039) );
  NAND2_X1 U2082 ( .A1(n2039), .A2(n2038), .ZN(n2040) );
  NAND2_X1 U2083 ( .A1(n2041), .A2(n2040), .ZN(G367) );
  NOR2_X1 U2084 ( .A1(G77), .A2(n2042), .ZN(G353) );
  XNOR2_X1 U2085 ( .A(n2044), .B(n2043), .ZN(G351) );
  XOR2_X1 U2086 ( .A(n2046), .B(n2045), .Z(G358) );
endmodule

