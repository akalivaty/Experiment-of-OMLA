//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1190, new_n1191, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XNOR2_X1  g0006(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G50), .B2(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G116), .ZN(new_n221));
  INV_X1    g0021(.A(G270), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n204), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(G58), .A2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n208), .B(new_n228), .C1(new_n231), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n222), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n254), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n257), .B1(new_n260), .B2(new_n225), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n261), .B(KEYINPUT71), .Z(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT68), .B(G1698), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n265), .B1(new_n210), .B2(new_n266), .C1(new_n267), .C2(new_n216), .ZN(new_n268));
  INV_X1    g0068(.A(new_n259), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n268), .B(new_n269), .C1(G107), .C2(new_n265), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G169), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n275), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT15), .B(G87), .Z(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n230), .A2(G33), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n229), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n253), .A2(G13), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n230), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n281), .A2(new_n283), .B1(new_n224), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(new_n253), .B2(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G77), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G179), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n262), .A2(new_n290), .A3(new_n270), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n273), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n209), .A2(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n276), .ZN(new_n295));
  INV_X1    g0095(.A(G50), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n294), .B1(new_n280), .B2(new_n224), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n283), .ZN(new_n298));
  XOR2_X1   g0098(.A(new_n298), .B(KEYINPUT11), .Z(new_n299));
  NOR2_X1   g0099(.A1(new_n284), .A2(new_n294), .ZN(new_n300));
  XOR2_X1   g0100(.A(new_n300), .B(KEYINPUT12), .Z(new_n301));
  INV_X1    g0101(.A(new_n287), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n209), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G226), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n267), .A2(new_n305), .B1(new_n216), .B2(new_n266), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n265), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G97), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n256), .B1(new_n309), .B2(new_n269), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT13), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n259), .A2(G238), .A3(new_n254), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n306), .A2(new_n265), .B1(G33), .B2(G97), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n312), .B(new_n257), .C1(new_n314), .C2(new_n259), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n304), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n313), .B2(new_n316), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n317), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT14), .B1(new_n323), .B2(new_n272), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(G179), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT14), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n317), .A2(new_n326), .A3(G169), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n304), .ZN(new_n329));
  AOI211_X1 g0129(.A(new_n293), .B(new_n322), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n260), .A2(new_n305), .ZN(new_n331));
  OR3_X1    g0131(.A1(new_n331), .A2(KEYINPUT67), .A3(new_n256), .ZN(new_n332));
  INV_X1    g0132(.A(G223), .ZN(new_n333));
  INV_X1    g0133(.A(G222), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n265), .B1(new_n333), .B2(new_n266), .C1(new_n267), .C2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(new_n269), .C1(G77), .C2(new_n265), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT67), .B1(new_n331), .B2(new_n256), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n272), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n230), .B1(new_n232), .B2(new_n296), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT69), .ZN(new_n341));
  INV_X1    g0141(.A(G150), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n274), .A2(new_n280), .B1(new_n342), .B2(new_n295), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n283), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n287), .A2(G50), .ZN(new_n345));
  INV_X1    g0145(.A(G13), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(G1), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G20), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n344), .B(new_n345), .C1(G50), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n339), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT70), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(G179), .B2(new_n338), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT9), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n338), .A2(new_n318), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n349), .A2(new_n353), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n338), .A2(G200), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n354), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT10), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n356), .A2(new_n357), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT10), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n360), .A2(new_n361), .A3(new_n354), .A4(new_n355), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n271), .A2(G200), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n262), .A2(G190), .A3(new_n270), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n364), .A2(new_n288), .A3(new_n286), .A4(new_n365), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n352), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n263), .A2(new_n230), .A3(new_n264), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT7), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n230), .A4(new_n264), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n209), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n215), .A2(new_n209), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n374), .B2(new_n232), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n276), .A2(G159), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n368), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g0178(.A1(KEYINPUT3), .A2(G33), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n381), .B2(new_n230), .ZN(new_n382));
  NOR4_X1   g0182(.A1(new_n379), .A2(new_n380), .A3(new_n370), .A4(G20), .ZN(new_n383));
  OAI21_X1  g0183(.A(G68), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n377), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n378), .A2(new_n386), .A3(new_n283), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n275), .A2(new_n348), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n287), .B2(new_n275), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n259), .A2(G232), .A3(new_n254), .ZN(new_n391));
  INV_X1    g0191(.A(G33), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n219), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G226), .A2(G1698), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n267), .B2(new_n333), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n395), .B2(new_n265), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n257), .B(new_n391), .C1(new_n396), .C2(new_n259), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n272), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT68), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G1698), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G223), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n381), .B1(new_n403), .B2(new_n394), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n269), .B1(new_n404), .B2(new_n393), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n405), .A2(new_n290), .A3(new_n257), .A4(new_n391), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n390), .A2(new_n398), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n407), .B(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n397), .A2(G200), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n405), .A2(G190), .A3(new_n257), .A4(new_n391), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n410), .A2(new_n387), .A3(new_n411), .A4(new_n389), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT17), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT72), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n409), .A2(new_n413), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT72), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n330), .B(new_n367), .C1(new_n414), .C2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n220), .B1(new_n263), .B2(new_n264), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n402), .ZN(new_n420));
  OAI211_X1 g0220(.A(G257), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT82), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n265), .A2(KEYINPUT82), .A3(G257), .A4(G1698), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G294), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n420), .A2(new_n423), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n269), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT5), .B(G41), .ZN(new_n428));
  INV_X1    g0228(.A(G45), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(G1), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G274), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n269), .B1(new_n430), .B2(new_n428), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G264), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n427), .A2(new_n318), .A3(new_n432), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT83), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n427), .A2(new_n432), .A3(new_n434), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n320), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n426), .A2(new_n269), .B1(G264), .B2(new_n433), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT83), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(new_n318), .A4(new_n432), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n436), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n211), .A2(G20), .ZN(new_n443));
  XOR2_X1   g0243(.A(new_n443), .B(KEYINPUT23), .Z(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G116), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n230), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n230), .B(G87), .C1(new_n379), .C2(new_n380), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n448), .A2(KEYINPUT22), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(KEYINPUT22), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n444), .B(new_n447), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT24), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n448), .B(KEYINPUT22), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n454), .A2(KEYINPUT24), .A3(new_n444), .A4(new_n447), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n455), .A3(new_n283), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n282), .A2(new_n229), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(new_n348), .C1(G1), .C2(new_n392), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G107), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n284), .A2(new_n443), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT25), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n456), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n442), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n419), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  OAI21_X1  g0266(.A(G244), .B1(new_n379), .B2(new_n380), .ZN(new_n467));
  OAI211_X1 g0267(.A(KEYINPUT75), .B(new_n466), .C1(new_n467), .C2(new_n267), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(KEYINPUT75), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n265), .A2(new_n402), .A3(G244), .A4(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n466), .A2(KEYINPUT75), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n465), .A2(new_n468), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(new_n269), .B1(G257), .B2(new_n433), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n432), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G200), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n348), .A2(G97), .ZN(new_n476));
  OAI21_X1  g0276(.A(G107), .B1(new_n382), .B2(new_n383), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT74), .ZN(new_n478));
  OR2_X1    g0278(.A1(KEYINPUT73), .A2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(KEYINPUT73), .A2(G97), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n479), .A2(KEYINPUT6), .A3(new_n211), .A4(new_n480), .ZN(new_n481));
  XOR2_X1   g0281(.A(G97), .B(G107), .Z(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(KEYINPUT6), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n483), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT74), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(G107), .C1(new_n382), .C2(new_n383), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n478), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n476), .B1(new_n487), .B2(new_n283), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n459), .A2(G97), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n473), .A2(G190), .A3(new_n432), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n475), .A2(new_n488), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n283), .ZN(new_n492));
  INV_X1    g0292(.A(new_n476), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n493), .A3(new_n489), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n474), .A2(new_n272), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n473), .A2(new_n290), .A3(new_n432), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n456), .A2(new_n460), .A3(new_n462), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n437), .A2(new_n272), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n439), .A2(new_n290), .A3(new_n432), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n464), .A2(new_n491), .A3(new_n497), .A4(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n230), .A2(G116), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT79), .B1(new_n457), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(G20), .B1(G33), .B2(G283), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n479), .A2(new_n480), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(G33), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT79), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n283), .B(new_n508), .C1(new_n230), .C2(G116), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT80), .B(KEYINPUT20), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n459), .A2(G116), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT80), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(KEYINPUT20), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n504), .A2(new_n507), .A3(new_n515), .A4(new_n509), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n347), .A2(new_n503), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n512), .A2(new_n513), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n433), .A2(G270), .B1(new_n431), .B2(G274), .ZN(new_n519));
  INV_X1    g0319(.A(G257), .ZN(new_n520));
  OAI221_X1 g0320(.A(new_n265), .B1(new_n212), .B2(new_n266), .C1(new_n267), .C2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G303), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n381), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n269), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n518), .A2(G169), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT21), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n518), .A2(new_n525), .A3(new_n528), .A4(G169), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n519), .A2(new_n524), .A3(G179), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n518), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT81), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT81), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n518), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n527), .A2(new_n529), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n480), .ZN(new_n536));
  NOR2_X1   g0336(.A1(KEYINPUT73), .A2(G97), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n219), .B(new_n211), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n230), .B1(new_n308), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n230), .B(G68), .C1(new_n379), .C2(new_n380), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT77), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n539), .B1(new_n506), .B2(new_n280), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n265), .A2(KEYINPUT77), .A3(new_n230), .A4(G68), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n541), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n283), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n279), .A2(new_n285), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n459), .A2(G87), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n210), .B1(new_n399), .B2(new_n401), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n225), .A2(new_n266), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n265), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n259), .B1(new_n554), .B2(new_n445), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n430), .A2(new_n255), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n220), .B1(new_n429), .B2(G1), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n259), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT76), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT76), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n267), .A2(new_n210), .B1(new_n225), .B2(new_n266), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n446), .B1(new_n562), .B2(new_n265), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n561), .B(new_n558), .C1(new_n563), .C2(new_n259), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n551), .B1(new_n565), .B2(G190), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n560), .A2(G200), .A3(new_n564), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n290), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n459), .A2(new_n278), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n548), .A2(new_n570), .A3(KEYINPUT78), .A4(new_n549), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n548), .A2(new_n549), .A3(new_n570), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT78), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n560), .A2(new_n272), .A3(new_n564), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n569), .A2(new_n571), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n525), .A2(new_n318), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n320), .B1(new_n519), .B2(new_n524), .ZN(new_n578));
  OR3_X1    g0378(.A1(new_n577), .A2(new_n518), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n535), .A2(new_n568), .A3(new_n576), .A4(new_n579), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n418), .A2(new_n502), .A3(new_n580), .ZN(G372));
  XNOR2_X1  g0381(.A(new_n407), .B(KEYINPUT18), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n328), .A2(new_n329), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n322), .B1(new_n583), .B2(new_n292), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n582), .B1(new_n584), .B2(new_n413), .ZN(new_n585));
  INV_X1    g0385(.A(new_n363), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n352), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n572), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n290), .B2(new_n565), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n555), .A2(new_n591), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n563), .A2(KEYINPUT84), .A3(new_n259), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n558), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n272), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(G200), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n590), .A2(new_n595), .B1(new_n566), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n597), .A2(new_n464), .A3(new_n497), .A4(new_n491), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n527), .A2(new_n529), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n532), .A2(new_n534), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT85), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT85), .B1(new_n600), .B2(new_n601), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n501), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n568), .A2(new_n576), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT26), .B1(new_n606), .B2(new_n497), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT26), .ZN(new_n608));
  INV_X1    g0408(.A(new_n497), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n597), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n590), .A2(new_n595), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n588), .B1(new_n418), .B2(new_n614), .ZN(G369));
  NAND2_X1  g0415(.A1(new_n600), .A2(new_n601), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n535), .A2(KEYINPUT85), .ZN(new_n619));
  OR3_X1    g0419(.A1(new_n284), .A2(KEYINPUT27), .A3(G20), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT27), .B1(new_n284), .B2(G20), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(G213), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(G343), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n618), .A2(new_n619), .A3(new_n518), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n518), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n535), .A2(new_n579), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g0428(.A(new_n628), .B(KEYINPUT86), .Z(new_n629));
  AND2_X1   g0429(.A1(new_n629), .A2(G330), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n501), .A2(new_n624), .ZN(new_n631));
  INV_X1    g0431(.A(new_n624), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n464), .B1(new_n463), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n631), .B1(new_n633), .B2(new_n501), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n535), .A2(new_n624), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(new_n631), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(G399));
  INV_X1    g0439(.A(new_n205), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G41), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n538), .A2(G116), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n641), .A2(new_n642), .A3(new_n253), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n235), .B2(new_n641), .ZN(new_n644));
  XOR2_X1   g0444(.A(new_n644), .B(KEYINPUT28), .Z(new_n645));
  NAND4_X1  g0445(.A1(new_n609), .A2(new_n608), .A3(new_n568), .A4(new_n576), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n600), .A2(new_n501), .A3(new_n601), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n566), .A2(new_n596), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n464), .A2(new_n491), .A3(new_n497), .A4(new_n648), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n646), .B(new_n611), .C1(new_n647), .C2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n608), .B1(new_n597), .B2(new_n609), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n632), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT29), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n613), .A2(new_n632), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(KEYINPUT29), .ZN(new_n655));
  INV_X1    g0455(.A(G330), .ZN(new_n656));
  INV_X1    g0456(.A(new_n473), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n427), .A2(new_n434), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n564), .B2(new_n560), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n657), .B1(new_n659), .B2(KEYINPUT87), .ZN(new_n660));
  INV_X1    g0460(.A(new_n530), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n565), .A2(new_n439), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT87), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT30), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n594), .A2(new_n290), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n668), .A2(new_n437), .A3(new_n474), .A4(new_n525), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n667), .A2(KEYINPUT88), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n660), .A2(new_n664), .A3(KEYINPUT30), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT88), .B1(new_n667), .B2(new_n669), .ZN(new_n673));
  OAI211_X1 g0473(.A(KEYINPUT31), .B(new_n624), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n667), .A2(new_n671), .A3(new_n669), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n624), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n580), .A2(new_n502), .A3(new_n624), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT31), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n656), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n655), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n645), .B1(new_n681), .B2(G1), .ZN(G364));
  NOR2_X1   g0482(.A1(new_n346), .A2(G20), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n253), .B1(new_n683), .B2(G45), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n641), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n630), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(G330), .B2(new_n629), .ZN(new_n688));
  NOR2_X1   g0488(.A1(G13), .A2(G33), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G20), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n625), .A2(new_n627), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n229), .B1(G20), .B2(new_n272), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n290), .A2(new_n320), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n230), .A2(G190), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n230), .A2(new_n318), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n320), .A2(G179), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n209), .A2(new_n696), .B1(new_n699), .B2(new_n219), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G179), .A2(G200), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n230), .B1(new_n701), .B2(G190), .ZN(new_n702));
  INV_X1    g0502(.A(G97), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n695), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n705), .B1(new_n211), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT32), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n695), .A2(new_n701), .ZN(new_n709));
  INV_X1    g0509(.A(G159), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n709), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(KEYINPUT32), .A3(G159), .ZN(new_n713));
  AOI211_X1 g0513(.A(new_n381), .B(new_n707), .C1(new_n711), .C2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n697), .A2(new_n694), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n290), .A2(G200), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n695), .ZN(new_n717));
  OAI221_X1 g0517(.A(new_n714), .B1(new_n296), .B2(new_n715), .C1(new_n224), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n697), .A2(new_n716), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n718), .B1(G58), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G326), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n715), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n699), .B(KEYINPUT89), .Z(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G303), .ZN(new_n726));
  INV_X1    g0526(.A(G311), .ZN(new_n727));
  INV_X1    g0527(.A(G329), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n717), .A2(new_n727), .B1(new_n709), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n706), .ZN(new_n730));
  AOI211_X1 g0530(.A(new_n265), .B(new_n729), .C1(G283), .C2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n702), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G294), .ZN(new_n733));
  INV_X1    g0533(.A(new_n696), .ZN(new_n734));
  INV_X1    g0534(.A(G317), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT33), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n735), .A2(KEYINPUT33), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n726), .A2(new_n731), .A3(new_n733), .A4(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n723), .B(new_n739), .C1(G322), .C2(new_n720), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n693), .B1(new_n721), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n205), .A2(G355), .A3(new_n265), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n640), .A2(new_n265), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G45), .B2(new_n234), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n248), .A2(new_n429), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n742), .B1(G116), .B2(new_n205), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n691), .A2(new_n693), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n692), .A2(new_n741), .A3(new_n748), .A4(new_n686), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n688), .A2(new_n749), .ZN(G396));
  INV_X1    g0550(.A(new_n680), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n289), .A2(new_n624), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n366), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n292), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n292), .A2(new_n624), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n618), .A2(new_n619), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n598), .B1(new_n759), .B2(new_n501), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n632), .B(new_n758), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n757), .B(KEYINPUT90), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n624), .B1(new_n605), .B2(new_n612), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n751), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT91), .Z(new_n767));
  INV_X1    g0567(.A(new_n686), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(new_n751), .C2(new_n765), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n704), .B1(new_n725), .B2(G107), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n706), .A2(new_n219), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n770), .B(new_n772), .C1(new_n727), .C2(new_n709), .ZN(new_n773));
  INV_X1    g0573(.A(G294), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n381), .B1(new_n717), .B2(new_n221), .C1(new_n774), .C2(new_n719), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n777), .B2(new_n696), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n715), .A2(new_n522), .ZN(new_n779));
  INV_X1    g0579(.A(new_n717), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G143), .A2(new_n720), .B1(new_n780), .B2(G159), .ZN(new_n781));
  INV_X1    g0581(.A(G137), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n781), .B1(new_n782), .B2(new_n715), .C1(new_n342), .C2(new_n696), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT34), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n706), .A2(new_n209), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n381), .B(new_n785), .C1(G132), .C2(new_n712), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n784), .B(new_n786), .C1(new_n296), .C2(new_n724), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n702), .A2(new_n215), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n778), .A2(new_n779), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n768), .B1(new_n789), .B2(new_n693), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n693), .A2(new_n689), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n790), .B1(G77), .B2(new_n792), .C1(new_n690), .C2(new_n758), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n769), .A2(new_n793), .ZN(G384));
  INV_X1    g0594(.A(new_n622), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n390), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n412), .B(KEYINPUT17), .Z(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n798), .B2(new_n582), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n407), .A2(new_n412), .A3(new_n796), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(KEYINPUT37), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT37), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n407), .A2(new_n796), .A3(new_n802), .A4(new_n412), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT38), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n799), .A2(KEYINPUT38), .A3(new_n804), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT39), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT93), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n387), .A2(new_n389), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n398), .A2(new_n406), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n412), .B(new_n812), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n796), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n812), .B1(new_n407), .B2(new_n412), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT37), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n803), .A2(KEYINPUT94), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT95), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT94), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n822), .B(KEYINPUT37), .C1(new_n816), .C2(new_n817), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n799), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n821), .B1(new_n820), .B2(new_n823), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n806), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n808), .A2(KEYINPUT96), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT96), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n799), .A2(new_n804), .A3(new_n829), .A4(KEYINPUT38), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n811), .B1(new_n832), .B2(new_n810), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n583), .A2(new_n624), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n322), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n329), .A2(new_n624), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n583), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n329), .B(new_n624), .C1(new_n328), .C2(new_n322), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n762), .B2(new_n756), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n841), .A2(new_n809), .B1(new_n582), .B2(new_n622), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n835), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n418), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n587), .B1(new_n655), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n843), .B(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n757), .B1(new_n838), .B2(new_n839), .ZN(new_n847));
  NAND2_X1  g0647(.A1(KEYINPUT97), .A2(KEYINPUT40), .ZN(new_n848));
  INV_X1    g0648(.A(new_n502), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n600), .A2(new_n601), .A3(new_n579), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n606), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n851), .A3(new_n632), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n852), .A2(KEYINPUT31), .B1(new_n624), .B2(new_n675), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n675), .A2(KEYINPUT31), .A3(new_n624), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n847), .B(new_n848), .C1(new_n853), .C2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n808), .B2(new_n807), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n847), .B1(new_n853), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT97), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n832), .A2(new_n859), .A3(new_n856), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n857), .B1(new_n860), .B2(KEYINPUT40), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n418), .B1(new_n679), .B2(new_n854), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(G330), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n846), .B(new_n864), .Z(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n253), .B2(new_n683), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n221), .B1(new_n483), .B2(KEYINPUT35), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n867), .B(new_n231), .C1(KEYINPUT35), .C2(new_n483), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT36), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n234), .A2(new_n224), .A3(new_n374), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT92), .Z(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(G50), .B2(new_n209), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(G1), .A3(new_n346), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n866), .A2(new_n869), .A3(new_n873), .ZN(G367));
  NAND2_X1  g0674(.A1(new_n609), .A2(new_n624), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n494), .A2(new_n624), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n491), .A2(new_n497), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n637), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n497), .B1(new_n877), .B2(new_n501), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n879), .A2(KEYINPUT42), .B1(new_n632), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT100), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(KEYINPUT42), .B2(new_n879), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT43), .ZN(new_n884));
  INV_X1    g0684(.A(new_n551), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n597), .B1(new_n885), .B2(new_n632), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n590), .A2(new_n551), .A3(new_n595), .A4(new_n624), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n883), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n635), .B1(new_n877), .B2(new_n875), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(KEYINPUT98), .B(KEYINPUT43), .Z(new_n895));
  NAND2_X1  g0695(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(KEYINPUT99), .B(KEYINPUT101), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n896), .B(new_n897), .Z(new_n898));
  XNOR2_X1  g0698(.A(new_n894), .B(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  OR3_X1    g0700(.A1(new_n638), .A2(KEYINPUT44), .A3(new_n878), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n638), .A2(new_n878), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT44), .B1(new_n638), .B2(new_n878), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n638), .A2(new_n878), .A3(new_n903), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n901), .A2(new_n905), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n635), .B(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n630), .A2(KEYINPUT104), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n634), .A2(new_n636), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n637), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n911), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n681), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n641), .B(new_n916), .Z(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(KEYINPUT105), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT105), .ZN(new_n920));
  INV_X1    g0720(.A(new_n681), .ZN(new_n921));
  INV_X1    g0721(.A(new_n913), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n911), .B(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n921), .B1(new_n923), .B2(new_n909), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n920), .B1(new_n924), .B2(new_n917), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n684), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n900), .A2(new_n927), .A3(KEYINPUT106), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT106), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n685), .B1(new_n919), .B2(new_n925), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n929), .B1(new_n930), .B2(new_n899), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n715), .A2(new_n727), .B1(new_n719), .B2(new_n522), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT46), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT107), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n934), .A2(KEYINPUT107), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n935), .B(new_n936), .C1(new_n699), .C2(new_n221), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n506), .B2(new_n706), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n933), .B(new_n938), .C1(G317), .C2(new_n712), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n265), .B1(new_n732), .B2(G107), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n725), .A2(KEYINPUT46), .A3(G116), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n942), .B1(new_n777), .B2(new_n717), .C1(new_n774), .C2(new_n696), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n696), .A2(new_n710), .B1(new_n717), .B2(new_n296), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT108), .Z(new_n945));
  INV_X1    g0745(.A(new_n715), .ZN(new_n946));
  AOI22_X1  g0746(.A1(G143), .A2(new_n946), .B1(new_n730), .B2(G77), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n342), .B2(new_n719), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n265), .B1(new_n709), .B2(new_n782), .C1(new_n215), .C2(new_n699), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n209), .B2(new_n702), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n943), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT47), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n693), .ZN(new_n954));
  INV_X1    g0754(.A(new_n743), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n747), .B1(new_n205), .B2(new_n279), .C1(new_n244), .C2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n954), .A2(new_n686), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n691), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n888), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n932), .A2(new_n961), .ZN(G387));
  NAND2_X1  g0762(.A1(new_n923), .A2(new_n681), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n914), .A2(new_n921), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n963), .A2(new_n964), .A3(new_n641), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G322), .A2(new_n946), .B1(new_n734), .B2(G311), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n522), .B2(new_n717), .C1(new_n735), .C2(new_n719), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT48), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n777), .B2(new_n702), .C1(new_n774), .C2(new_n699), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT49), .Z(new_n970));
  OAI221_X1 g0770(.A(new_n381), .B1(new_n709), .B2(new_n722), .C1(new_n221), .C2(new_n706), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n719), .A2(new_n296), .B1(new_n706), .B2(new_n703), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n279), .A2(new_n702), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(new_n275), .C2(new_n734), .ZN(new_n974));
  INV_X1    g0774(.A(new_n699), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(G77), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n974), .B(new_n976), .C1(new_n710), .C2(new_n715), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n265), .B1(new_n709), .B2(new_n342), .C1(new_n209), .C2(new_n717), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n970), .A2(new_n971), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n768), .B1(new_n979), .B2(new_n693), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n640), .A2(G107), .ZN(new_n981));
  OR3_X1    g0781(.A1(new_n274), .A2(KEYINPUT50), .A3(G50), .ZN(new_n982));
  OAI21_X1  g0782(.A(KEYINPUT50), .B1(new_n274), .B2(G50), .ZN(new_n983));
  NAND2_X1  g0783(.A1(G68), .A2(G77), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n429), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n642), .B1(new_n985), .B2(new_n381), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n241), .A2(new_n429), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n986), .B1(new_n987), .B2(new_n381), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n747), .B(new_n981), .C1(new_n988), .C2(new_n640), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n980), .B(new_n989), .C1(new_n634), .C2(new_n958), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n965), .B(new_n990), .C1(new_n684), .C2(new_n914), .ZN(G393));
  AOI211_X1 g0791(.A(G41), .B(new_n640), .C1(new_n963), .C2(new_n910), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n910), .B2(new_n963), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n909), .A2(new_n685), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n747), .B1(new_n205), .B2(new_n506), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n743), .B2(new_n251), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n715), .A2(new_n342), .B1(new_n719), .B2(new_n710), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT51), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n699), .A2(new_n209), .B1(new_n717), .B2(new_n274), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G50), .B2(new_n734), .ZN(new_n1000));
  AND4_X1   g0800(.A1(new_n265), .A2(new_n998), .A3(new_n772), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n712), .A2(G143), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(new_n224), .C2(new_n702), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT109), .Z(new_n1004));
  OAI22_X1  g0804(.A1(new_n715), .A2(new_n735), .B1(new_n719), .B2(new_n727), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT52), .Z(new_n1006));
  AOI211_X1 g0806(.A(new_n265), .B(new_n1006), .C1(G294), .C2(new_n780), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n734), .A2(G303), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G283), .A2(new_n975), .B1(new_n712), .B2(G322), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT110), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G107), .B2(new_n730), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n732), .A2(G116), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1007), .A2(new_n1008), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1004), .A2(new_n1013), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n768), .B(new_n996), .C1(new_n1014), .C2(new_n693), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n958), .B2(new_n878), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n993), .A2(new_n994), .A3(new_n1016), .ZN(G390));
  AOI21_X1  g0817(.A(KEYINPUT114), .B1(new_n862), .B2(G330), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n679), .A2(new_n854), .ZN(new_n1019));
  AND4_X1   g0819(.A1(KEYINPUT114), .A2(new_n844), .A3(G330), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n845), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n755), .B1(new_n764), .B2(new_n758), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n840), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n680), .B2(new_n758), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1019), .A2(G330), .A3(new_n847), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1023), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n632), .B(new_n754), .C1(new_n650), .C2(new_n651), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n756), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT111), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1029), .A2(KEYINPUT111), .A3(new_n756), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n680), .A2(new_n758), .A3(new_n1024), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n1019), .A2(G330), .A3(new_n763), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1034), .B(new_n1035), .C1(new_n1024), .C2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1021), .B1(new_n1028), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1032), .A2(new_n1024), .A3(new_n1033), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n834), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n832), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT112), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n841), .B2(new_n834), .ZN(new_n1043));
  OAI211_X1 g0843(.A(KEYINPUT112), .B(new_n1040), .C1(new_n1022), .C2(new_n840), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1041), .B(new_n1035), .C1(new_n1045), .C2(new_n833), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(KEYINPUT113), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT39), .B1(new_n827), .B2(new_n831), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1043), .B(new_n1044), .C1(new_n1048), .C2(new_n811), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT113), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1049), .A2(new_n1050), .A3(new_n1041), .A4(new_n1035), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1041), .B1(new_n1045), .B2(new_n833), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n1027), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1038), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1047), .A2(new_n1054), .A3(new_n1051), .A4(new_n1038), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n641), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1052), .A2(new_n685), .A3(new_n1054), .ZN(new_n1059));
  XOR2_X1   g0859(.A(KEYINPUT54), .B(G143), .Z(new_n1060));
  AOI22_X1  g0860(.A1(new_n734), .A2(G137), .B1(new_n780), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT115), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G50), .B2(new_n730), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n975), .A2(G150), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT53), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n946), .A2(G128), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n712), .A2(G125), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n265), .B(new_n1067), .C1(new_n1064), .C2(KEYINPUT53), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G159), .B2(new_n732), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(G132), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n719), .A2(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n715), .A2(new_n777), .B1(new_n717), .B2(new_n506), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G107), .B2(new_n734), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT116), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n224), .B2(new_n702), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n381), .B1(new_n724), .B2(new_n219), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n709), .A2(new_n774), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n719), .A2(new_n221), .ZN(new_n1079));
  OR4_X1    g0879(.A1(new_n785), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1070), .A2(new_n1072), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n768), .B1(new_n1081), .B2(new_n693), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n275), .B2(new_n792), .C1(new_n833), .C2(new_n690), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1059), .A2(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1058), .A2(new_n1084), .ZN(G378));
  INV_X1    g0885(.A(new_n1021), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1056), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n843), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n352), .A2(new_n363), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n349), .A2(new_n795), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n857), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n828), .A2(new_n830), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n820), .A2(new_n823), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(KEYINPUT95), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1098), .A2(new_n799), .A3(new_n824), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1096), .B1(new_n1099), .B2(new_n806), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n856), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT97), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1019), .B2(new_n847), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT40), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1095), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1094), .B1(new_n1106), .B2(G330), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n861), .A2(new_n656), .A3(new_n1093), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1088), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1093), .B1(new_n861), .B2(new_n656), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n827), .A2(new_n831), .B1(new_n858), .B2(KEYINPUT97), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1105), .B1(new_n1111), .B2(new_n856), .ZN(new_n1112));
  OAI211_X1 g0912(.A(G330), .B(new_n1094), .C1(new_n1112), .C2(new_n857), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1110), .A2(new_n843), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1109), .A2(KEYINPUT57), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(KEYINPUT120), .B1(new_n1087), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT57), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1087), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1110), .A2(new_n843), .A3(new_n1113), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n843), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT120), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1056), .A2(new_n1086), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .A4(KEYINPUT57), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1116), .A2(new_n1119), .A3(new_n641), .A4(new_n1125), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1120), .A2(new_n1121), .A3(new_n684), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n976), .B1(new_n211), .B2(new_n719), .ZN(new_n1128));
  AOI211_X1 g0928(.A(G41), .B(new_n1128), .C1(G68), .C2(new_n732), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n265), .B1(new_n730), .B2(G58), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n780), .A2(new_n278), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G97), .A2(new_n734), .B1(new_n712), .B2(G283), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G116), .B2(new_n946), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1135));
  XNOR2_X1  g0935(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n296), .B1(new_n379), .B2(G41), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G128), .A2(new_n720), .B1(new_n780), .B2(G137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n975), .A2(new_n1060), .B1(new_n732), .B2(G150), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n946), .A2(G125), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G132), .B2(new_n734), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT59), .ZN(new_n1143));
  AOI21_X1  g0943(.A(G33), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(G41), .B1(new_n712), .B2(G124), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n710), .C2(new_n706), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1137), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n693), .B1(new_n1136), .B2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT118), .Z(new_n1150));
  AOI21_X1  g0950(.A(new_n768), .B1(new_n296), .B2(new_n791), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n1093), .C2(new_n690), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(KEYINPUT119), .B1(new_n1127), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT119), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n1152), .C1(new_n1118), .C2(new_n684), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1126), .A2(new_n1157), .ZN(G375));
  INV_X1    g0958(.A(new_n1038), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1021), .A2(new_n1028), .A3(new_n1037), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n918), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n684), .B1(new_n1028), .B2(new_n1037), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n840), .A2(new_n689), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n792), .A2(G68), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n265), .B1(new_n706), .B2(new_n215), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n724), .A2(new_n710), .B1(new_n1071), .B2(new_n715), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(G50), .C2(new_n732), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n734), .A2(new_n1060), .B1(new_n712), .B2(G128), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n782), .B2(new_n719), .C1(new_n342), .C2(new_n717), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n381), .B1(new_n706), .B2(new_n224), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT121), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n973), .B(new_n1172), .C1(G294), .C2(new_n946), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n734), .A2(G116), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n725), .A2(G97), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G283), .A2(new_n720), .B1(new_n712), .B2(G303), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n717), .A2(new_n211), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1170), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n768), .B(new_n1164), .C1(new_n1179), .C2(new_n693), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1162), .B1(new_n1163), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1161), .A2(new_n1181), .ZN(G381));
  INV_X1    g0982(.A(G390), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n932), .A2(new_n961), .A3(new_n1183), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1184), .A2(G396), .A3(G393), .ZN(new_n1185));
  INV_X1    g0985(.A(G384), .ZN(new_n1186));
  INV_X1    g0986(.A(G381), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(G375), .A2(G378), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(G407));
  INV_X1    g0989(.A(G213), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1188), .B2(new_n623), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(G407), .A2(new_n1191), .ZN(G409));
  NAND3_X1  g0992(.A1(new_n1126), .A2(G378), .A3(new_n1157), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(KEYINPUT122), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT122), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1126), .A2(G378), .A3(new_n1195), .A4(new_n1157), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(G378), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1122), .A2(new_n918), .A3(new_n1124), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1199), .B(new_n1152), .C1(new_n684), .C2(new_n1118), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1197), .A2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1190), .A2(G343), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT123), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1160), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT60), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT60), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1160), .A2(new_n1205), .A3(new_n1208), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1159), .A2(new_n1207), .A3(new_n641), .A4(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G384), .B1(new_n1210), .B2(new_n1181), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(G384), .A3(new_n1181), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1202), .A2(new_n1204), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(KEYINPUT124), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1203), .A2(G2897), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT124), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1212), .A2(new_n1219), .A3(new_n1213), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1220), .A2(new_n1218), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT63), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1216), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(G387), .A2(G390), .ZN(new_n1228));
  XOR2_X1   g1028(.A(G393), .B(G396), .Z(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1184), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1183), .B1(new_n932), .B2(new_n961), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n960), .B(G390), .C1(new_n928), .C2(new_n931), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1229), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT61), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1231), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1202), .A2(KEYINPUT63), .A3(new_n1204), .A4(new_n1215), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT125), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1194), .A2(new_n1196), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1239), .A2(new_n1203), .A3(new_n1214), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT125), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1241), .A3(KEYINPUT63), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1227), .A2(new_n1236), .A3(new_n1238), .A4(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1223), .B1(new_n1239), .B2(new_n1203), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT62), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1245), .B1(new_n1240), .B2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1202), .A2(new_n1246), .A3(new_n1204), .A4(new_n1215), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1235), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1244), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1243), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT126), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1243), .A2(new_n1250), .A3(KEYINPUT126), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(G405));
  NAND2_X1  g1055(.A1(G375), .A2(new_n1198), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1197), .A2(new_n1256), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(new_n1214), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(KEYINPUT127), .B2(new_n1244), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1244), .A2(KEYINPUT127), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1259), .B(new_n1260), .Z(G402));
endmodule


