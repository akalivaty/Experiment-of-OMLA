

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U557 ( .A(KEYINPUT86), .B(n537), .ZN(G164) );
  NOR2_X2 U558 ( .A1(n532), .A2(G2105), .ZN(n538) );
  INV_X2 U559 ( .A(G2104), .ZN(n532) );
  NOR2_X2 U560 ( .A1(G1384), .A2(G164), .ZN(n782) );
  INV_X1 U561 ( .A(n738), .ZN(n722) );
  BUF_X1 U562 ( .A(n621), .Z(n622) );
  XNOR2_X1 U563 ( .A(n539), .B(KEYINPUT66), .ZN(n540) );
  XNOR2_X1 U564 ( .A(n526), .B(KEYINPUT65), .ZN(n619) );
  INV_X1 U565 ( .A(KEYINPUT97), .ZN(n714) );
  NOR2_X1 U566 ( .A1(n766), .A2(n765), .ZN(n767) );
  AND2_X1 U567 ( .A1(n692), .A2(G40), .ZN(n780) );
  XNOR2_X1 U568 ( .A(n541), .B(n540), .ZN(n543) );
  NOR2_X1 U569 ( .A1(n587), .A2(n586), .ZN(n589) );
  AND2_X1 U570 ( .A1(n821), .A2(n812), .ZN(n522) );
  AND2_X1 U571 ( .A1(n522), .A2(n813), .ZN(n523) );
  OR2_X1 U572 ( .A1(n778), .A2(n777), .ZN(n524) );
  NOR2_X1 U573 ( .A1(n778), .A2(n760), .ZN(n525) );
  AND2_X1 U574 ( .A1(n738), .A2(G1341), .ZN(n694) );
  NOR2_X1 U575 ( .A1(n710), .A2(n709), .ZN(n716) );
  INV_X1 U576 ( .A(KEYINPUT32), .ZN(n747) );
  INV_X1 U577 ( .A(n992), .ZN(n765) );
  INV_X1 U578 ( .A(KEYINPUT68), .ZN(n527) );
  XNOR2_X1 U579 ( .A(n527), .B(KEYINPUT17), .ZN(n529) );
  XNOR2_X1 U580 ( .A(n529), .B(n528), .ZN(n621) );
  BUF_X1 U581 ( .A(n619), .Z(n891) );
  BUF_X1 U582 ( .A(n538), .Z(n896) );
  XNOR2_X1 U583 ( .A(n599), .B(n598), .ZN(n996) );
  NAND2_X1 U584 ( .A1(n589), .A2(n588), .ZN(n985) );
  NAND2_X1 U585 ( .A1(n532), .A2(G2105), .ZN(n526) );
  NAND2_X1 U586 ( .A1(G126), .A2(n619), .ZN(n531) );
  NOR2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n621), .A2(G138), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n531), .A2(n530), .ZN(n536) );
  NAND2_X1 U590 ( .A1(G102), .A2(n896), .ZN(n534) );
  AND2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n892) );
  NAND2_X1 U592 ( .A1(G114), .A2(n892), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U595 ( .A1(G101), .A2(n538), .ZN(n541) );
  INV_X1 U596 ( .A(KEYINPUT23), .ZN(n539) );
  NAND2_X1 U597 ( .A1(G125), .A2(n619), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n545) );
  INV_X1 U599 ( .A(KEYINPUT67), .ZN(n544) );
  XNOR2_X1 U600 ( .A(n545), .B(n544), .ZN(n549) );
  NAND2_X1 U601 ( .A1(n892), .A2(G113), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G137), .A2(n621), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U605 ( .A(n550), .B(KEYINPUT64), .ZN(n692) );
  BUF_X1 U606 ( .A(n692), .Z(G160) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  INV_X1 U611 ( .A(G651), .ZN(n555) );
  NOR2_X1 U612 ( .A1(G543), .A2(n555), .ZN(n551) );
  XOR2_X2 U613 ( .A(KEYINPUT1), .B(n551), .Z(n657) );
  NAND2_X1 U614 ( .A1(G64), .A2(n657), .ZN(n553) );
  XOR2_X1 U615 ( .A(KEYINPUT0), .B(G543), .Z(n654) );
  NOR2_X2 U616 ( .A1(n654), .A2(G651), .ZN(n665) );
  NAND2_X1 U617 ( .A1(G52), .A2(n665), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U619 ( .A(KEYINPUT71), .B(n554), .Z(n560) );
  NOR2_X2 U620 ( .A1(G543), .A2(G651), .ZN(n658) );
  NAND2_X1 U621 ( .A1(G90), .A2(n658), .ZN(n557) );
  NOR2_X4 U622 ( .A1(n654), .A2(n555), .ZN(n661) );
  NAND2_X1 U623 ( .A1(G77), .A2(n661), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(G171) );
  NAND2_X1 U627 ( .A1(n658), .A2(G88), .ZN(n563) );
  NAND2_X1 U628 ( .A1(G75), .A2(n661), .ZN(n561) );
  XOR2_X1 U629 ( .A(KEYINPUT83), .B(n561), .Z(n562) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G62), .A2(n657), .ZN(n565) );
  NAND2_X1 U632 ( .A1(G50), .A2(n665), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U634 ( .A1(n567), .A2(n566), .ZN(G166) );
  NAND2_X1 U635 ( .A1(G63), .A2(n657), .ZN(n569) );
  NAND2_X1 U636 ( .A1(G51), .A2(n665), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U638 ( .A(KEYINPUT6), .B(n570), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n658), .A2(G89), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n571), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U641 ( .A1(G76), .A2(n661), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U643 ( .A(n574), .B(KEYINPUT5), .Z(n575) );
  NOR2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U645 ( .A(KEYINPUT7), .B(n577), .Z(n578) );
  XNOR2_X1 U646 ( .A(KEYINPUT78), .B(n578), .ZN(G168) );
  XOR2_X1 U647 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U648 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U649 ( .A(n579), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U650 ( .A(G223), .ZN(n842) );
  NAND2_X1 U651 ( .A1(n842), .A2(G567), .ZN(n580) );
  XOR2_X1 U652 ( .A(KEYINPUT11), .B(n580), .Z(G234) );
  NAND2_X1 U653 ( .A1(G56), .A2(n657), .ZN(n581) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(n581), .Z(n587) );
  NAND2_X1 U655 ( .A1(n658), .A2(G81), .ZN(n582) );
  XNOR2_X1 U656 ( .A(n582), .B(KEYINPUT12), .ZN(n584) );
  NAND2_X1 U657 ( .A1(G68), .A2(n661), .ZN(n583) );
  NAND2_X1 U658 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U659 ( .A(KEYINPUT13), .B(n585), .Z(n586) );
  NAND2_X1 U660 ( .A1(n665), .A2(G43), .ZN(n588) );
  INV_X1 U661 ( .A(G860), .ZN(n613) );
  OR2_X1 U662 ( .A1(n985), .A2(n613), .ZN(G153) );
  INV_X1 U663 ( .A(G171), .ZN(G301) );
  NAND2_X1 U664 ( .A1(G868), .A2(G301), .ZN(n601) );
  XNOR2_X1 U665 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n599) );
  NAND2_X1 U666 ( .A1(G54), .A2(n665), .ZN(n590) );
  XNOR2_X1 U667 ( .A(n590), .B(KEYINPUT76), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G66), .A2(n657), .ZN(n592) );
  NAND2_X1 U669 ( .A1(G92), .A2(n658), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U671 ( .A1(G79), .A2(n661), .ZN(n593) );
  XNOR2_X1 U672 ( .A(KEYINPUT75), .B(n593), .ZN(n594) );
  NOR2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n598) );
  INV_X1 U675 ( .A(G868), .ZN(n610) );
  NAND2_X1 U676 ( .A1(n996), .A2(n610), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(G284) );
  NAND2_X1 U678 ( .A1(G91), .A2(n658), .ZN(n602) );
  XNOR2_X1 U679 ( .A(n602), .B(KEYINPUT72), .ZN(n605) );
  NAND2_X1 U680 ( .A1(G53), .A2(n665), .ZN(n603) );
  XOR2_X1 U681 ( .A(KEYINPUT73), .B(n603), .Z(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U683 ( .A1(G65), .A2(n657), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G78), .A2(n661), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n973) );
  XOR2_X1 U687 ( .A(KEYINPUT74), .B(n973), .Z(G299) );
  NAND2_X1 U688 ( .A1(G868), .A2(G286), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G299), .A2(n610), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(G297) );
  NAND2_X1 U691 ( .A1(n613), .A2(G559), .ZN(n614) );
  INV_X1 U692 ( .A(n996), .ZN(n912) );
  NAND2_X1 U693 ( .A1(n614), .A2(n912), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n615), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U695 ( .A1(G868), .A2(n985), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n912), .A2(G868), .ZN(n616) );
  NOR2_X1 U697 ( .A1(G559), .A2(n616), .ZN(n617) );
  NOR2_X1 U698 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U699 ( .A1(G123), .A2(n891), .ZN(n620) );
  XNOR2_X1 U700 ( .A(n620), .B(KEYINPUT18), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G99), .A2(n896), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G135), .A2(n622), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G111), .A2(n892), .ZN(n625) );
  XNOR2_X1 U705 ( .A(KEYINPUT79), .B(n625), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U708 ( .A(KEYINPUT80), .B(n630), .Z(n932) );
  XNOR2_X1 U709 ( .A(n932), .B(G2096), .ZN(n632) );
  INV_X1 U710 ( .A(G2100), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(G156) );
  NAND2_X1 U712 ( .A1(G559), .A2(n912), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n985), .B(n633), .ZN(n676) );
  NOR2_X1 U714 ( .A1(n676), .A2(G860), .ZN(n642) );
  NAND2_X1 U715 ( .A1(n661), .A2(G80), .ZN(n634) );
  XOR2_X1 U716 ( .A(KEYINPUT81), .B(n634), .Z(n636) );
  NAND2_X1 U717 ( .A1(n658), .A2(G93), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U719 ( .A(KEYINPUT82), .B(n637), .ZN(n641) );
  NAND2_X1 U720 ( .A1(G67), .A2(n657), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G55), .A2(n665), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n669) );
  XNOR2_X1 U724 ( .A(n642), .B(n669), .ZN(G145) );
  NAND2_X1 U725 ( .A1(G60), .A2(n657), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G47), .A2(n665), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U728 ( .A(KEYINPUT70), .B(n645), .ZN(n648) );
  NAND2_X1 U729 ( .A1(G85), .A2(n658), .ZN(n646) );
  XNOR2_X1 U730 ( .A(KEYINPUT69), .B(n646), .ZN(n647) );
  NOR2_X1 U731 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n661), .A2(G72), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n650), .A2(n649), .ZN(G290) );
  NAND2_X1 U734 ( .A1(G49), .A2(n665), .ZN(n652) );
  NAND2_X1 U735 ( .A1(G74), .A2(G651), .ZN(n651) );
  NAND2_X1 U736 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U737 ( .A1(n657), .A2(n653), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n654), .A2(G87), .ZN(n655) );
  NAND2_X1 U739 ( .A1(n656), .A2(n655), .ZN(G288) );
  NAND2_X1 U740 ( .A1(G61), .A2(n657), .ZN(n660) );
  NAND2_X1 U741 ( .A1(G86), .A2(n658), .ZN(n659) );
  NAND2_X1 U742 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n661), .A2(G73), .ZN(n662) );
  XOR2_X1 U744 ( .A(KEYINPUT2), .B(n662), .Z(n663) );
  NOR2_X1 U745 ( .A1(n664), .A2(n663), .ZN(n667) );
  NAND2_X1 U746 ( .A1(n665), .A2(G48), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n667), .A2(n666), .ZN(G305) );
  NOR2_X1 U748 ( .A1(G868), .A2(n669), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n668), .B(KEYINPUT85), .ZN(n679) );
  XNOR2_X1 U750 ( .A(G299), .B(n669), .ZN(n675) );
  XNOR2_X1 U751 ( .A(KEYINPUT84), .B(G290), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n670), .B(G288), .ZN(n671) );
  XNOR2_X1 U753 ( .A(KEYINPUT19), .B(n671), .ZN(n673) );
  XNOR2_X1 U754 ( .A(G305), .B(G166), .ZN(n672) );
  XNOR2_X1 U755 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U756 ( .A(n675), .B(n674), .ZN(n911) );
  XOR2_X1 U757 ( .A(n911), .B(n676), .Z(n677) );
  NAND2_X1 U758 ( .A1(G868), .A2(n677), .ZN(n678) );
  NAND2_X1 U759 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U760 ( .A1(G2078), .A2(G2084), .ZN(n680) );
  XOR2_X1 U761 ( .A(KEYINPUT20), .B(n680), .Z(n681) );
  NAND2_X1 U762 ( .A1(G2090), .A2(n681), .ZN(n682) );
  XNOR2_X1 U763 ( .A(KEYINPUT21), .B(n682), .ZN(n683) );
  NAND2_X1 U764 ( .A1(n683), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n684) );
  XOR2_X1 U767 ( .A(KEYINPUT22), .B(n684), .Z(n685) );
  NOR2_X1 U768 ( .A1(G218), .A2(n685), .ZN(n686) );
  NAND2_X1 U769 ( .A1(G96), .A2(n686), .ZN(n847) );
  NAND2_X1 U770 ( .A1(n847), .A2(G2106), .ZN(n690) );
  NAND2_X1 U771 ( .A1(G69), .A2(G120), .ZN(n687) );
  NOR2_X1 U772 ( .A1(G237), .A2(n687), .ZN(n688) );
  NAND2_X1 U773 ( .A1(G108), .A2(n688), .ZN(n848) );
  NAND2_X1 U774 ( .A1(n848), .A2(G567), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n690), .A2(n689), .ZN(n849) );
  NAND2_X1 U776 ( .A1(G661), .A2(G483), .ZN(n691) );
  NOR2_X1 U777 ( .A1(n849), .A2(n691), .ZN(n846) );
  NAND2_X1 U778 ( .A1(n846), .A2(G36), .ZN(G176) );
  INV_X1 U779 ( .A(G166), .ZN(G303) );
  NAND2_X2 U780 ( .A1(n782), .A2(n780), .ZN(n738) );
  NAND2_X1 U781 ( .A1(G1996), .A2(n722), .ZN(n693) );
  XNOR2_X1 U782 ( .A(n693), .B(KEYINPUT26), .ZN(n703) );
  NOR2_X2 U783 ( .A1(n694), .A2(n985), .ZN(n702) );
  AND2_X1 U784 ( .A1(n702), .A2(n912), .ZN(n695) );
  NAND2_X1 U785 ( .A1(n703), .A2(n695), .ZN(n696) );
  XNOR2_X1 U786 ( .A(n696), .B(KEYINPUT94), .ZN(n701) );
  INV_X1 U787 ( .A(G2067), .ZN(n953) );
  NOR2_X1 U788 ( .A1(n738), .A2(n953), .ZN(n697) );
  XNOR2_X1 U789 ( .A(n697), .B(KEYINPUT95), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n738), .A2(G1348), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n706) );
  NAND2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U794 ( .A1(n996), .A2(n704), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n706), .A2(n705), .ZN(n713) );
  NAND2_X1 U796 ( .A1(n722), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U797 ( .A(KEYINPUT27), .B(n707), .ZN(n710) );
  NAND2_X1 U798 ( .A1(G1956), .A2(n738), .ZN(n708) );
  XNOR2_X1 U799 ( .A(KEYINPUT93), .B(n708), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n716), .A2(n973), .ZN(n711) );
  XNOR2_X1 U801 ( .A(n711), .B(KEYINPUT96), .ZN(n712) );
  NAND2_X1 U802 ( .A1(n713), .A2(n712), .ZN(n715) );
  XNOR2_X1 U803 ( .A(n715), .B(n714), .ZN(n719) );
  OR2_X1 U804 ( .A1(n973), .A2(n716), .ZN(n717) );
  XNOR2_X1 U805 ( .A(KEYINPUT28), .B(n717), .ZN(n718) );
  NAND2_X1 U806 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U807 ( .A(n720), .B(KEYINPUT29), .ZN(n726) );
  XOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .Z(n956) );
  NOR2_X1 U809 ( .A1(n956), .A2(n738), .ZN(n721) );
  XNOR2_X1 U810 ( .A(n721), .B(KEYINPUT92), .ZN(n724) );
  NOR2_X1 U811 ( .A1(n722), .A2(G1961), .ZN(n723) );
  NOR2_X1 U812 ( .A1(n724), .A2(n723), .ZN(n730) );
  NOR2_X1 U813 ( .A1(G301), .A2(n730), .ZN(n725) );
  NOR2_X1 U814 ( .A1(n726), .A2(n725), .ZN(n735) );
  NAND2_X1 U815 ( .A1(G8), .A2(n738), .ZN(n778) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n778), .ZN(n752) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n738), .ZN(n749) );
  NOR2_X1 U818 ( .A1(n752), .A2(n749), .ZN(n727) );
  NAND2_X1 U819 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n728), .ZN(n729) );
  NOR2_X1 U821 ( .A1(G168), .A2(n729), .ZN(n732) );
  AND2_X1 U822 ( .A1(G301), .A2(n730), .ZN(n731) );
  NOR2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U824 ( .A(n733), .B(KEYINPUT31), .ZN(n734) );
  NOR2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n737) );
  INV_X1 U826 ( .A(KEYINPUT98), .ZN(n736) );
  XNOR2_X1 U827 ( .A(n737), .B(n736), .ZN(n750) );
  NAND2_X1 U828 ( .A1(n750), .A2(G286), .ZN(n746) );
  INV_X1 U829 ( .A(G8), .ZN(n744) );
  NOR2_X1 U830 ( .A1(G2090), .A2(n738), .ZN(n739) );
  XNOR2_X1 U831 ( .A(KEYINPUT99), .B(n739), .ZN(n742) );
  NOR2_X1 U832 ( .A1(G1971), .A2(n778), .ZN(n740) );
  NOR2_X1 U833 ( .A1(G166), .A2(n740), .ZN(n741) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n743) );
  OR2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n748) );
  XNOR2_X1 U837 ( .A(n748), .B(n747), .ZN(n756) );
  NAND2_X1 U838 ( .A1(G8), .A2(n749), .ZN(n754) );
  INV_X1 U839 ( .A(n750), .ZN(n751) );
  NOR2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n756), .A2(n755), .ZN(n771) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n976) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n757) );
  NOR2_X1 U845 ( .A1(n976), .A2(n757), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n771), .A2(n758), .ZN(n759) );
  XNOR2_X1 U847 ( .A(n759), .B(KEYINPUT100), .ZN(n761) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n977) );
  INV_X1 U849 ( .A(n977), .ZN(n760) );
  AND2_X1 U850 ( .A1(n761), .A2(n525), .ZN(n762) );
  NOR2_X1 U851 ( .A1(n762), .A2(KEYINPUT33), .ZN(n763) );
  INV_X1 U852 ( .A(n763), .ZN(n768) );
  NAND2_X1 U853 ( .A1(n976), .A2(KEYINPUT33), .ZN(n764) );
  NOR2_X1 U854 ( .A1(n764), .A2(n778), .ZN(n766) );
  XOR2_X1 U855 ( .A(G1981), .B(G305), .Z(n992) );
  NAND2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n774) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U858 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n772), .A2(n778), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U862 ( .A(n775), .B(KEYINPUT101), .ZN(n779) );
  NOR2_X1 U863 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U864 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NAND2_X1 U865 ( .A1(n779), .A2(n524), .ZN(n814) );
  INV_X1 U866 ( .A(n780), .ZN(n781) );
  NOR2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n825) );
  XNOR2_X1 U868 ( .A(G2067), .B(KEYINPUT37), .ZN(n823) );
  NAND2_X1 U869 ( .A1(n896), .A2(G104), .ZN(n783) );
  XOR2_X1 U870 ( .A(KEYINPUT87), .B(n783), .Z(n785) );
  NAND2_X1 U871 ( .A1(G140), .A2(n622), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U873 ( .A(KEYINPUT34), .B(n786), .ZN(n794) );
  NAND2_X1 U874 ( .A1(n892), .A2(G116), .ZN(n787) );
  XNOR2_X1 U875 ( .A(KEYINPUT89), .B(n787), .ZN(n790) );
  NAND2_X1 U876 ( .A1(n891), .A2(G128), .ZN(n788) );
  XOR2_X1 U877 ( .A(n788), .B(KEYINPUT88), .Z(n789) );
  NOR2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U879 ( .A(KEYINPUT35), .B(n791), .Z(n792) );
  XOR2_X1 U880 ( .A(KEYINPUT90), .B(n792), .Z(n793) );
  NOR2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U882 ( .A(KEYINPUT36), .B(n795), .ZN(n908) );
  NOR2_X1 U883 ( .A1(n823), .A2(n908), .ZN(n944) );
  NAND2_X1 U884 ( .A1(n825), .A2(n944), .ZN(n821) );
  NAND2_X1 U885 ( .A1(G95), .A2(n896), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G131), .A2(n622), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G119), .A2(n891), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G107), .A2(n892), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n877) );
  INV_X1 U892 ( .A(G1991), .ZN(n952) );
  NOR2_X1 U893 ( .A1(n877), .A2(n952), .ZN(n810) );
  NAND2_X1 U894 ( .A1(G129), .A2(n891), .ZN(n803) );
  NAND2_X1 U895 ( .A1(G141), .A2(n622), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n896), .A2(G105), .ZN(n804) );
  XOR2_X1 U898 ( .A(KEYINPUT38), .B(n804), .Z(n805) );
  NOR2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n892), .A2(G117), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n902) );
  AND2_X1 U902 ( .A1(G1996), .A2(n902), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n924) );
  XNOR2_X1 U904 ( .A(KEYINPUT91), .B(n825), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n924), .A2(n811), .ZN(n818) );
  INV_X1 U906 ( .A(n818), .ZN(n812) );
  XNOR2_X1 U907 ( .A(G1986), .B(G290), .ZN(n981) );
  NAND2_X1 U908 ( .A1(n981), .A2(n825), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n814), .A2(n523), .ZN(n828) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n902), .ZN(n928) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n952), .A2(n877), .ZN(n923) );
  INV_X1 U913 ( .A(n923), .ZN(n815) );
  NOR2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U916 ( .A1(n928), .A2(n819), .ZN(n820) );
  XNOR2_X1 U917 ( .A(KEYINPUT39), .B(n820), .ZN(n822) );
  NAND2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n823), .A2(n908), .ZN(n941) );
  NAND2_X1 U920 ( .A1(n824), .A2(n941), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U923 ( .A(n829), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U924 ( .A(G1348), .B(G1341), .ZN(n830) );
  XNOR2_X1 U925 ( .A(n830), .B(G2451), .ZN(n840) );
  XOR2_X1 U926 ( .A(G2435), .B(G2430), .Z(n832) );
  XNOR2_X1 U927 ( .A(G2454), .B(G2438), .ZN(n831) );
  XNOR2_X1 U928 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U929 ( .A(G2427), .B(KEYINPUT103), .Z(n834) );
  XNOR2_X1 U930 ( .A(G2443), .B(G2446), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U932 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U933 ( .A(KEYINPUT104), .B(KEYINPUT102), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U935 ( .A(n840), .B(n839), .ZN(n841) );
  NAND2_X1 U936 ( .A1(n841), .A2(G14), .ZN(n917) );
  XNOR2_X1 U937 ( .A(KEYINPUT105), .B(n917), .ZN(G401) );
  NAND2_X1 U938 ( .A1(n842), .A2(G2106), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n843), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U941 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U943 ( .A1(n846), .A2(n845), .ZN(G188) );
  XNOR2_X1 U944 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  NOR2_X1 U945 ( .A1(n848), .A2(n847), .ZN(G325) );
  XOR2_X1 U946 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U948 ( .A(G120), .ZN(G236) );
  INV_X1 U949 ( .A(G69), .ZN(G235) );
  INV_X1 U950 ( .A(n849), .ZN(G319) );
  XOR2_X1 U951 ( .A(G2100), .B(G2096), .Z(n851) );
  XNOR2_X1 U952 ( .A(KEYINPUT42), .B(G2678), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U954 ( .A(KEYINPUT43), .B(G2072), .Z(n853) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2090), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U957 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U958 ( .A(G2078), .B(G2084), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(G227) );
  XOR2_X1 U960 ( .A(G1976), .B(G1971), .Z(n859) );
  XNOR2_X1 U961 ( .A(G1986), .B(G1956), .ZN(n858) );
  XNOR2_X1 U962 ( .A(n859), .B(n858), .ZN(n869) );
  XOR2_X1 U963 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n861) );
  XNOR2_X1 U964 ( .A(G1996), .B(KEYINPUT111), .ZN(n860) );
  XNOR2_X1 U965 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U966 ( .A(G1961), .B(G1966), .Z(n863) );
  XNOR2_X1 U967 ( .A(G1991), .B(G1981), .ZN(n862) );
  XNOR2_X1 U968 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U969 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U970 ( .A(KEYINPUT110), .B(G2474), .ZN(n866) );
  XNOR2_X1 U971 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U972 ( .A(n869), .B(n868), .Z(G229) );
  NAND2_X1 U973 ( .A1(G100), .A2(n896), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G112), .A2(n892), .ZN(n870) );
  NAND2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n891), .A2(G124), .ZN(n872) );
  XNOR2_X1 U977 ( .A(n872), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U978 ( .A1(G136), .A2(n622), .ZN(n873) );
  NAND2_X1 U979 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U980 ( .A1(n876), .A2(n875), .ZN(G162) );
  XNOR2_X1 U981 ( .A(n877), .B(G164), .ZN(n878) );
  XNOR2_X1 U982 ( .A(n878), .B(G160), .ZN(n882) );
  XOR2_X1 U983 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n880) );
  XNOR2_X1 U984 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n879) );
  XNOR2_X1 U985 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U986 ( .A(n882), .B(n881), .Z(n907) );
  NAND2_X1 U987 ( .A1(G130), .A2(n891), .ZN(n884) );
  NAND2_X1 U988 ( .A1(G118), .A2(n892), .ZN(n883) );
  NAND2_X1 U989 ( .A1(n884), .A2(n883), .ZN(n889) );
  NAND2_X1 U990 ( .A1(G106), .A2(n896), .ZN(n886) );
  NAND2_X1 U991 ( .A1(G142), .A2(n622), .ZN(n885) );
  NAND2_X1 U992 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U993 ( .A(n887), .B(KEYINPUT45), .Z(n888) );
  NOR2_X1 U994 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U995 ( .A(n890), .B(n932), .ZN(n905) );
  NAND2_X1 U996 ( .A1(G127), .A2(n891), .ZN(n894) );
  NAND2_X1 U997 ( .A1(G115), .A2(n892), .ZN(n893) );
  NAND2_X1 U998 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U999 ( .A(n895), .B(KEYINPUT47), .ZN(n898) );
  NAND2_X1 U1000 ( .A1(G103), .A2(n896), .ZN(n897) );
  NAND2_X1 U1001 ( .A1(n898), .A2(n897), .ZN(n901) );
  NAND2_X1 U1002 ( .A1(n622), .A2(G139), .ZN(n899) );
  XOR2_X1 U1003 ( .A(KEYINPUT112), .B(n899), .Z(n900) );
  NOR2_X1 U1004 ( .A1(n901), .A2(n900), .ZN(n935) );
  XOR2_X1 U1005 ( .A(n902), .B(n935), .Z(n903) );
  XNOR2_X1 U1006 ( .A(n903), .B(G162), .ZN(n904) );
  XNOR2_X1 U1007 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1009 ( .A(n909), .B(n908), .Z(n910) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1011 ( .A(n985), .B(n911), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(G171), .B(n912), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n915), .B(G286), .ZN(n916) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n916), .ZN(G397) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n917), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n926) );
  XOR2_X1 U1025 ( .A(G2084), .B(G160), .Z(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(G2090), .B(G162), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(n927), .B(KEYINPUT115), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(KEYINPUT51), .B(n930), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n940) );
  XOR2_X1 U1033 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1036 ( .A(KEYINPUT50), .B(n938), .Z(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(KEYINPUT52), .B(n945), .ZN(n946) );
  XOR2_X1 U1041 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n967) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n967), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n947), .A2(G29), .ZN(n1033) );
  XOR2_X1 U1044 ( .A(G2072), .B(G33), .Z(n948) );
  NAND2_X1 U1045 ( .A1(n948), .A2(G28), .ZN(n951) );
  XOR2_X1 U1046 ( .A(KEYINPUT117), .B(G1996), .Z(n949) );
  XNOR2_X1 U1047 ( .A(G32), .B(n949), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n960) );
  XNOR2_X1 U1049 ( .A(n952), .B(G25), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n953), .B(G26), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G27), .B(n956), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n961), .B(KEYINPUT53), .ZN(n964) );
  XOR2_X1 U1056 ( .A(G2084), .B(G34), .Z(n962) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n962), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(G35), .B(G2090), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1061 ( .A(KEYINPUT118), .B(n967), .Z(n968) );
  XNOR2_X1 U1062 ( .A(n969), .B(n968), .ZN(n971) );
  INV_X1 U1063 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n972), .A2(G11), .ZN(n1031) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  XOR2_X1 U1067 ( .A(n973), .B(G1956), .Z(n975) );
  XOR2_X1 U1068 ( .A(G166), .B(G1971), .Z(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n983) );
  INV_X1 U1070 ( .A(n976), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(KEYINPUT120), .B(n979), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(n984), .B(KEYINPUT121), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(G301), .B(G1961), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(n985), .B(G1341), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n995) );
  XOR2_X1 U1080 ( .A(G1966), .B(KEYINPUT119), .Z(n990) );
  XNOR2_X1 U1081 ( .A(G168), .B(n990), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1083 ( .A(KEYINPUT57), .B(n993), .Z(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n998) );
  XOR2_X1 U1085 ( .A(G1348), .B(n996), .Z(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1029) );
  INV_X1 U1088 ( .A(G16), .ZN(n1027) );
  XOR2_X1 U1089 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n1025) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G21), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(G5), .B(G1961), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1023) );
  XNOR2_X1 U1093 ( .A(G1981), .B(G6), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G1341), .B(G19), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1096 ( .A(KEYINPUT122), .B(n1005), .Z(n1007) );
  XNOR2_X1 U1097 ( .A(G1956), .B(G20), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1099 ( .A(KEYINPUT123), .B(n1008), .Z(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT59), .B(G4), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(n1009), .B(KEYINPUT124), .ZN(n1010) );
  XNOR2_X1 U1102 ( .A(G1348), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n1013) );
  XNOR2_X1 U1105 ( .A(n1014), .B(n1013), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1016) );
  XNOR2_X1 U1107 ( .A(G23), .B(G1976), .ZN(n1015) );
  NOR2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XOR2_X1 U1109 ( .A(G1986), .B(G24), .Z(n1017) );
  NAND2_X1 U1110 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1114 ( .A(n1025), .B(n1024), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1119 ( .A(n1034), .B(KEYINPUT62), .ZN(n1035) );
  XNOR2_X1 U1120 ( .A(KEYINPUT127), .B(n1035), .ZN(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

