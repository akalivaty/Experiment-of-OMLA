//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n599, new_n601, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT64), .Z(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G137), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n465), .A2(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n464), .A2(new_n466), .B1(new_n467), .B2(G101), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(new_n465), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  XNOR2_X1  g046(.A(new_n464), .B(KEYINPUT65), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n465), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT66), .Z(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n472), .A2(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G124), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(G126), .A2(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G102), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(new_n465), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n485), .B2(new_n486), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n495), .B(new_n498), .C1(new_n486), .C2(new_n485), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(G164));
  NAND3_X1  g075(.A1(KEYINPUT67), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(G543), .B1(KEYINPUT67), .B2(KEYINPUT5), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OAI21_X1  g083(.A(G543), .B1(new_n504), .B2(new_n505), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(G62), .B1(new_n502), .B2(new_n503), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n510), .A2(new_n514), .ZN(G166));
  XOR2_X1   g090(.A(KEYINPUT68), .B(KEYINPUT7), .Z(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n509), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G51), .ZN(new_n520));
  INV_X1    g095(.A(new_n503), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(new_n501), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n518), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n506), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n511), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n506), .A2(new_n530), .B1(new_n531), .B2(new_n509), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G171));
  AOI22_X1  g108(.A1(new_n525), .A2(G81), .B1(G43), .B2(new_n519), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT70), .ZN(new_n535));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n502), .A2(new_n503), .ZN(new_n537));
  INV_X1    g112(.A(G56), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n511), .B1(new_n539), .B2(KEYINPUT69), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n540), .B1(KEYINPUT69), .B2(new_n539), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n535), .A2(G860), .A3(new_n541), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT71), .ZN(G188));
  NAND2_X1  g122(.A1(new_n519), .A2(G53), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G65), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n537), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G651), .B1(new_n525), .B2(G91), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G299));
  INV_X1    g129(.A(G171), .ZN(G301));
  INV_X1    g130(.A(G168), .ZN(G286));
  INV_X1    g131(.A(G166), .ZN(G303));
  NAND2_X1  g132(.A1(new_n525), .A2(G87), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n519), .A2(G49), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(G288));
  INV_X1    g136(.A(G86), .ZN(new_n562));
  INV_X1    g137(.A(G48), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n506), .A2(new_n562), .B1(new_n563), .B2(new_n509), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(G61), .B1(new_n502), .B2(new_n503), .ZN(new_n566));
  NAND2_X1  g141(.A1(G73), .A2(G543), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n511), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI211_X1 g145(.A(KEYINPUT72), .B(new_n511), .C1(new_n566), .C2(new_n567), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n565), .B1(new_n570), .B2(new_n571), .ZN(G305));
  AOI22_X1  g147(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n511), .ZN(new_n574));
  INV_X1    g149(.A(G85), .ZN(new_n575));
  INV_X1    g150(.A(G47), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n506), .A2(new_n575), .B1(new_n576), .B2(new_n509), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G290));
  INV_X1    g154(.A(G868), .ZN(new_n580));
  NOR2_X1   g155(.A1(G301), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n525), .A2(G92), .ZN(new_n582));
  XOR2_X1   g157(.A(KEYINPUT73), .B(KEYINPUT10), .Z(new_n583));
  XNOR2_X1  g158(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G79), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G66), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n537), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(new_n519), .B2(G54), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(KEYINPUT74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(KEYINPUT74), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n581), .B1(new_n593), .B2(new_n580), .ZN(G284));
  AOI21_X1  g169(.A(new_n581), .B1(new_n593), .B2(new_n580), .ZN(G321));
  NAND2_X1  g170(.A1(G299), .A2(new_n580), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(G168), .B2(new_n580), .ZN(G297));
  OAI21_X1  g172(.A(new_n596), .B1(G168), .B2(new_n580), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n593), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n535), .A2(new_n541), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n592), .A2(KEYINPUT75), .A3(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT75), .B1(new_n592), .B2(G559), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  MUX2_X1   g179(.A(new_n601), .B(new_n604), .S(G868), .Z(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g181(.A(G111), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n607), .A2(KEYINPUT77), .A3(G2105), .ZN(new_n608));
  AOI21_X1  g183(.A(KEYINPUT77), .B1(new_n607), .B2(G2105), .ZN(new_n609));
  OAI21_X1  g184(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n474), .A2(G135), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT76), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n480), .A2(new_n613), .A3(G123), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n480), .B2(G123), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(G2096), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(G2096), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n464), .A2(new_n467), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(G156));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT14), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n627), .B(new_n633), .Z(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(G14), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n635), .ZN(G401));
  XOR2_X1   g214(.A(G2072), .B(G2078), .Z(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(KEYINPUT78), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(KEYINPUT78), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n640), .B(KEYINPUT17), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n647), .C1(new_n648), .C2(new_n644), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT79), .Z(new_n650));
  NOR3_X1   g225(.A1(new_n647), .A2(new_n640), .A3(new_n644), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT18), .Z(new_n652));
  NOR2_X1   g227(.A1(new_n647), .A2(new_n643), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n652), .B1(new_n648), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2096), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n662), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT20), .Z(new_n666));
  AOI211_X1 g241(.A(new_n664), .B(new_n666), .C1(new_n659), .C2(new_n663), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G22), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G166), .B2(new_n674), .ZN(new_n676));
  INV_X1    g251(.A(G1971), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(G16), .A2(G23), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT82), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G288), .B2(new_n674), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT83), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT33), .B(G1976), .Z(new_n683));
  OAI21_X1  g258(.A(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(G6), .B(G305), .S(G16), .Z(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT32), .B(G1981), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI211_X1 g264(.A(new_n684), .B(new_n689), .C1(new_n686), .C2(new_n685), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT84), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(KEYINPUT34), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n690), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT34), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(G16), .A2(G24), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n578), .B(KEYINPUT81), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1986), .ZN(new_n700));
  OR2_X1    g275(.A1(G95), .A2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n701), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT80), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n480), .B2(G119), .ZN(new_n704));
  INV_X1    g279(.A(G131), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n473), .ZN(new_n706));
  MUX2_X1   g281(.A(G25), .B(new_n706), .S(G29), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n711));
  AOI211_X1 g286(.A(new_n700), .B(new_n710), .C1(new_n711), .C2(KEYINPUT36), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n692), .A2(new_n696), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(KEYINPUT36), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G32), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n474), .A2(G141), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT89), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT26), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n467), .A2(G105), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n722), .B(new_n723), .C1(new_n480), .C2(G129), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n718), .B1(new_n726), .B2(new_n717), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT27), .B(G1996), .Z(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT90), .Z(new_n730));
  NAND3_X1  g305(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT25), .Z(new_n732));
  AOI22_X1  g307(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n465), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n474), .B2(G139), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT87), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(new_n717), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n717), .B2(G33), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n738), .A2(new_n442), .B1(new_n727), .B2(new_n728), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n442), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n674), .A2(G5), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G171), .B2(new_n674), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(G1961), .ZN(new_n743));
  AND2_X1   g318(.A1(KEYINPUT24), .A2(G34), .ZN(new_n744));
  NOR2_X1   g319(.A1(KEYINPUT24), .A2(G34), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n717), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT88), .Z(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n470), .B2(new_n717), .ZN(new_n748));
  INV_X1    g323(.A(G2084), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n717), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n717), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2078), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n743), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  AND3_X1   g329(.A1(new_n739), .A2(new_n740), .A3(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n616), .A2(new_n717), .ZN(new_n756));
  OR2_X1    g331(.A1(KEYINPUT30), .A2(G28), .ZN(new_n757));
  NAND2_X1  g332(.A1(KEYINPUT30), .A2(G28), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT31), .B(G11), .Z(new_n760));
  AOI211_X1 g335(.A(new_n759), .B(new_n760), .C1(new_n742), .C2(G1961), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n674), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n674), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT91), .B(G1966), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n763), .A2(new_n765), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n756), .A2(new_n761), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(KEYINPUT92), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(KEYINPUT92), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n730), .A2(new_n755), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT93), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n717), .A2(G35), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n482), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT29), .ZN(new_n775));
  INV_X1    g350(.A(G2090), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n674), .A2(G20), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT23), .Z(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G1956), .Z(new_n781));
  OAI21_X1  g356(.A(KEYINPUT94), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  OR3_X1    g357(.A1(new_n777), .A2(KEYINPUT94), .A3(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n674), .A2(G4), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n593), .B2(new_n674), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT86), .B(G1348), .Z(new_n786));
  XOR2_X1   g361(.A(new_n785), .B(new_n786), .Z(new_n787));
  AND2_X1   g362(.A1(new_n674), .A2(G19), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n601), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1341), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n717), .A2(G26), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT28), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n474), .A2(G140), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n480), .A2(G128), .ZN(new_n795));
  OR2_X1    g370(.A1(G104), .A2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n796), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n793), .B1(new_n798), .B2(G29), .ZN(new_n799));
  INV_X1    g374(.A(G2067), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n789), .A2(new_n790), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n787), .A2(new_n791), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n775), .A2(new_n776), .ZN(new_n804));
  AND4_X1   g379(.A1(new_n782), .A2(new_n783), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n715), .A2(new_n716), .A3(new_n772), .A4(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  XOR2_X1   g382(.A(KEYINPUT96), .B(G860), .Z(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n593), .A2(G559), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT38), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n522), .A2(G67), .ZN(new_n812));
  AND2_X1   g387(.A1(G80), .A2(G543), .ZN(new_n813));
  OAI21_X1  g388(.A(G651), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT95), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n525), .A2(G93), .B1(G55), .B2(new_n519), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n601), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n601), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n811), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n809), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n824), .B2(new_n823), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n819), .A2(new_n809), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(G145));
  XNOR2_X1  g404(.A(new_n482), .B(new_n616), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n470), .B(KEYINPUT97), .Z(new_n831));
  XOR2_X1   g406(.A(new_n830), .B(new_n831), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n474), .A2(G142), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT99), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n480), .A2(G130), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n465), .A2(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n706), .B(new_n620), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n464), .A2(new_n484), .B1(new_n843), .B2(new_n491), .ZN(new_n844));
  INV_X1    g419(.A(new_n499), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n498), .B1(new_n464), .B2(new_n495), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n736), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n726), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n725), .A2(new_n848), .A3(new_n736), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n798), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n798), .B1(new_n850), .B2(new_n851), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n847), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(G164), .A3(new_n852), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n841), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n857), .A3(new_n841), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI211_X1 g436(.A(KEYINPUT100), .B(new_n841), .C1(new_n855), .C2(new_n857), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n832), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n858), .A2(new_n832), .ZN(new_n864));
  AOI21_X1  g439(.A(G37), .B1(new_n864), .B2(new_n860), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n863), .A2(KEYINPUT40), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT40), .B1(new_n863), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(G395));
  NAND2_X1  g443(.A1(new_n819), .A2(new_n580), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n604), .A2(new_n822), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n589), .A2(new_n549), .A3(new_n553), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT102), .ZN(new_n872));
  NAND3_X1  g447(.A1(G299), .A2(new_n588), .A3(new_n584), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n873), .A2(KEYINPUT41), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n871), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n602), .A2(new_n603), .A3(new_n821), .A4(new_n820), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n870), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT103), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n870), .A2(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n871), .A2(new_n873), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT101), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n870), .A2(new_n879), .A3(new_n889), .A4(new_n880), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n882), .A2(new_n883), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(G290), .B(G305), .ZN(new_n892));
  XNOR2_X1  g467(.A(G303), .B(G288), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n892), .B(new_n893), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT42), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n882), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n888), .A2(new_n890), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT104), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g475(.A(KEYINPUT104), .B(new_n895), .C1(new_n897), .C2(new_n898), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n869), .B1(new_n902), .B2(new_n580), .ZN(G295));
  OAI21_X1  g478(.A(new_n869), .B1(new_n902), .B2(new_n580), .ZN(G331));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  INV_X1    g481(.A(new_n894), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n908));
  NAND2_X1  g483(.A1(G301), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(G171), .A2(KEYINPUT105), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(G168), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(G286), .A2(new_n908), .A3(G301), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n822), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n820), .A2(new_n821), .A3(new_n912), .A4(new_n911), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n885), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT106), .B1(new_n914), .B2(new_n915), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n822), .B2(new_n913), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n874), .A2(new_n875), .B1(new_n871), .B2(new_n877), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n907), .B(new_n916), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n879), .B1(new_n917), .B2(new_n919), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n907), .B1(new_n925), .B2(new_n916), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n906), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n917), .A2(new_n886), .A3(new_n919), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n872), .A2(new_n877), .B1(new_n875), .B2(new_n885), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n914), .B2(new_n915), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n894), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n931), .A2(new_n922), .A3(KEYINPUT43), .A4(new_n923), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n905), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n924), .B2(new_n926), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n931), .A2(new_n922), .A3(new_n906), .A4(new_n923), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n905), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT44), .B1(new_n935), .B2(new_n936), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT107), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(G397));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(G164), .B2(G1384), .ZN(new_n945));
  OAI211_X1 g520(.A(G40), .B(new_n468), .C1(new_n469), .C2(new_n465), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1996), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT46), .Z(new_n950));
  XNOR2_X1  g525(.A(new_n798), .B(new_n800), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n952), .B2(new_n947), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n953), .B(KEYINPUT47), .Z(new_n954));
  INV_X1    g529(.A(new_n947), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n725), .B(new_n948), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n956), .A2(new_n951), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n706), .B(new_n708), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR4_X1   g534(.A1(G290), .A2(new_n945), .A3(G1986), .A4(new_n946), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT48), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n798), .A2(G2067), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n706), .A2(new_n709), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n957), .B2(new_n963), .ZN(new_n964));
  OAI221_X1 g539(.A(new_n954), .B1(new_n959), .B2(new_n961), .C1(new_n964), .C2(new_n955), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n965), .B(KEYINPUT127), .Z(new_n966));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(G164), .B2(G1384), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n847), .A2(KEYINPUT109), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n847), .A2(new_n970), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n946), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1961), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n847), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n978));
  INV_X1    g553(.A(new_n946), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n945), .A2(new_n978), .A3(new_n443), .A4(new_n979), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n975), .A2(new_n976), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n978), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n847), .A2(KEYINPUT114), .A3(KEYINPUT45), .A4(new_n970), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(G164), .A2(new_n967), .A3(G1384), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT109), .B1(new_n847), .B2(new_n970), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n944), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n977), .A2(G2078), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n985), .A2(new_n988), .A3(new_n979), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(G301), .B1(new_n981), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n972), .A2(new_n776), .A3(new_n974), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n945), .A2(new_n979), .A3(new_n978), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n677), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G166), .B2(new_n992), .ZN(new_n998));
  OAI211_X1 g573(.A(KEYINPUT55), .B(G8), .C1(new_n510), .C2(new_n514), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n998), .A2(KEYINPUT110), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT110), .B1(new_n998), .B2(new_n999), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n996), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT111), .B(G8), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n969), .B1(new_n968), .B2(new_n971), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n979), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1008), .A3(new_n776), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1004), .B1(new_n1009), .B2(new_n995), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n998), .A2(new_n999), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1003), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT112), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1015), .B(new_n565), .C1(new_n570), .C2(new_n571), .ZN(new_n1016));
  OAI21_X1  g591(.A(G1981), .B1(new_n564), .B2(new_n568), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1004), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n968), .A2(new_n979), .A3(new_n971), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1016), .A2(new_n1017), .A3(new_n1014), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G288), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(G1976), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(G288), .B2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1021), .A2(new_n1025), .A3(new_n1027), .A4(new_n1020), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1021), .A2(new_n1025), .A3(new_n1020), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT52), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1023), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1012), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n985), .A2(new_n988), .A3(new_n979), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n764), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n972), .A2(new_n974), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n749), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(KEYINPUT123), .A3(new_n1020), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT123), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1033), .A2(new_n764), .B1(new_n1035), .B2(new_n749), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(new_n1004), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G168), .A2(new_n1004), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(KEYINPUT51), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1040), .A2(new_n992), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT51), .B1(new_n1045), .B2(new_n1042), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1044), .A2(new_n1046), .B1(new_n1042), .B2(new_n1037), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT62), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n991), .B(new_n1032), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n975), .A2(new_n976), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n980), .A2(new_n977), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n990), .A2(new_n1051), .A3(G301), .A4(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n980), .A2(new_n977), .ZN(new_n1054));
  AOI21_X1  g629(.A(G1961), .B1(new_n972), .B2(new_n974), .ZN(new_n1055));
  INV_X1    g630(.A(new_n989), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n994), .A2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1053), .B(KEYINPUT54), .C1(new_n1058), .C2(G301), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1031), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1005), .A2(G2090), .A3(new_n1007), .ZN(new_n1061));
  INV_X1    g636(.A(new_n995), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1020), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1011), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1063), .A2(new_n1064), .B1(new_n996), .B2(new_n1002), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1059), .A2(new_n1060), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n990), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G171), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1057), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n981), .A2(G301), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1067), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI211_X1 g649(.A(KEYINPUT124), .B(KEYINPUT54), .C1(new_n1069), .C2(new_n1071), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1066), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT125), .B1(new_n1076), .B2(new_n1047), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1037), .A2(new_n1042), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1059), .A2(new_n1060), .A3(new_n1065), .ZN(new_n1081));
  NOR4_X1   g656(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .A4(G171), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1073), .B1(new_n1082), .B2(new_n991), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT124), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1072), .A2(new_n1067), .A3(new_n1073), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1081), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1080), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n1089));
  XNOR2_X1  g664(.A(G299), .B(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1091), .B(KEYINPUT118), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n945), .A2(new_n978), .A3(new_n979), .A4(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(G1956), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1090), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1096), .B2(new_n1095), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1021), .A2(G2067), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n786), .B2(new_n975), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(new_n589), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1090), .B(new_n1093), .C1(G1956), .C2(new_n1094), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(G299), .B(KEYINPUT57), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1095), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT61), .B1(new_n1106), .B2(new_n1102), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT122), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1102), .A2(KEYINPUT61), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1098), .A2(new_n1109), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n589), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n589), .B1(new_n1100), .B2(KEYINPUT60), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1111), .A2(new_n1112), .B1(KEYINPUT60), .B2(new_n1100), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n945), .A2(new_n978), .A3(new_n948), .A4(new_n979), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  AOI22_X1  g690(.A1(KEYINPUT120), .A2(new_n1114), .B1(new_n1021), .B2(new_n1115), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1114), .A2(KEYINPUT120), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n601), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(KEYINPUT121), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1122));
  NOR2_X1   g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1110), .A2(new_n1113), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1104), .B1(new_n1108), .B2(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1077), .A2(new_n1088), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1030), .A2(new_n1028), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1022), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(new_n1018), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT113), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT113), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1023), .A2(new_n1132), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1003), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1021), .A2(new_n1020), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1023), .A2(new_n1026), .A3(new_n1024), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(new_n1136), .B2(new_n1016), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n968), .A2(new_n971), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n946), .B1(new_n1139), .B2(new_n944), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n765), .B1(new_n1140), .B2(new_n985), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n975), .A2(G2084), .ZN(new_n1142));
  OAI211_X1 g717(.A(G168), .B(new_n1020), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1037), .A2(KEYINPUT115), .A3(G168), .A4(new_n1020), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1003), .A2(KEYINPUT63), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n996), .A2(new_n1011), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1149), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1147), .B(new_n1148), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT63), .B1(new_n1032), .B2(new_n1147), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT116), .ZN(new_n1156));
  OAI22_X1  g731(.A1(new_n1152), .A2(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1138), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT126), .B1(new_n1127), .B2(new_n1159), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1077), .A2(new_n1126), .A3(new_n1088), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1138), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1050), .B1(new_n1160), .B2(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n578), .B(G1986), .Z(new_n1169));
  AOI21_X1  g744(.A(new_n959), .B1(new_n947), .B2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT108), .Z(new_n1171));
  OAI21_X1  g746(.A(new_n966), .B1(new_n1168), .B2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g747(.A1(new_n863), .A2(new_n865), .ZN(new_n1174));
  NOR4_X1   g748(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n1174), .A2(new_n1175), .A3(new_n937), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


