//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AND2_X1   g0009(.A1(G68), .A2(G238), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G97), .A2(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n210), .B(new_n214), .C1(G107), .C2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G116), .A2(G270), .ZN(new_n216));
  AND2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(G58), .A2(G232), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n204), .ZN(new_n227));
  NOR2_X1   g0027(.A1(G58), .A2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n209), .B(new_n225), .C1(new_n227), .C2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n239), .B(G270), .Z(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NOR2_X1   g0048(.A1(KEYINPUT8), .A2(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT66), .B(G58), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n249), .B1(new_n250), .B2(KEYINPUT8), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n251), .A2(new_n253), .B1(G150), .B2(new_n254), .ZN(new_n255));
  OR2_X1    g0055(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n256));
  OAI21_X1  g0056(.A(G20), .B1(new_n229), .B2(G50), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n226), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n260), .B1(new_n205), .B2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n203), .A2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G50), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n261), .A2(new_n264), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n218), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n263), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT65), .B1(new_n276), .B2(new_n226), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT65), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n260), .A2(new_n278), .A3(new_n275), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n274), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n277), .B2(new_n279), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G226), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT3), .B(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G222), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G223), .A2(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n276), .A2(new_n226), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n291), .B(new_n292), .C1(G77), .C2(new_n287), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n284), .A2(new_n286), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G179), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n294), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n273), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n287), .A2(G232), .A3(new_n288), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT68), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G107), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n287), .A2(G238), .A3(G1698), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n287), .A2(KEYINPUT68), .A3(G232), .A4(new_n288), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n301), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n292), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n285), .A2(G244), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n284), .A3(new_n311), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n312), .A2(G179), .ZN(new_n313));
  XOR2_X1   g0113(.A(KEYINPUT15), .B(G87), .Z(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n253), .ZN(new_n315));
  INV_X1    g0115(.A(new_n254), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT8), .B(G58), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n315), .B1(new_n204), .B2(new_n220), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(new_n262), .B1(new_n220), .B2(new_n266), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n261), .A2(G77), .A3(new_n264), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n312), .A2(new_n296), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n313), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n321), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n312), .A2(G200), .ZN(new_n325));
  INV_X1    g0125(.A(G190), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n324), .B(new_n325), .C1(new_n326), .C2(new_n312), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n263), .A2(KEYINPUT9), .A3(new_n269), .A4(new_n272), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n294), .A2(new_n326), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT10), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n268), .B1(new_n259), .B2(new_n262), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT9), .B1(new_n333), .B2(new_n272), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n294), .A2(G200), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n331), .A2(new_n332), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n329), .A2(new_n336), .A3(new_n330), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT10), .B1(new_n338), .B2(new_n334), .ZN(new_n339));
  AOI211_X1 g0139(.A(new_n298), .B(new_n328), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT14), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n285), .A2(G238), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n219), .A2(new_n288), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(G232), .B2(new_n288), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n343), .B1(new_n345), .B2(new_n305), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n292), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n284), .A2(new_n342), .A3(new_n347), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n348), .A2(KEYINPUT13), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(KEYINPUT13), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n341), .B1(new_n351), .B2(G169), .ZN(new_n352));
  AOI211_X1 g0152(.A(KEYINPUT14), .B(new_n296), .C1(new_n349), .C2(new_n350), .ZN(new_n353));
  INV_X1    g0153(.A(G179), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n253), .A2(G77), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n358), .B1(new_n204), .B2(G68), .C1(new_n316), .C2(new_n218), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n262), .ZN(new_n360));
  XOR2_X1   g0160(.A(new_n360), .B(KEYINPUT11), .Z(new_n361));
  INV_X1    g0161(.A(G68), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n270), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n266), .A2(new_n362), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT12), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n361), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n357), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n351), .A2(G200), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n367), .B(new_n370), .C1(new_n326), .C2(new_n351), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n228), .B1(new_n250), .B2(G68), .ZN(new_n374));
  INV_X1    g0174(.A(G159), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n374), .A2(new_n204), .B1(new_n375), .B2(new_n316), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n287), .B2(G20), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n302), .A2(G33), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT7), .B(new_n204), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n362), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n373), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT70), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT69), .B1(new_n302), .B2(G33), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT69), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(new_n252), .A3(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n303), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(new_n377), .A3(new_n204), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n379), .B1(new_n385), .B2(new_n387), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT7), .B1(new_n391), .B2(G20), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(G68), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n376), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT70), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n396), .B(new_n373), .C1(new_n376), .C2(new_n382), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n384), .A2(new_n262), .A3(new_n395), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n285), .A2(G232), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n284), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT72), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n288), .A2(G223), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n401), .B1(new_n389), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n219), .A2(new_n288), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n391), .A2(new_n404), .B1(G33), .B2(G87), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n391), .A2(KEYINPUT72), .A3(G223), .A4(new_n288), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n400), .B1(new_n407), .B2(new_n292), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G190), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n270), .A2(new_n251), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n251), .B2(new_n266), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n398), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n407), .A2(new_n292), .ZN(new_n413));
  INV_X1    g0213(.A(new_n400), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G200), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n412), .A2(KEYINPUT73), .A3(KEYINPUT17), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n416), .A2(new_n398), .A3(new_n409), .A4(new_n411), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT73), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n413), .A2(G179), .A3(new_n414), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n296), .B2(new_n408), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT71), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n398), .A2(new_n425), .A3(new_n411), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n398), .B2(new_n411), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(KEYINPUT18), .B(new_n424), .C1(new_n426), .C2(new_n427), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n422), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n340), .A2(new_n372), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT74), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n340), .A2(new_n372), .A3(KEYINPUT74), .A4(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n287), .A2(new_n204), .A3(G87), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT22), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT23), .B1(new_n204), .B2(G107), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT83), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n204), .A2(KEYINPUT23), .A3(G107), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n444), .B1(KEYINPUT82), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n440), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n391), .A2(KEYINPUT22), .A3(new_n204), .A4(G87), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n445), .A2(KEYINPUT82), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n447), .A2(KEYINPUT24), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT24), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n440), .A2(new_n443), .A3(new_n449), .A4(new_n446), .ZN(new_n452));
  INV_X1    g0252(.A(new_n448), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(new_n454), .A3(new_n262), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n252), .A2(G1), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n262), .A2(new_n266), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G107), .ZN(new_n458));
  INV_X1    g0258(.A(G107), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n266), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g0260(.A(new_n460), .B(KEYINPUT25), .Z(new_n461));
  NAND3_X1  g0261(.A1(new_n455), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n281), .A2(KEYINPUT5), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n203), .A2(G45), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT78), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n281), .A2(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G41), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT78), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n203), .A4(G45), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n465), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n277), .A2(new_n279), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(KEYINPUT85), .A3(G264), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(G264), .A3(new_n472), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT85), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n391), .B1(G257), .B2(new_n288), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G250), .A2(G1698), .ZN(new_n479));
  INV_X1    g0279(.A(G294), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n478), .A2(new_n479), .B1(new_n252), .B2(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n474), .A2(new_n477), .B1(new_n292), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n472), .A2(G274), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT79), .B1(new_n483), .B2(new_n471), .ZN(new_n484));
  INV_X1    g0284(.A(new_n471), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT79), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(new_n280), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G200), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n481), .A2(new_n292), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n492), .A3(new_n475), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n493), .A2(G190), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n462), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n462), .A2(KEYINPUT84), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT84), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n455), .A2(new_n497), .A3(new_n458), .A4(new_n461), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n493), .A2(G169), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n489), .B2(new_n354), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n495), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n305), .A2(G303), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n391), .B1(G264), .B2(new_n288), .ZN(new_n504));
  NOR2_X1   g0304(.A1(G257), .A2(G1698), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n292), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n473), .A2(G270), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n488), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G200), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n326), .B2(new_n509), .ZN(new_n511));
  INV_X1    g0311(.A(G116), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n266), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n457), .A2(G116), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(G20), .ZN(new_n515));
  AOI21_X1  g0315(.A(G20), .B1(G33), .B2(G283), .ZN(new_n516));
  INV_X1    g0316(.A(G97), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(G33), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n262), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT20), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n513), .B(new_n514), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n511), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n523), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n488), .A2(new_n507), .A3(G179), .A4(new_n508), .ZN(new_n526));
  OR2_X1    g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n509), .A2(new_n523), .A3(G169), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT21), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n509), .A2(new_n523), .A3(KEYINPUT21), .A4(G169), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n464), .A2(new_n213), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n203), .A2(new_n274), .A3(G45), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n472), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G238), .A2(G1698), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n221), .B2(G1698), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n391), .A2(new_n538), .B1(G33), .B2(G116), .ZN(new_n539));
  INV_X1    g0339(.A(new_n292), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G190), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n391), .A2(new_n204), .A3(G68), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n204), .B1(new_n343), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G97), .A2(G107), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n212), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n204), .A2(G33), .A3(G97), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n546), .A2(new_n548), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n314), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n551), .A2(new_n262), .B1(new_n266), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n541), .A2(G200), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n457), .A2(G87), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n543), .A2(new_n553), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n541), .A2(G169), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n536), .B(G179), .C1(new_n539), .C2(new_n540), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n457), .A2(new_n314), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n553), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT81), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n221), .A2(G1698), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n391), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g0367(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n305), .A2(new_n288), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n287), .A2(KEYINPUT4), .A3(new_n566), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT77), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n287), .A2(KEYINPUT77), .A3(KEYINPUT4), .A4(new_n566), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n569), .A2(new_n571), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n292), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n473), .A2(G257), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n577), .A2(G190), .A3(new_n488), .A4(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT80), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n577), .A2(new_n488), .A3(new_n578), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G200), .ZN(new_n583));
  XNOR2_X1  g0383(.A(G97), .B(G107), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT6), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n585), .B2(new_n459), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n587), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(G20), .B1(G77), .B2(new_n254), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n378), .A2(new_n381), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G107), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n261), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n457), .A2(G97), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n267), .A2(G97), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n576), .A2(new_n292), .B1(new_n484), .B2(new_n487), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n598), .A2(KEYINPUT80), .A3(G190), .A4(new_n578), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n581), .A2(new_n583), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n597), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n582), .A2(new_n296), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(new_n354), .A3(new_n578), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n556), .A2(KEYINPUT81), .A3(new_n562), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n565), .A2(new_n600), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n437), .A2(new_n502), .A3(new_n533), .A4(new_n606), .ZN(G372));
  NAND2_X1  g0407(.A1(new_n565), .A2(new_n605), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT26), .B1(new_n608), .B2(new_n604), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT86), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n559), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n557), .A2(KEYINPUT86), .A3(new_n558), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n561), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n553), .A2(new_n555), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(G200), .B2(new_n541), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n613), .A2(new_n561), .B1(new_n616), .B2(new_n543), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n609), .B(new_n614), .C1(KEYINPUT26), .C2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n501), .A2(new_n462), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(new_n532), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n455), .A2(new_n458), .A3(new_n461), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n493), .A2(G190), .ZN(new_n624));
  AOI21_X1  g0424(.A(G200), .B1(new_n482), .B2(new_n488), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n626), .A2(new_n617), .A3(new_n604), .A4(new_n600), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n620), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n437), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n298), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n337), .A2(new_n339), .ZN(new_n632));
  INV_X1    g0432(.A(new_n323), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n357), .A2(new_n368), .B1(new_n633), .B2(new_n371), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(new_n422), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n398), .A2(new_n411), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n424), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n637), .B(KEYINPUT18), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n632), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n630), .A2(new_n631), .A3(new_n639), .ZN(G369));
  NOR2_X1   g0440(.A1(new_n265), .A2(G20), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n203), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n523), .A2(new_n647), .ZN(new_n648));
  MUX2_X1   g0448(.A(new_n532), .B(new_n533), .S(new_n648), .Z(new_n649));
  NAND2_X1  g0449(.A1(new_n499), .A2(new_n647), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n502), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n499), .A2(new_n501), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n647), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n649), .A2(new_n654), .A3(G330), .ZN(new_n655));
  INV_X1    g0455(.A(new_n647), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n532), .A2(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n502), .A2(new_n657), .B1(new_n621), .B2(new_n656), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n658), .ZN(G399));
  INV_X1    g0459(.A(new_n207), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(G41), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n548), .A2(G116), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G1), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n230), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n619), .A2(KEYINPUT26), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n532), .B1(new_n499), .B2(new_n501), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n667), .B(new_n614), .C1(new_n668), .C2(new_n627), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n608), .A2(KEYINPUT26), .A3(new_n604), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(KEYINPUT88), .A3(KEYINPUT29), .A4(new_n656), .ZN(new_n672));
  OAI211_X1 g0472(.A(KEYINPUT29), .B(new_n656), .C1(new_n669), .C2(new_n670), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT88), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n656), .B1(new_n620), .B2(new_n628), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT29), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n672), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n606), .A2(new_n502), .A3(new_n533), .A4(new_n656), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n526), .A2(KEYINPUT87), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n484), .A2(new_n487), .B1(G270), .B2(new_n473), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT87), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(G179), .A4(new_n507), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n482), .A2(new_n598), .A3(new_n578), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n542), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n685), .A2(KEYINPUT30), .A3(new_n686), .A4(new_n542), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n542), .B1(new_n598), .B2(new_n578), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n354), .A3(new_n489), .A4(new_n509), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n647), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n680), .A2(new_n694), .A3(KEYINPUT31), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT31), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(new_n696), .A3(new_n647), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n679), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n666), .B1(new_n701), .B2(G1), .ZN(G364));
  OR2_X1    g0502(.A1(new_n649), .A2(G330), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT89), .B1(new_n649), .B2(G330), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n641), .A2(G45), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n662), .A2(G1), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(G13), .A2(G33), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G20), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n226), .B1(G20), .B2(new_n296), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n660), .A2(new_n391), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n282), .B2(new_n231), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n244), .A2(G45), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(new_n512), .B2(new_n660), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n207), .A2(G355), .A3(new_n287), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n714), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n490), .A2(G179), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n204), .A2(G190), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n459), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n354), .A2(new_n490), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n723), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G179), .A2(G200), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n204), .B1(new_n728), .B2(G190), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n727), .A2(new_n362), .B1(new_n729), .B2(new_n517), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT92), .Z(new_n731));
  NOR2_X1   g0531(.A1(new_n204), .A2(new_n326), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n726), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n725), .B(new_n731), .C1(G50), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n732), .A2(new_n722), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G87), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n354), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n732), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n723), .A2(new_n739), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n745), .A2(new_n250), .B1(G77), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n723), .A2(new_n728), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  XOR2_X1   g0550(.A(KEYINPUT91), .B(G159), .Z(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT32), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n305), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n735), .A2(new_n738), .A3(new_n748), .A4(new_n754), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT93), .B(G317), .Z(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT33), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n727), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G311), .A2(new_n747), .B1(new_n750), .B2(G329), .ZN(new_n759));
  INV_X1    g0559(.A(G283), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n759), .B1(new_n760), .B2(new_n724), .C1(new_n480), .C2(new_n729), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n758), .B(new_n761), .C1(G322), .C2(new_n745), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n734), .A2(G326), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n737), .A2(G303), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n762), .A2(new_n305), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n755), .A2(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n707), .B(new_n721), .C1(new_n766), .C2(new_n712), .ZN(new_n767));
  INV_X1    g0567(.A(new_n711), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n649), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n708), .A2(new_n769), .ZN(G396));
  NAND2_X1  g0570(.A1(new_n321), .A2(new_n647), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n323), .A2(new_n327), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT94), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n323), .A2(new_n327), .A3(KEYINPUT94), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n656), .B(new_n777), .C1(new_n620), .C2(new_n628), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n633), .A2(new_n647), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT95), .Z(new_n781));
  INV_X1    g0581(.A(new_n676), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n778), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(new_n699), .Z(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n707), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n736), .A2(new_n218), .ZN(new_n786));
  INV_X1    g0586(.A(new_n727), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G137), .A2(new_n734), .B1(new_n787), .B2(G150), .ZN(new_n788));
  INV_X1    g0588(.A(new_n751), .ZN(new_n789));
  INV_X1    g0589(.A(G143), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n788), .B1(new_n746), .B2(new_n789), .C1(new_n744), .C2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT34), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n389), .B1(G132), .B2(new_n750), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n792), .B(new_n793), .C1(new_n362), .C2(new_n724), .ZN(new_n794));
  INV_X1    g0594(.A(new_n729), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n786), .B(new_n794), .C1(new_n250), .C2(new_n795), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n305), .B1(new_n746), .B2(new_n512), .C1(new_n459), .C2(new_n736), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n745), .A2(G294), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n734), .A2(G303), .ZN(new_n799));
  INV_X1    g0599(.A(new_n724), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G87), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G311), .A2(new_n750), .B1(new_n795), .B2(G97), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n798), .A2(new_n799), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n797), .B(new_n803), .C1(G283), .C2(new_n787), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n712), .B1(new_n796), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n707), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n712), .A2(new_n709), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n220), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n776), .A2(new_n709), .A3(new_n779), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n805), .A2(new_n806), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n785), .A2(new_n810), .ZN(G384));
  INV_X1    g0611(.A(new_n645), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n426), .A2(new_n427), .B1(new_n424), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT37), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n419), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT96), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n395), .A2(new_n262), .ZN(new_n818));
  AOI21_X1  g0618(.A(KEYINPUT16), .B1(new_n393), .B2(new_n394), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n411), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n424), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n812), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n821), .A2(new_n419), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT37), .ZN(new_n824));
  AND3_X1   g0624(.A1(new_n816), .A2(new_n817), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n817), .B1(new_n816), .B2(new_n824), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n430), .A2(new_n431), .ZN(new_n828));
  INV_X1    g0628(.A(new_n422), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n822), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT38), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n822), .B1(new_n828), .B2(new_n829), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n834), .A2(new_n825), .A3(new_n826), .A4(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT97), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n826), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n816), .A2(new_n817), .A3(new_n824), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n835), .B1(new_n840), .B2(new_n834), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n827), .A2(new_n832), .A3(KEYINPUT38), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT97), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n357), .A2(new_n368), .A3(new_n647), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n368), .A2(new_n647), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n371), .B(new_n846), .C1(new_n356), .C2(new_n367), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n845), .A2(new_n847), .B1(new_n776), .B2(new_n779), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n695), .A2(new_n697), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n837), .A2(new_n844), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT40), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT98), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n637), .A2(new_n419), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n812), .B1(new_n426), .B2(new_n427), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n814), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n813), .A2(new_n815), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n427), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n398), .A2(new_n425), .A3(new_n411), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n645), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n638), .B2(new_n422), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n863), .B2(new_n855), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(KEYINPUT98), .A3(new_n816), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n860), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n835), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n852), .B(new_n849), .C1(new_n842), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n853), .A2(G330), .A3(new_n870), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n437), .A2(G330), .A3(new_n698), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n869), .B1(new_n851), .B2(new_n852), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n437), .A2(new_n698), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n871), .A2(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n639), .A2(new_n631), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n672), .A2(new_n675), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT99), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(new_n437), .A4(new_n678), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n435), .A2(new_n436), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT99), .B1(new_n679), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n877), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n876), .B(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT39), .B1(new_n868), .B2(new_n842), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n369), .A2(new_n647), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT39), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n638), .A2(new_n645), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n845), .A2(new_n847), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n323), .A2(new_n647), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(new_n778), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n837), .A2(new_n844), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n889), .A2(new_n890), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n884), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n203), .B2(new_n641), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n512), .B1(new_n590), .B2(KEYINPUT35), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n227), .C1(KEYINPUT35), .C2(new_n590), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT36), .ZN(new_n903));
  INV_X1    g0703(.A(new_n250), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n231), .B(G77), .C1(new_n362), .C2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(G50), .B2(new_n362), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(G1), .A3(new_n265), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n900), .A2(new_n903), .A3(new_n907), .ZN(G367));
  AND2_X1   g0708(.A1(new_n600), .A2(new_n604), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n597), .B2(new_n656), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n618), .A2(new_n647), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT102), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT102), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n910), .A2(new_n914), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n655), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n615), .A2(new_n647), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n614), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n617), .A2(new_n920), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n913), .A2(new_n652), .A3(new_n915), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n647), .B1(new_n925), .B2(new_n604), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n502), .A2(new_n657), .A3(new_n909), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT42), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n924), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT101), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT101), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(new_n924), .C1(new_n926), .C2(new_n928), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n919), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n923), .ZN(new_n935));
  XNOR2_X1  g0735(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n930), .A2(new_n919), .A3(new_n932), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n934), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n930), .A2(new_n919), .A3(new_n932), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n937), .B1(new_n941), .B2(new_n933), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n661), .B(KEYINPUT41), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n502), .A2(new_n657), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n654), .B2(new_n657), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n649), .A2(G330), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT104), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT104), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n949), .A2(new_n655), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n700), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT105), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT105), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n700), .B2(new_n952), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT103), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n912), .A2(new_n957), .A3(new_n658), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n957), .B1(new_n912), .B2(new_n658), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT45), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n912), .A2(new_n658), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT44), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n960), .B1(new_n958), .B2(new_n959), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n961), .A2(new_n963), .A3(new_n655), .A4(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n918), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n954), .A2(new_n956), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n944), .B1(new_n968), .B2(new_n701), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n706), .A2(G1), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n940), .B(new_n942), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n787), .A2(G294), .B1(new_n795), .B2(G107), .ZN(new_n972));
  INV_X1    g0772(.A(G311), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n972), .B1(new_n973), .B2(new_n733), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n724), .A2(new_n517), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n746), .A2(new_n760), .ZN(new_n976));
  NOR4_X1   g0776(.A1(new_n974), .A2(new_n391), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT106), .B1(new_n737), .B2(G116), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT46), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n745), .A2(G303), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n750), .A2(G317), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n977), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT107), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n724), .A2(new_n220), .ZN(new_n984));
  XOR2_X1   g0784(.A(KEYINPUT109), .B(G137), .Z(new_n985));
  AOI21_X1  g0785(.A(new_n305), .B1(new_n750), .B2(new_n985), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n218), .B2(new_n746), .C1(new_n790), .C2(new_n733), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n984), .B(new_n987), .C1(new_n787), .C2(new_n751), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n904), .B2(new_n736), .ZN(new_n989));
  INV_X1    g0789(.A(G150), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n744), .A2(new_n990), .B1(new_n362), .B2(new_n729), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT108), .Z(new_n992));
  OAI21_X1  g0792(.A(new_n983), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n712), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n935), .A2(new_n711), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n713), .B1(new_n207), .B2(new_n552), .C1(new_n240), .C2(new_n716), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n995), .A2(new_n806), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n971), .A2(new_n998), .ZN(G387));
  XOR2_X1   g0799(.A(new_n661), .B(KEYINPUT113), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n953), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n952), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1001), .B1(new_n701), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n651), .A2(new_n653), .A3(new_n711), .ZN(new_n1004));
  OR3_X1    g0804(.A1(new_n317), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT50), .B1(new_n317), .B2(G50), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1005), .A2(new_n282), .A3(new_n663), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n362), .A2(new_n220), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n715), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT111), .Z(new_n1010));
  INV_X1    g0810(.A(new_n237), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1010), .B1(new_n282), .B2(new_n1011), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n660), .A2(new_n663), .A3(new_n305), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n459), .B2(new_n660), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT110), .Z(new_n1015));
  AOI21_X1  g0815(.A(new_n714), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n734), .A2(G159), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT112), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n389), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n1018), .B2(new_n1017), .C1(new_n362), .C2(new_n746), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n736), .A2(new_n220), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n552), .A2(new_n729), .ZN(new_n1022));
  OR4_X1    g0822(.A1(new_n975), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G150), .B2(new_n750), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n251), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1024), .B1(new_n218), .B2(new_n744), .C1(new_n1025), .C2(new_n727), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G311), .A2(new_n787), .B1(new_n747), .B2(G303), .ZN(new_n1027));
  INV_X1    g0827(.A(G322), .ZN(new_n1028));
  INV_X1    g0828(.A(G317), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n733), .C1(new_n744), .C2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT48), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n760), .B2(new_n729), .C1(new_n480), .C2(new_n736), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n750), .A2(G326), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n800), .A2(G116), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1034), .A2(new_n389), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1026), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n707), .B(new_n1016), .C1(new_n1039), .C2(new_n712), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1002), .A2(new_n970), .B1(new_n1004), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1003), .A2(new_n1041), .ZN(G393));
  INV_X1    g0842(.A(new_n1000), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT114), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n967), .A2(new_n1044), .A3(new_n965), .ZN(new_n1045));
  OR3_X1    g0845(.A1(new_n966), .A2(new_n1044), .A3(new_n918), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n968), .B(new_n1043), .C1(new_n1047), .C2(new_n953), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n970), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n744), .A2(new_n973), .B1(new_n1029), .B2(new_n733), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT115), .Z(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT52), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n787), .A2(G303), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n736), .A2(new_n760), .B1(new_n749), .B2(new_n1028), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT116), .Z(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G294), .B2(new_n747), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n729), .A2(new_n512), .ZN(new_n1058));
  NOR4_X1   g0858(.A1(new_n1057), .A2(new_n287), .A3(new_n725), .A4(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n744), .A2(new_n375), .B1(new_n990), .B2(new_n733), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n737), .A2(G68), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n787), .A2(G50), .B1(new_n795), .B2(G77), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1061), .A2(new_n801), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n746), .A2(new_n317), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n391), .B1(new_n790), .B2(new_n749), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n712), .B1(new_n1059), .B2(new_n1067), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n713), .B1(new_n517), .B2(new_n207), .C1(new_n716), .C2(new_n247), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n806), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT117), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1070), .A2(new_n1071), .B1(new_n711), .B2(new_n916), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n1071), .B2(new_n1070), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1048), .A2(new_n1049), .A3(new_n1073), .ZN(G390));
  NAND2_X1  g0874(.A1(new_n883), .A2(new_n873), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n778), .A2(new_n894), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n698), .A2(G330), .A3(new_n780), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1077), .A2(new_n892), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n892), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1077), .A2(new_n892), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n656), .B(new_n777), .C1(new_n669), .C2(new_n670), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n894), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n781), .A2(G330), .A3(new_n698), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n892), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1081), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1080), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1075), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n895), .A2(new_n887), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n886), .B2(new_n888), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n887), .B1(new_n1083), .B2(new_n891), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n868), .A2(new_n842), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1079), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n888), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1097), .A2(new_n885), .B1(new_n887), .B2(new_n895), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1098), .A2(new_n1081), .A3(new_n1094), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1089), .A2(new_n1101), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n877), .B(new_n872), .C1(new_n880), .C2(new_n882), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1080), .A2(new_n1087), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n1100), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1102), .A2(new_n1043), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1101), .A2(new_n970), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n709), .B1(new_n1097), .B2(new_n885), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1025), .A2(new_n807), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n738), .B1(new_n220), .B2(new_n729), .C1(new_n480), .C2(new_n749), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G116), .B2(new_n745), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n727), .A2(new_n459), .B1(new_n724), .B2(new_n362), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n287), .B(new_n1113), .C1(G97), .C2(new_n747), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1112), .B(new_n1114), .C1(new_n760), .C2(new_n733), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n737), .A2(G150), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT118), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT53), .Z(new_n1118));
  NAND2_X1  g0918(.A1(new_n745), .A2(G132), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n734), .A2(G128), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n787), .A2(new_n985), .B1(new_n750), .B2(G125), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n724), .A2(new_n218), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n287), .B1(new_n729), .B2(new_n375), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT54), .B(G143), .Z(new_n1124));
  AOI211_X1 g0924(.A(new_n1122), .B(new_n1123), .C1(new_n747), .C2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1115), .B1(new_n1118), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n712), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1109), .A2(new_n806), .A3(new_n1110), .A4(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1107), .A2(new_n1108), .A3(new_n1129), .ZN(G378));
  NAND2_X1  g0930(.A1(new_n632), .A2(new_n631), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1132));
  XOR2_X1   g0932(.A(new_n1131), .B(new_n1132), .Z(new_n1133));
  NAND2_X1  g0933(.A1(new_n273), .A2(new_n812), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1133), .B(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n874), .A2(G330), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n874), .B2(G330), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n897), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1103), .B1(new_n1100), .B2(new_n1088), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n871), .A2(new_n1135), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n874), .A2(G330), .A3(new_n1136), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n898), .A3(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1139), .A2(new_n1140), .A3(new_n1143), .A4(KEYINPUT57), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1043), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT121), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1137), .A2(new_n1138), .A3(new_n897), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n898), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1139), .A2(KEYINPUT121), .A3(new_n1143), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n1140), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1145), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1149), .A2(new_n970), .A3(new_n1150), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1136), .A2(new_n709), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n807), .A2(new_n218), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n904), .A2(new_n724), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n281), .B1(new_n744), .B2(new_n459), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(G283), .C2(new_n750), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n314), .A2(new_n747), .B1(new_n795), .B2(G68), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n517), .B2(new_n727), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n391), .B(new_n1161), .C1(G116), .C2(new_n734), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1159), .B(new_n1162), .C1(new_n220), .C2(new_n736), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT58), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n281), .B1(new_n389), .B2(new_n252), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1163), .A2(new_n1164), .B1(new_n218), .B2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT119), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n745), .A2(G128), .B1(new_n737), .B2(new_n1124), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n734), .A2(G125), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G137), .A2(new_n747), .B1(new_n795), .B2(G150), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G132), .B2(new_n787), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT59), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G33), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G41), .B1(new_n750), .B2(G124), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n724), .C2(new_n789), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1167), .B1(new_n1164), .B2(new_n1163), .C1(new_n1174), .C2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT120), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n712), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1155), .A2(new_n806), .A3(new_n1156), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1154), .A2(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1153), .A2(new_n1182), .ZN(G375));
  OAI21_X1  g0983(.A(KEYINPUT122), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT122), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1075), .A2(new_n1185), .A3(new_n1088), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1187), .A2(new_n943), .A3(new_n1105), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n892), .A2(new_n709), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n807), .A2(new_n362), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n746), .A2(new_n990), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n745), .A2(new_n985), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n736), .A2(new_n375), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1193), .B(new_n1157), .C1(new_n787), .C2(new_n1124), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n795), .A2(G50), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n389), .B1(G128), .B2(new_n750), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1192), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1191), .B(new_n1197), .C1(G132), .C2(new_n734), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n727), .A2(new_n512), .B1(new_n746), .B2(new_n459), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT123), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n745), .A2(G283), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1022), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n287), .B1(new_n750), .B2(G303), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n984), .B1(G97), .B2(new_n737), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1200), .B(new_n1205), .C1(G294), .C2(new_n734), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n712), .B1(new_n1198), .B2(new_n1206), .ZN(new_n1207));
  AND4_X1   g1007(.A1(new_n806), .A2(new_n1189), .A3(new_n1190), .A4(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1104), .B2(new_n970), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1188), .A2(new_n1209), .ZN(G381));
  NOR2_X1   g1010(.A1(G375), .A2(G378), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G381), .A2(G384), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1048), .A2(new_n1049), .A3(new_n1073), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(new_n998), .A3(new_n971), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(G396), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1003), .A2(new_n1216), .A3(new_n1041), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1211), .A2(new_n1212), .A3(new_n1215), .A4(new_n1218), .ZN(G407));
  NAND2_X1  g1019(.A1(new_n1211), .A2(new_n646), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(G407), .A2(G213), .A3(new_n1220), .ZN(G409));
  INV_X1    g1021(.A(KEYINPUT127), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT124), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1216), .B1(new_n1003), .B2(new_n1041), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1223), .B1(new_n1225), .B2(new_n1217), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1218), .A2(KEYINPUT124), .A3(new_n1224), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1213), .B1(new_n998), .B2(new_n971), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1228), .B1(new_n1215), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G387), .A2(G390), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1214), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(G378), .B1(new_n1153), .B2(new_n1182), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n646), .A2(G213), .ZN(new_n1237));
  INV_X1    g1037(.A(G378), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1149), .A2(new_n943), .A3(new_n1140), .A4(new_n1150), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1139), .A2(new_n970), .A3(new_n1143), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1238), .A2(new_n1181), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1184), .A2(new_n1186), .B1(new_n1105), .B2(KEYINPUT60), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1075), .A2(KEYINPUT60), .A3(new_n1088), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1043), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1209), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G384), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G384), .B(new_n1209), .C1(new_n1242), .C2(new_n1244), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1236), .A2(new_n1237), .A3(new_n1241), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT62), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1250), .B(new_n1251), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1236), .A2(new_n1237), .A3(new_n1241), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n646), .A2(G213), .A3(G2897), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1247), .A2(new_n1248), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1255), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1253), .B1(new_n1254), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1235), .B1(new_n1252), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT63), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1254), .A2(new_n1258), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(new_n1250), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1250), .A2(new_n1261), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT61), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1230), .A2(new_n1266), .A3(new_n1233), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(KEYINPUT125), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT125), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1230), .A2(new_n1269), .A3(new_n1266), .A4(new_n1233), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1263), .A2(new_n1265), .A3(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1222), .B1(new_n1260), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1262), .A2(new_n1250), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT63), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1275), .A2(new_n1264), .A3(new_n1268), .A4(new_n1270), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1250), .A2(KEYINPUT62), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1250), .A2(KEYINPUT62), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n1259), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1234), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1276), .A2(new_n1280), .A3(KEYINPUT127), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1273), .A2(new_n1281), .ZN(G405));
  XNOR2_X1  g1082(.A(G375), .B(new_n1238), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(new_n1234), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1249), .ZN(G402));
endmodule


