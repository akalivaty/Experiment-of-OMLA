

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592;

  NAND2_X1 U326 ( .A1(n295), .A2(n423), .ZN(n424) );
  XOR2_X1 U327 ( .A(n385), .B(n411), .Z(n294) );
  XOR2_X1 U328 ( .A(n379), .B(n378), .Z(n295) );
  INV_X1 U329 ( .A(n561), .ZN(n422) );
  AND2_X1 U330 ( .A1(n572), .A2(n422), .ZN(n423) );
  INV_X1 U331 ( .A(KEYINPUT33), .ZN(n350) );
  XNOR2_X1 U332 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U333 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U334 ( .A(n357), .B(n356), .ZN(n581) );
  NOR2_X1 U335 ( .A1(n526), .A2(n457), .ZN(n570) );
  XNOR2_X1 U336 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U337 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(G134GAT), .B(G43GAT), .Z(n410) );
  XOR2_X1 U339 ( .A(G120GAT), .B(G176GAT), .Z(n345) );
  XOR2_X1 U340 ( .A(n410), .B(n345), .Z(n297) );
  NAND2_X1 U341 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U343 ( .A(KEYINPUT86), .B(G71GAT), .Z(n299) );
  XNOR2_X1 U344 ( .A(KEYINPUT20), .B(KEYINPUT85), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U346 ( .A(n301), .B(n300), .Z(n305) );
  XOR2_X1 U347 ( .A(KEYINPUT0), .B(G113GAT), .Z(n436) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(KEYINPUT84), .ZN(n302) );
  XOR2_X1 U349 ( .A(G127GAT), .B(G15GAT), .Z(n389) );
  XNOR2_X1 U350 ( .A(n302), .B(n389), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n436), .B(n303), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n310) );
  XOR2_X1 U353 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n307) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G183GAT), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n309) );
  XOR2_X1 U356 ( .A(G190GAT), .B(KEYINPUT19), .Z(n308) );
  XOR2_X1 U357 ( .A(n309), .B(n308), .Z(n338) );
  XNOR2_X1 U358 ( .A(n310), .B(n338), .ZN(n535) );
  INV_X1 U359 ( .A(n535), .ZN(n526) );
  XOR2_X1 U360 ( .A(G162GAT), .B(G50GAT), .Z(n412) );
  XOR2_X1 U361 ( .A(G141GAT), .B(KEYINPUT2), .Z(n312) );
  XNOR2_X1 U362 ( .A(KEYINPUT3), .B(KEYINPUT91), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n440) );
  XOR2_X1 U364 ( .A(n412), .B(n440), .Z(n314) );
  NAND2_X1 U365 ( .A1(G228GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n327) );
  XOR2_X1 U367 ( .A(KEYINPUT22), .B(KEYINPUT94), .Z(n316) );
  XNOR2_X1 U368 ( .A(G211GAT), .B(KEYINPUT88), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U370 ( .A(KEYINPUT23), .B(KEYINPUT93), .Z(n318) );
  XNOR2_X1 U371 ( .A(KEYINPUT92), .B(KEYINPUT24), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U373 ( .A(n320), .B(n319), .Z(n325) );
  XNOR2_X1 U374 ( .A(G155GAT), .B(G22GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n321), .B(G78GAT), .ZN(n386) );
  XOR2_X1 U376 ( .A(KEYINPUT71), .B(G106GAT), .Z(n323) );
  XNOR2_X1 U377 ( .A(G148GAT), .B(G204GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n349) );
  XNOR2_X1 U379 ( .A(n386), .B(n349), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U382 ( .A(KEYINPUT21), .B(G218GAT), .Z(n329) );
  XNOR2_X1 U383 ( .A(KEYINPUT89), .B(G197GAT), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U385 ( .A(KEYINPUT90), .B(n330), .Z(n342) );
  XOR2_X1 U386 ( .A(n331), .B(n342), .Z(n469) );
  XOR2_X1 U387 ( .A(G211GAT), .B(G8GAT), .Z(n390) );
  XOR2_X1 U388 ( .A(G92GAT), .B(G64GAT), .Z(n346) );
  XOR2_X1 U389 ( .A(n390), .B(n346), .Z(n333) );
  NAND2_X1 U390 ( .A1(G226GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U392 ( .A(KEYINPUT78), .B(G36GAT), .Z(n413) );
  XOR2_X1 U393 ( .A(n334), .B(n413), .Z(n340) );
  XOR2_X1 U394 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n336) );
  XNOR2_X1 U395 ( .A(G204GAT), .B(G176GAT), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n524) );
  XOR2_X1 U400 ( .A(KEYINPUT46), .B(KEYINPUT118), .Z(n379) );
  INV_X1 U401 ( .A(KEYINPUT41), .ZN(n358) );
  XOR2_X1 U402 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n344) );
  XNOR2_X1 U403 ( .A(G78GAT), .B(KEYINPUT72), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n357) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n355) );
  XNOR2_X1 U406 ( .A(G57GAT), .B(G71GAT), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n347), .B(KEYINPUT13), .ZN(n385) );
  XOR2_X1 U408 ( .A(G85GAT), .B(G99GAT), .Z(n411) );
  NAND2_X1 U409 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n294), .B(n348), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n349), .B(KEYINPUT32), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n358), .B(n581), .ZN(n553) );
  INV_X1 U414 ( .A(n553), .ZN(n566) );
  XOR2_X1 U415 ( .A(KEYINPUT67), .B(G8GAT), .Z(n360) );
  XNOR2_X1 U416 ( .A(G1GAT), .B(G169GAT), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U418 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n362) );
  XNOR2_X1 U419 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n377) );
  XNOR2_X1 U422 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n365), .B(KEYINPUT7), .ZN(n407) );
  XOR2_X1 U424 ( .A(n407), .B(KEYINPUT68), .Z(n367) );
  NAND2_X1 U425 ( .A1(G229GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U427 ( .A(G15GAT), .B(G197GAT), .Z(n369) );
  XNOR2_X1 U428 ( .A(G141GAT), .B(G113GAT), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U431 ( .A(G43GAT), .B(G50GAT), .Z(n373) );
  XNOR2_X1 U432 ( .A(G36GAT), .B(G22GAT), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n576) );
  NAND2_X1 U436 ( .A1(n566), .A2(n576), .ZN(n378) );
  XOR2_X1 U437 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n381) );
  XNOR2_X1 U438 ( .A(KEYINPUT12), .B(KEYINPUT82), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n398) );
  XOR2_X1 U440 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n383) );
  NAND2_X1 U441 ( .A1(G231GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U443 ( .A(n384), .B(KEYINPUT80), .Z(n388) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n394) );
  XOR2_X1 U446 ( .A(n389), .B(G64GAT), .Z(n392) );
  XNOR2_X1 U447 ( .A(G183GAT), .B(n390), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U449 ( .A(n394), .B(n393), .Z(n396) );
  XNOR2_X1 U450 ( .A(G1GAT), .B(KEYINPUT14), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n558) );
  XOR2_X1 U453 ( .A(KEYINPUT117), .B(n558), .Z(n572) );
  XOR2_X1 U454 ( .A(KEYINPUT75), .B(KEYINPUT65), .Z(n400) );
  XNOR2_X1 U455 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n421) );
  XOR2_X1 U457 ( .A(KEYINPUT74), .B(G106GAT), .Z(n402) );
  XNOR2_X1 U458 ( .A(KEYINPUT77), .B(G218GAT), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U460 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n404) );
  XNOR2_X1 U461 ( .A(G92GAT), .B(KEYINPUT76), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U463 ( .A(n406), .B(n405), .Z(n419) );
  XOR2_X1 U464 ( .A(G190GAT), .B(n407), .Z(n409) );
  NAND2_X1 U465 ( .A1(G232GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n417) );
  XOR2_X1 U467 ( .A(n411), .B(n410), .Z(n415) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U472 ( .A(n421), .B(n420), .Z(n561) );
  XNOR2_X1 U473 ( .A(n424), .B(KEYINPUT47), .ZN(n430) );
  XOR2_X1 U474 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n426) );
  INV_X1 U475 ( .A(n558), .ZN(n585) );
  XNOR2_X1 U476 ( .A(n561), .B(KEYINPUT36), .ZN(n588) );
  NAND2_X1 U477 ( .A1(n585), .A2(n588), .ZN(n425) );
  XNOR2_X1 U478 ( .A(n426), .B(n425), .ZN(n427) );
  NAND2_X1 U479 ( .A1(n427), .A2(n581), .ZN(n428) );
  NOR2_X1 U480 ( .A1(n428), .A2(n576), .ZN(n429) );
  NOR2_X1 U481 ( .A1(n430), .A2(n429), .ZN(n431) );
  XNOR2_X1 U482 ( .A(KEYINPUT48), .B(n431), .ZN(n533) );
  NOR2_X1 U483 ( .A1(n524), .A2(n533), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n432), .B(KEYINPUT54), .ZN(n455) );
  XOR2_X1 U485 ( .A(G134GAT), .B(G85GAT), .Z(n434) );
  XNOR2_X1 U486 ( .A(KEYINPUT77), .B(G29GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U488 ( .A(n436), .B(n435), .Z(n438) );
  NAND2_X1 U489 ( .A1(G225GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U491 ( .A(n439), .B(KEYINPUT1), .Z(n442) );
  XNOR2_X1 U492 ( .A(n440), .B(KEYINPUT97), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U494 ( .A(G120GAT), .B(G148GAT), .Z(n444) );
  XNOR2_X1 U495 ( .A(G162GAT), .B(G155GAT), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U497 ( .A(n446), .B(n445), .Z(n454) );
  XOR2_X1 U498 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n448) );
  XNOR2_X1 U499 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U501 ( .A(KEYINPUT6), .B(G57GAT), .Z(n450) );
  XNOR2_X1 U502 ( .A(G1GAT), .B(G127GAT), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n454), .B(n453), .ZN(n522) );
  NAND2_X1 U506 ( .A1(n455), .A2(n522), .ZN(n574) );
  NOR2_X1 U507 ( .A1(n469), .A2(n574), .ZN(n456) );
  XNOR2_X1 U508 ( .A(n456), .B(KEYINPUT55), .ZN(n457) );
  AND2_X1 U509 ( .A1(n570), .A2(n561), .ZN(n461) );
  XNOR2_X1 U510 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n459) );
  INV_X1 U511 ( .A(G190GAT), .ZN(n458) );
  XNOR2_X1 U512 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n486) );
  NAND2_X1 U513 ( .A1(n576), .A2(n581), .ZN(n496) );
  XNOR2_X1 U514 ( .A(KEYINPUT27), .B(KEYINPUT100), .ZN(n462) );
  XNOR2_X1 U515 ( .A(n462), .B(n524), .ZN(n472) );
  NOR2_X1 U516 ( .A1(n522), .A2(n472), .ZN(n463) );
  XOR2_X1 U517 ( .A(KEYINPUT101), .B(n463), .Z(n532) );
  XNOR2_X1 U518 ( .A(KEYINPUT28), .B(n469), .ZN(n537) );
  XNOR2_X1 U519 ( .A(KEYINPUT87), .B(n526), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n537), .A2(n464), .ZN(n465) );
  NAND2_X1 U521 ( .A1(n532), .A2(n465), .ZN(n478) );
  NOR2_X1 U522 ( .A1(n526), .A2(n524), .ZN(n466) );
  XOR2_X1 U523 ( .A(KEYINPUT103), .B(n466), .Z(n467) );
  NOR2_X1 U524 ( .A1(n469), .A2(n467), .ZN(n468) );
  XNOR2_X1 U525 ( .A(n468), .B(KEYINPUT25), .ZN(n474) );
  AND2_X1 U526 ( .A1(n469), .A2(n526), .ZN(n471) );
  XNOR2_X1 U527 ( .A(KEYINPUT102), .B(KEYINPUT26), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n471), .B(n470), .ZN(n549) );
  INV_X1 U529 ( .A(n549), .ZN(n575) );
  OR2_X1 U530 ( .A1(n575), .A2(n472), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n522), .A2(n475), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT104), .B(n476), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n479), .B(KEYINPUT105), .ZN(n494) );
  NOR2_X1 U536 ( .A1(n561), .A2(n558), .ZN(n480) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(n480), .Z(n481) );
  NOR2_X1 U538 ( .A1(n494), .A2(n481), .ZN(n482) );
  XOR2_X1 U539 ( .A(KEYINPUT106), .B(n482), .Z(n510) );
  NOR2_X1 U540 ( .A1(n496), .A2(n510), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n483), .B(KEYINPUT107), .ZN(n491) );
  NOR2_X1 U542 ( .A1(n522), .A2(n491), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT108), .B(n484), .Z(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(G1324GAT) );
  NOR2_X1 U545 ( .A1(n524), .A2(n491), .ZN(n488) );
  XNOR2_X1 U546 ( .A(G8GAT), .B(KEYINPUT109), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(G1325GAT) );
  NOR2_X1 U548 ( .A1(n526), .A2(n491), .ZN(n490) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  INV_X1 U551 ( .A(n537), .ZN(n529) );
  NOR2_X1 U552 ( .A1(n529), .A2(n491), .ZN(n492) );
  XOR2_X1 U553 ( .A(G22GAT), .B(n492), .Z(G1327GAT) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  NAND2_X1 U555 ( .A1(n558), .A2(n588), .ZN(n493) );
  NOR2_X1 U556 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U557 ( .A(KEYINPUT37), .B(n495), .ZN(n521) );
  NOR2_X1 U558 ( .A1(n496), .A2(n521), .ZN(n497) );
  XOR2_X1 U559 ( .A(KEYINPUT38), .B(n497), .Z(n505) );
  NOR2_X1 U560 ( .A1(n522), .A2(n505), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U562 ( .A1(n505), .A2(n524), .ZN(n500) );
  XOR2_X1 U563 ( .A(KEYINPUT110), .B(n500), .Z(n501) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  XNOR2_X1 U565 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n503) );
  NOR2_X1 U566 ( .A1(n526), .A2(n505), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  NOR2_X1 U569 ( .A1(n505), .A2(n529), .ZN(n507) );
  XNOR2_X1 U570 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(n508), .ZN(G1331GAT) );
  INV_X1 U573 ( .A(n576), .ZN(n550) );
  NAND2_X1 U574 ( .A1(n550), .A2(n566), .ZN(n509) );
  XOR2_X1 U575 ( .A(KEYINPUT115), .B(n509), .Z(n520) );
  OR2_X1 U576 ( .A1(n510), .A2(n520), .ZN(n517) );
  NOR2_X1 U577 ( .A1(n517), .A2(n522), .ZN(n514) );
  XOR2_X1 U578 ( .A(KEYINPUT114), .B(KEYINPUT116), .Z(n512) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U582 ( .A1(n524), .A2(n517), .ZN(n515) );
  XOR2_X1 U583 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U584 ( .A1(n526), .A2(n517), .ZN(n516) );
  XOR2_X1 U585 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U586 ( .A1(n529), .A2(n517), .ZN(n519) );
  XNOR2_X1 U587 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U588 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  OR2_X1 U589 ( .A1(n521), .A2(n520), .ZN(n528) );
  NOR2_X1 U590 ( .A1(n522), .A2(n528), .ZN(n523) );
  XOR2_X1 U591 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U592 ( .A1(n524), .A2(n528), .ZN(n525) );
  XOR2_X1 U593 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U594 ( .A1(n526), .A2(n528), .ZN(n527) );
  XOR2_X1 U595 ( .A(G99GAT), .B(n527), .Z(G1338GAT) );
  NOR2_X1 U596 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(n530), .Z(n531) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  INV_X1 U599 ( .A(n532), .ZN(n534) );
  NOR2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n548), .A2(n535), .ZN(n536) );
  NOR2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n576), .A2(n545), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U606 ( .A1(n545), .A2(n566), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(G120GAT), .B(n541), .Z(G1341GAT) );
  INV_X1 U609 ( .A(n545), .ZN(n542) );
  NOR2_X1 U610 ( .A1(n572), .A2(n542), .ZN(n543) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(n543), .Z(n544) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U614 ( .A1(n545), .A2(n561), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n562) );
  NOR2_X1 U617 ( .A1(n550), .A2(n562), .ZN(n551) );
  XOR2_X1 U618 ( .A(G141GAT), .B(n551), .Z(n552) );
  XNOR2_X1 U619 ( .A(KEYINPUT120), .B(n552), .ZN(G1344GAT) );
  NOR2_X1 U620 ( .A1(n562), .A2(n553), .ZN(n557) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n558), .A2(n562), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT122), .B(n559), .Z(n560) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n560), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n422), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(KEYINPUT123), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n576), .A2(n570), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n568) );
  NAND2_X1 U634 ( .A1(n570), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(n569), .ZN(G1349GAT) );
  INV_X1 U637 ( .A(n570), .ZN(n571) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(G183GAT), .B(n573), .Z(G1350GAT) );
  XOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT60), .Z(n578) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n589) );
  NAND2_X1 U642 ( .A1(n589), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U647 ( .A(n581), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n589), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(KEYINPUT126), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(n587), .ZN(G1354GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n591) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

