//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942;
  NOR2_X1   g000(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G120gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n207));
  OAI21_X1  g006(.A(G120gat), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G127gat), .B(G134gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n209), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G113gat), .B2(G120gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n219));
  AND2_X1   g018(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n218), .A2(new_n219), .B1(new_n220), .B2(G190gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(KEYINPUT23), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G176gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G169gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228));
  NOR4_X1   g027(.A1(new_n221), .A2(new_n224), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230));
  AND2_X1   g029(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n226), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n230), .B1(new_n233), .B2(new_n224), .ZN(new_n234));
  OR2_X1    g033(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n235), .A2(KEYINPUT23), .A3(new_n225), .A4(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n222), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT23), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n240), .A3(KEYINPUT65), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n219), .A2(new_n218), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n220), .A2(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n234), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n229), .B1(new_n245), .B2(new_n228), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT26), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n238), .A2(new_n247), .A3(new_n223), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n222), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT68), .ZN(new_n251));
  INV_X1    g050(.A(G183gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT27), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT27), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G183gat), .ZN(new_n255));
  INV_X1    g054(.A(G190gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n248), .A2(new_n249), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n257), .A3(KEYINPUT66), .ZN(new_n264));
  AND4_X1   g063(.A1(new_n251), .A2(new_n261), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n217), .B1(new_n246), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G227gat), .A2(G233gat), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n251), .A2(new_n261), .A3(new_n263), .A4(new_n264), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n237), .A2(new_n240), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n221), .B1(new_n269), .B2(new_n230), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT25), .B1(new_n270), .B2(new_n241), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n216), .B(new_n268), .C1(new_n271), .C2(new_n229), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n266), .A2(new_n267), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT32), .ZN(new_n274));
  XNOR2_X1  g073(.A(G15gat), .B(G43gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G71gat), .B(G99gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n274), .B1(KEYINPUT33), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT33), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n273), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n278), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n285), .B1(new_n273), .B2(KEYINPUT32), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n273), .A2(new_n285), .A3(KEYINPUT32), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n281), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n277), .B1(new_n273), .B2(new_n282), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n290), .A2(new_n281), .A3(new_n288), .A4(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n280), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n267), .B1(new_n266), .B2(new_n272), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT34), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(new_n296), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n290), .A2(new_n288), .A3(new_n291), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT72), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n279), .B1(new_n302), .B2(new_n292), .ZN(new_n303));
  INV_X1    g102(.A(new_n299), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(G228gat), .A2(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G197gat), .B(G204gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT22), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n308), .A3(new_n312), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(KEYINPUT75), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n313), .A2(new_n319), .A3(new_n315), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n318), .A2(KEYINPUT76), .A3(new_n320), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(G155gat), .ZN(new_n327));
  INV_X1    g126(.A(G162gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G141gat), .B(G148gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n326), .B(new_n329), .C1(new_n330), .C2(KEYINPUT2), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332));
  INV_X1    g131(.A(G141gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G148gat), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G141gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n326), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n326), .A2(KEYINPUT2), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n331), .A2(new_n332), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n307), .B1(new_n325), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n332), .B1(new_n321), .B2(KEYINPUT29), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n331), .A2(new_n340), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n321), .A2(new_n343), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT84), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(KEYINPUT29), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n316), .A2(KEYINPUT84), .A3(new_n317), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT3), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n346), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n349), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n307), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n348), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(KEYINPUT86), .A3(G22gat), .ZN(new_n358));
  INV_X1    g157(.A(G22gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n348), .A2(new_n359), .A3(new_n356), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT85), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n344), .A2(new_n347), .B1(new_n307), .B2(new_n355), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(new_n359), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(KEYINPUT85), .A3(new_n359), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n358), .A2(new_n362), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT31), .B(G50gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n360), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n364), .A2(new_n359), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n372), .A2(new_n373), .A3(new_n370), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n300), .A2(new_n305), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT87), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n216), .A2(new_n346), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n211), .A2(new_n331), .A3(new_n215), .A4(new_n340), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n384), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n381), .A2(KEYINPUT4), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n346), .A2(KEYINPUT3), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n216), .A3(new_n341), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n386), .B1(new_n392), .B2(new_n383), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT82), .B1(new_n381), .B2(KEYINPUT4), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n381), .A2(new_n387), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n381), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n397));
  OAI211_X1 g196(.A(KEYINPUT5), .B(new_n391), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n385), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G1gat), .B(G29gat), .Z(new_n400));
  XNOR2_X1  g199(.A(G57gat), .B(G85gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  OAI21_X1  g203(.A(new_n379), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n404), .ZN(new_n406));
  AOI211_X1 g205(.A(new_n406), .B(new_n385), .C1(new_n393), .C2(new_n398), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n378), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n398), .ZN(new_n409));
  INV_X1    g208(.A(new_n385), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n406), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n399), .A2(new_n404), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n412), .A2(KEYINPUT87), .A3(new_n379), .A4(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n406), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n408), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G8gat), .B(G36gat), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT80), .ZN(new_n418));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT77), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n246), .A2(new_n265), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(KEYINPUT29), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n321), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n423), .B1(new_n246), .B2(new_n265), .ZN(new_n430));
  OAI211_X1 g229(.A(KEYINPUT79), .B(new_n424), .C1(new_n425), .C2(KEYINPUT29), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT78), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(KEYINPUT78), .B(new_n423), .C1(new_n246), .C2(new_n265), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n426), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n325), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n421), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n432), .A2(new_n421), .A3(new_n437), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n440), .B2(KEYINPUT30), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT35), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n416), .A2(new_n441), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT88), .B1(new_n377), .B2(new_n445), .ZN(new_n446));
  AND4_X1   g245(.A1(new_n442), .A2(new_n416), .A3(new_n444), .A4(new_n441), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n302), .A2(new_n292), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n304), .B1(new_n448), .B2(new_n280), .ZN(new_n449));
  AOI211_X1 g248(.A(new_n279), .B(new_n299), .C1(new_n302), .C2(new_n292), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n447), .A2(new_n451), .A3(new_n452), .A4(new_n376), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n446), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT73), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n294), .A2(new_n455), .A3(new_n299), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT73), .B1(new_n303), .B2(new_n304), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n305), .A4(new_n376), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT89), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n450), .B1(new_n449), .B2(new_n455), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n461), .A2(KEYINPUT89), .A3(new_n457), .A4(new_n376), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n441), .A2(new_n444), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n412), .A2(new_n379), .A3(new_n413), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n464), .A2(new_n415), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n460), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n454), .B1(new_n467), .B2(KEYINPUT35), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT74), .B1(new_n451), .B2(KEYINPUT36), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT36), .A4(new_n305), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT74), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT36), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n471), .B(new_n472), .C1(new_n449), .C2(new_n450), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n466), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n374), .B1(new_n367), .B2(new_n370), .ZN(new_n476));
  INV_X1    g275(.A(new_n416), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n478), .A2(new_n321), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n436), .A2(new_n325), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT37), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT38), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT37), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n432), .A2(new_n483), .A3(new_n437), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n481), .A2(new_n482), .A3(new_n420), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n420), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n483), .B1(new_n432), .B2(new_n437), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT38), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n477), .A2(new_n485), .A3(new_n488), .A4(new_n439), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n392), .A2(new_n386), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(KEYINPUT39), .C1(new_n386), .C2(new_n382), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n491), .B(new_n404), .C1(KEYINPUT39), .C2(new_n490), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT40), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n412), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n493), .B2(new_n492), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n476), .B1(new_n463), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n475), .A2(new_n476), .B1(new_n489), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n474), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n468), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT95), .ZN(new_n500));
  INV_X1    g299(.A(G29gat), .ZN(new_n501));
  INV_X1    g300(.A(G36gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT14), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(G29gat), .B2(G36gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n506), .B(KEYINPUT91), .Z(new_n507));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n510));
  NAND2_X1  g309(.A1(G29gat), .A2(G36gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT92), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n511), .ZN(new_n515));
  OAI211_X1 g314(.A(KEYINPUT15), .B(new_n508), .C1(new_n506), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT16), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(G1gat), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(G1gat), .B2(new_n518), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G8gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT93), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n517), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n517), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n522), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n514), .A2(KEYINPUT17), .A3(new_n516), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n527), .A2(KEYINPUT18), .A3(new_n528), .A4(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n517), .A2(new_n525), .A3(new_n522), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n525), .B1(new_n517), .B2(new_n522), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n533), .B(new_n528), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n517), .A2(new_n522), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n535), .B2(new_n536), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n524), .A2(KEYINPUT94), .A3(new_n526), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n528), .B(KEYINPUT13), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n534), .B(new_n539), .C1(new_n544), .C2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G197gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT11), .B(G169gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n551), .B(KEYINPUT12), .Z(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT90), .Z(new_n553));
  AOI21_X1  g352(.A(new_n500), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n542), .A2(new_n543), .ZN(new_n555));
  INV_X1    g354(.A(new_n540), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n545), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n558), .A2(new_n534), .A3(new_n539), .A4(new_n552), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n547), .A2(new_n500), .A3(new_n553), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n499), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n564), .B(new_n565), .Z(new_n566));
  XOR2_X1   g365(.A(G99gat), .B(G106gat), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT99), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(G85gat), .ZN(new_n570));
  INV_X1    g369(.A(G92gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(KEYINPUT8), .A2(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n566), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n567), .A2(KEYINPUT99), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n530), .A2(new_n532), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G190gat), .B(G218gat), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  AND3_X1   g378(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n576), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(new_n517), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n577), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n579), .B1(new_n577), .B2(new_n582), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n589), .A2(KEYINPUT100), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(KEYINPUT100), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n585), .A2(new_n591), .ZN(new_n593));
  AND2_X1   g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  XOR2_X1   g394(.A(G57gat), .B(G64gat), .Z(new_n596));
  AOI211_X1 g395(.A(new_n594), .B(new_n595), .C1(new_n596), .C2(KEYINPUT9), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n594), .B1(KEYINPUT9), .B2(new_n595), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT96), .B(G57gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G64gat), .ZN(new_n600));
  INV_X1    g399(.A(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G57gat), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n598), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n604), .A2(new_n607), .A3(new_n605), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(G127gat), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n603), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n522), .B1(KEYINPUT21), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n609), .A2(new_n612), .A3(new_n610), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n611), .A2(new_n612), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n615), .B1(new_n620), .B2(new_n617), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n327), .ZN(new_n623));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  NAND3_X1  g424(.A1(new_n619), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n619), .B2(new_n621), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n592), .B(new_n593), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n576), .A2(new_n604), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n573), .A2(new_n574), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n573), .A2(new_n574), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n614), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n630), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n581), .A2(KEYINPUT10), .A3(new_n614), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n581), .A2(KEYINPUT101), .A3(KEYINPUT10), .A4(new_n614), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT102), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n638), .A2(new_n643), .A3(new_n639), .A4(new_n640), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n639), .B1(new_n630), .B2(new_n634), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n644), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n641), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n649), .B1(new_n652), .B2(new_n645), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n629), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n563), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n465), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(G1gat), .Z(G1324gat));
  NAND3_X1  g458(.A1(new_n563), .A2(new_n463), .A3(new_n655), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR4_X1   g462(.A1(new_n660), .A2(KEYINPUT103), .A3(new_n661), .A4(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n661), .B1(new_n660), .B2(G8gat), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n660), .A2(new_n663), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n666), .B2(KEYINPUT42), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n664), .B1(new_n667), .B2(new_n669), .ZN(G1325gat));
  INV_X1    g469(.A(G15gat), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n656), .A2(new_n671), .A3(new_n474), .ZN(new_n672));
  INV_X1    g471(.A(new_n451), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n656), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(KEYINPUT104), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(KEYINPUT104), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n672), .B1(new_n675), .B2(new_n676), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n656), .A2(new_n376), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  AND3_X1   g479(.A1(new_n547), .A2(new_n500), .A3(new_n553), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n559), .B2(new_n554), .ZN(new_n682));
  INV_X1    g481(.A(new_n628), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n626), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n654), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n593), .A2(new_n592), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT105), .Z(new_n688));
  OAI211_X1 g487(.A(new_n682), .B(new_n688), .C1(new_n468), .C2(new_n498), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(G29gat), .A3(new_n657), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT45), .Z(new_n691));
  OAI21_X1  g490(.A(new_n686), .B1(new_n468), .B2(new_n498), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g493(.A(KEYINPUT44), .B(new_n686), .C1(new_n468), .C2(new_n498), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n682), .A2(new_n685), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n696), .A2(new_n465), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n691), .B1(new_n501), .B2(new_n698), .ZN(G1328gat));
  INV_X1    g498(.A(new_n463), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n689), .A2(G36gat), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT46), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n696), .A2(new_n463), .A3(new_n697), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n703), .B2(new_n502), .ZN(G1329gat));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT106), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n673), .A2(G43gat), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n689), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n474), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n694), .A2(new_n710), .A3(new_n695), .A4(new_n697), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(G43gat), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n705), .A2(KEYINPUT106), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1330gat));
  OR3_X1    g513(.A1(new_n689), .A2(G50gat), .A3(new_n376), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(KEYINPUT48), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n694), .A2(new_n476), .A3(new_n695), .A4(new_n697), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT107), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G50gat), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n717), .A2(KEYINPUT107), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(G50gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n715), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n721), .A2(new_n725), .ZN(G1331gat));
  INV_X1    g525(.A(new_n686), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n562), .A2(new_n684), .A3(new_n727), .A4(new_n654), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n499), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n465), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(new_n599), .Z(G1332gat));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n463), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT49), .B(G64gat), .Z(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(G1333gat));
  NAND2_X1  g534(.A1(new_n729), .A2(new_n451), .ZN(new_n736));
  INV_X1    g535(.A(G71gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n474), .A2(new_n737), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n729), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n739), .B1(new_n729), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n738), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n476), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n682), .A2(new_n684), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n654), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT109), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n694), .A2(new_n465), .A3(new_n695), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT110), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G85gat), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n750), .A2(KEYINPUT110), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n474), .A2(new_n497), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n467), .A2(KEYINPUT35), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(new_n454), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n756), .A2(KEYINPUT51), .A3(new_n686), .A4(new_n747), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n686), .B(new_n747), .C1(new_n468), .C2(new_n498), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n465), .A2(new_n570), .A3(new_n654), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT111), .Z(new_n764));
  OAI22_X1  g563(.A1(new_n752), .A2(new_n753), .B1(new_n762), .B2(new_n764), .ZN(G1336gat));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT112), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n694), .A2(new_n463), .A3(new_n695), .A4(new_n749), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n766), .A2(KEYINPUT112), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n654), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n700), .A2(G92gat), .A3(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n758), .A2(new_n759), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND4_X1   g575(.A1(new_n767), .A2(new_n769), .A3(new_n771), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n770), .B1(new_n761), .B2(new_n773), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n767), .B1(new_n778), .B2(new_n769), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n777), .A2(new_n779), .ZN(G1337gat));
  NAND3_X1  g579(.A1(new_n696), .A2(new_n710), .A3(new_n749), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G99gat), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n772), .A2(G99gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n761), .A2(new_n451), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1338gat));
  NAND4_X1  g584(.A1(new_n694), .A2(new_n476), .A3(new_n695), .A4(new_n749), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n376), .A2(new_n772), .A3(G106gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n762), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT53), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n787), .B(new_n791), .C1(new_n762), .C2(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1339gat));
  NAND2_X1  g592(.A1(new_n638), .A2(new_n640), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(G230gat), .A3(G233gat), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n642), .A2(new_n795), .A3(KEYINPUT54), .A4(new_n644), .ZN(new_n796));
  XNOR2_X1  g595(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n648), .B1(new_n652), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n555), .A2(new_n556), .A3(new_n546), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n527), .A2(new_n533), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(G229gat), .A3(G233gat), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n551), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n547), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n552), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n796), .A2(KEYINPUT55), .A3(new_n798), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n801), .A2(new_n807), .A3(new_n808), .A4(new_n651), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n684), .B1(new_n809), .B2(new_n686), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n686), .B1(new_n807), .B2(new_n654), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n801), .A2(new_n651), .A3(new_n808), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n562), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n727), .A2(new_n772), .A3(new_n684), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n682), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n655), .A2(new_n562), .A3(KEYINPUT113), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n810), .A2(new_n813), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n818), .A2(new_n657), .A3(new_n463), .ZN(new_n819));
  INV_X1    g618(.A(new_n377), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n562), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n460), .A2(new_n462), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n562), .A2(new_n207), .A3(new_n206), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT115), .Z(new_n827));
  OAI21_X1  g626(.A(new_n823), .B1(new_n825), .B2(new_n827), .ZN(G1340gat));
  INV_X1    g627(.A(new_n825), .ZN(new_n829));
  AOI21_X1  g628(.A(G120gat), .B1(new_n829), .B2(new_n654), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n772), .A2(new_n204), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n821), .B2(new_n831), .ZN(G1341gat));
  INV_X1    g631(.A(new_n684), .ZN(new_n833));
  OAI21_X1  g632(.A(G127gat), .B1(new_n822), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n829), .A2(new_n612), .A3(new_n684), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1342gat));
  OR3_X1    g635(.A1(new_n825), .A2(G134gat), .A3(new_n727), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n686), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n837), .A2(KEYINPUT56), .B1(new_n838), .B2(G134gat), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n837), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G1343gat));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n818), .B2(new_n376), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n810), .A2(new_n813), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n816), .A2(new_n817), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(KEYINPUT57), .A3(new_n476), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n463), .A2(new_n657), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n474), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT117), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n855), .A3(new_n682), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n856), .A2(G141gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n818), .A2(new_n376), .ZN(new_n858));
  INV_X1    g657(.A(new_n854), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(G141gat), .A3(new_n562), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n845), .B(KEYINPUT58), .C1(new_n857), .C2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n856), .B2(G141gat), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT118), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT58), .B1(new_n861), .B2(KEYINPUT119), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(KEYINPUT119), .B2(new_n861), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n862), .B(new_n865), .C1(new_n857), .C2(new_n867), .ZN(G1344gat));
  NAND4_X1  g667(.A1(new_n858), .A2(new_n335), .A3(new_n654), .A4(new_n859), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G148gat), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n852), .A2(new_n855), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n654), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n655), .A2(new_n562), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n376), .B1(new_n848), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n851), .B1(KEYINPUT57), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n654), .A3(new_n855), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n870), .B1(new_n877), .B2(G148gat), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n869), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(KEYINPUT120), .B(new_n869), .C1(new_n873), .C2(new_n878), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1345gat));
  AOI21_X1  g682(.A(new_n327), .B1(new_n872), .B2(new_n684), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n860), .A2(G155gat), .A3(new_n833), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n884), .A2(new_n885), .ZN(G1346gat));
  NAND2_X1  g685(.A1(new_n872), .A2(new_n686), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n328), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n888), .B2(new_n887), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n376), .A2(new_n727), .A3(G162gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n819), .A2(new_n474), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1347gat));
  NOR3_X1   g692(.A1(new_n818), .A2(new_n465), .A3(new_n700), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n820), .ZN(new_n895));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895), .B2(new_n562), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n824), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n682), .A2(new_n235), .A3(new_n236), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(G1348gat));
  NAND4_X1  g698(.A1(new_n894), .A2(G176gat), .A3(new_n820), .A4(new_n654), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n894), .A2(new_n824), .A3(new_n654), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n901), .A2(KEYINPUT122), .A3(new_n225), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT122), .B1(new_n901), .B2(new_n225), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n904), .B(KEYINPUT123), .Z(G1349gat));
  NOR2_X1   g704(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n906));
  INV_X1    g705(.A(new_n897), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n907), .A2(new_n253), .A3(new_n255), .A4(new_n684), .ZN(new_n908));
  OAI21_X1  g707(.A(G183gat), .B1(new_n895), .B2(new_n833), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT125), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n910), .B(new_n912), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n895), .B2(new_n727), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT61), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n907), .A2(new_n256), .A3(new_n686), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1351gat));
  NOR3_X1   g716(.A1(new_n710), .A2(new_n465), .A3(new_n700), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n858), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(G197gat), .B1(new_n920), .B2(new_n682), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n876), .A2(new_n918), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n682), .A2(G197gat), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(G1352gat));
  NOR3_X1   g723(.A1(new_n919), .A2(G204gat), .A3(new_n772), .ZN(new_n925));
  XNOR2_X1  g724(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n876), .A2(new_n654), .A3(new_n918), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G204gat), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1353gat));
  NAND3_X1  g729(.A1(new_n876), .A2(new_n684), .A3(new_n918), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G211gat), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n934), .A2(KEYINPUT127), .A3(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n932), .A2(new_n937), .A3(new_n933), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n920), .A2(new_n310), .A3(new_n684), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(G1354gat));
  NAND3_X1  g739(.A1(new_n920), .A2(new_n311), .A3(new_n686), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n922), .A2(new_n686), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n311), .ZN(G1355gat));
endmodule


