//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n441, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n565, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G108), .ZN(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n441), .A2(G57), .A3(G69), .A4(G120), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT67), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n454));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G2106), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n453), .A2(G567), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n467), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n471), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT69), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n464), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n477), .A2(new_n479), .A3(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT70), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n477), .A2(new_n479), .A3(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n468), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n484), .A2(G136), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND3_X1  g065(.A1(new_n463), .A2(G102), .A3(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n464), .B2(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n491), .B1(new_n494), .B2(new_n463), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(new_n464), .B2(new_n499), .ZN(new_n500));
  AND4_X1   g075(.A1(new_n469), .A2(new_n499), .A3(new_n471), .A4(new_n497), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n495), .A2(new_n502), .ZN(G164));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT72), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n504), .A2(KEYINPUT72), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n505), .B(new_n506), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT73), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n508), .B(new_n510), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(G543), .B1(new_n516), .B2(new_n517), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n513), .A2(new_n524), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n515), .A2(new_n523), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  INV_X1    g102(.A(new_n518), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT76), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n532), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n508), .A2(new_n510), .A3(G63), .A4(G651), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n537));
  OR2_X1    g112(.A1(KEYINPUT74), .A2(G51), .ZN(new_n538));
  NAND2_X1  g113(.A1(KEYINPUT74), .A2(G51), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n536), .B(new_n537), .C1(new_n520), .C2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT6), .B(G651), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n543), .A2(G543), .A3(new_n538), .A4(new_n539), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n537), .B1(new_n544), .B2(new_n536), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n529), .B(new_n535), .C1(new_n542), .C2(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  XNOR2_X1  g122(.A(KEYINPUT5), .B(G543), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n543), .A2(new_n548), .A3(G90), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT77), .B(G52), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n548), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G651), .ZN(new_n552));
  OAI221_X1 g127(.A(new_n549), .B1(new_n520), .B2(new_n550), .C1(new_n551), .C2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND3_X1  g129(.A1(new_n508), .A2(new_n510), .A3(G56), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n555), .A2(KEYINPUT78), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT78), .B1(new_n555), .B2(new_n556), .ZN(new_n558));
  NOR3_X1   g133(.A1(new_n557), .A2(new_n558), .A3(new_n552), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  INV_X1    g135(.A(G43), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n518), .A2(new_n560), .B1(new_n520), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(G188));
  INV_X1    g144(.A(G78), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT79), .B1(new_n570), .B2(new_n507), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n572), .A2(G78), .A3(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n571), .B(new_n573), .C1(new_n511), .C2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(G651), .B1(new_n528), .B2(G91), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n543), .A2(G53), .A3(G543), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n520), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n580), .A2(KEYINPUT9), .A3(G53), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n576), .A2(new_n579), .A3(new_n581), .ZN(G299));
  OAI21_X1  g157(.A(G651), .B1(new_n548), .B2(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n543), .A2(new_n548), .A3(G87), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n543), .A2(G49), .A3(G543), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(KEYINPUT80), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G288));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n548), .B2(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n591), .B1(new_n594), .B2(new_n552), .ZN(new_n595));
  OAI211_X1 g170(.A(G48), .B(G543), .C1(new_n516), .C2(new_n517), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n518), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n508), .A2(new_n510), .A3(G61), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(new_n592), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n601), .A2(KEYINPUT81), .A3(G651), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n595), .A2(new_n599), .A3(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n548), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(new_n552), .ZN(new_n605));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  INV_X1    g181(.A(G47), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n518), .A2(new_n606), .B1(new_n520), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n511), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(new_n580), .B2(G54), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT10), .B1(new_n518), .B2(new_n616), .ZN(new_n617));
  OR3_X1    g192(.A1(new_n518), .A2(KEYINPUT10), .A3(new_n616), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n611), .B1(new_n620), .B2(G868), .ZN(G284));
  OAI21_X1  g196(.A(new_n611), .B1(new_n620), .B2(G868), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  XNOR2_X1  g198(.A(G299), .B(KEYINPUT82), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G297));
  OAI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n620), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n484), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n480), .A2(G123), .ZN(new_n634));
  OR2_X1    g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n635), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND3_X1  g213(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  OR2_X1    g220(.A1(G2451), .A2(G2454), .ZN(new_n646));
  NAND2_X1  g221(.A1(G2451), .A2(G2454), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT16), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT16), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n646), .A2(new_n650), .A3(new_n647), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n649), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n653), .B1(new_n649), .B2(new_n651), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n645), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n649), .A2(new_n651), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(new_n652), .ZN(new_n658));
  INV_X1    g233(.A(new_n645), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n649), .A2(new_n651), .A3(new_n653), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2427), .B(G2430), .ZN(new_n663));
  OR2_X1    g238(.A1(KEYINPUT15), .A2(G2435), .ZN(new_n664));
  NAND2_X1  g239(.A1(KEYINPUT15), .A2(G2435), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT83), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n664), .A2(new_n668), .A3(new_n665), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n667), .A2(G2438), .A3(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(G2438), .B1(new_n667), .B2(new_n669), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n663), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(new_n669), .ZN(new_n674));
  INV_X1    g249(.A(G2438), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n663), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(new_n677), .A3(new_n670), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n673), .A2(new_n678), .A3(KEYINPUT14), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n662), .B(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(KEYINPUT84), .B1(new_n680), .B2(G14), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n656), .A2(new_n661), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n682), .ZN(new_n684));
  AND4_X1   g259(.A1(KEYINPUT84), .A2(new_n683), .A3(G14), .A4(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n685), .ZN(G401));
  XOR2_X1   g261(.A(G2072), .B(G2078), .Z(new_n687));
  XOR2_X1   g262(.A(G2084), .B(G2090), .Z(new_n688));
  XNOR2_X1  g263(.A(G2067), .B(G2678), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n687), .B1(new_n690), .B2(KEYINPUT18), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G2096), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G2100), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT18), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n688), .A2(new_n689), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n695), .A2(new_n690), .A3(KEYINPUT17), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n692), .B(new_n642), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n694), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G227));
  XNOR2_X1  g277(.A(KEYINPUT22), .B(G1981), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(G1986), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1971), .B(G1976), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT19), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1956), .B(G2474), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1961), .B(G1966), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n711), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  NOR3_X1   g292(.A1(new_n711), .A2(KEYINPUT20), .A3(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT20), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n707), .B(new_n708), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n715), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n717), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n714), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n723), .B(new_n724), .C1(new_n709), .C2(new_n710), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n724), .B1(new_n720), .B2(new_n723), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n706), .B1(new_n722), .B2(new_n728), .ZN(new_n729));
  NOR3_X1   g304(.A1(new_n720), .A2(new_n723), .A3(new_n715), .ZN(new_n730));
  OAI21_X1  g305(.A(KEYINPUT20), .B1(new_n711), .B2(new_n716), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n720), .A2(new_n719), .A3(new_n715), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n727), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(new_n725), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n733), .A2(new_n735), .A3(new_n705), .ZN(new_n736));
  XNOR2_X1  g311(.A(G1991), .B(G1996), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n729), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n729), .B2(new_n736), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n704), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n722), .A2(new_n728), .A3(new_n706), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n705), .B1(new_n733), .B2(new_n735), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n737), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n729), .A2(new_n736), .A3(new_n738), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n744), .A2(new_n703), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n741), .A2(new_n746), .ZN(G229));
  XOR2_X1   g322(.A(KEYINPUT31), .B(G11), .Z(new_n748));
  NOR2_X1   g323(.A1(G5), .A2(G16), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G171), .B2(G16), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G1961), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G28), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT96), .ZN(new_n756));
  INV_X1    g331(.A(G29), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n756), .B(new_n757), .C1(new_n754), .C2(G28), .ZN(new_n758));
  OR2_X1    g333(.A1(KEYINPUT24), .A2(G34), .ZN(new_n759));
  NAND2_X1  g334(.A1(KEYINPUT24), .A2(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G160), .B2(G29), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n753), .B(new_n758), .C1(G2084), .C2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G1961), .B2(new_n750), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G16), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n766), .A2(KEYINPUT23), .A3(G20), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT23), .ZN(new_n768));
  INV_X1    g343(.A(G20), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(G16), .ZN(new_n770));
  INV_X1    g345(.A(G299), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n767), .B(new_n770), .C1(new_n771), .C2(new_n766), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT27), .B(G1996), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT93), .ZN(new_n775));
  NOR2_X1   g350(.A1(G29), .A2(G32), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n477), .A2(new_n479), .A3(G141), .A4(new_n463), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n477), .A2(new_n479), .A3(G129), .A4(G2105), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT26), .Z(new_n781));
  AND4_X1   g356(.A1(new_n777), .A2(new_n778), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n776), .B1(new_n782), .B2(G29), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n773), .B1(new_n775), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G4), .A2(G16), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n620), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT87), .B(G1348), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n766), .A2(G21), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G168), .B2(new_n766), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1966), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n757), .A2(G27), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G164), .B2(new_n757), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2078), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n757), .A2(G26), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n477), .A2(new_n479), .A3(G128), .A4(G2105), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n477), .A2(new_n479), .A3(G140), .A4(new_n463), .ZN(new_n800));
  OR2_X1    g375(.A1(G104), .A2(G2105), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n801), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n798), .B1(new_n803), .B2(new_n757), .ZN(new_n804));
  INV_X1    g379(.A(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n784), .A2(new_n788), .A3(new_n795), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n762), .A2(G2084), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT25), .Z(new_n810));
  INV_X1    g385(.A(G139), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n483), .B2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT90), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g389(.A(KEYINPUT90), .B(new_n810), .C1(new_n483), .C2(new_n811), .ZN(new_n815));
  NAND2_X1  g390(.A1(G115), .A2(G2104), .ZN(new_n816));
  INV_X1    g391(.A(G127), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n476), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G2105), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT91), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(KEYINPUT91), .A3(G2105), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n814), .A2(new_n815), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT92), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT92), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n814), .A2(new_n823), .A3(new_n826), .A4(new_n815), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n757), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(G29), .A2(G33), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT89), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(G2072), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(KEYINPUT89), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n831), .B1(new_n830), .B2(new_n833), .ZN(new_n835));
  OAI221_X1 g410(.A(new_n808), .B1(new_n775), .B2(new_n783), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT94), .ZN(new_n837));
  AOI211_X1 g412(.A(new_n765), .B(new_n807), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n757), .A2(G25), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n484), .A2(G131), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n480), .A2(G119), .ZN(new_n841));
  OR2_X1    g416(.A1(G95), .A2(G2105), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n842), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n839), .B1(new_n845), .B2(new_n757), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT35), .B(G1991), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n766), .A2(G24), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n609), .B2(new_n766), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G1986), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n848), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT86), .ZN(new_n854));
  INV_X1    g429(.A(G22), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(G16), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(G16), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(G303), .B2(G16), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n858), .B2(new_n854), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n859), .A2(G1971), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n766), .A2(G6), .ZN(new_n861));
  INV_X1    g436(.A(G305), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(new_n766), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT32), .B(G1981), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(G1971), .ZN(new_n866));
  NOR2_X1   g441(.A1(G16), .A2(G23), .ZN(new_n867));
  INV_X1    g442(.A(new_n586), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(G16), .ZN(new_n869));
  XNOR2_X1  g444(.A(KEYINPUT33), .B(G1976), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n860), .A2(new_n865), .A3(new_n866), .A4(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT34), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n853), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT36), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT36), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n878), .B(new_n853), .C1(new_n874), .C2(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n836), .A2(new_n837), .ZN(new_n881));
  INV_X1    g456(.A(G35), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT97), .B1(new_n882), .B2(G29), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n882), .A2(KEYINPUT97), .A3(G29), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n883), .B(new_n884), .C1(G162), .C2(new_n757), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT29), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(G2090), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n838), .A2(new_n880), .A3(new_n881), .A4(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n886), .A2(G2090), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(KEYINPUT98), .Z(new_n890));
  OR2_X1    g465(.A1(new_n637), .A2(new_n757), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT95), .Z(new_n892));
  NAND2_X1  g467(.A1(new_n766), .A2(G19), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n563), .B2(new_n766), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(G1341), .Z(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR4_X1   g471(.A1(new_n888), .A2(new_n890), .A3(new_n892), .A4(new_n896), .ZN(G311));
  INV_X1    g472(.A(new_n888), .ZN(new_n898));
  INV_X1    g473(.A(new_n892), .ZN(new_n899));
  INV_X1    g474(.A(new_n890), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .A4(new_n895), .ZN(G150));
  NAND3_X1  g476(.A1(new_n543), .A2(G55), .A3(G543), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n543), .A2(new_n548), .A3(G93), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n548), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n902), .B(new_n903), .C1(new_n904), .C2(new_n552), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n559), .B2(new_n562), .ZN(new_n907));
  INV_X1    g482(.A(new_n558), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n555), .A2(KEYINPUT78), .A3(new_n556), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(G651), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n562), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n905), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n619), .A2(new_n627), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(KEYINPUT39), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT100), .ZN(new_n919));
  AOI21_X1  g494(.A(G860), .B1(new_n917), .B2(KEYINPUT39), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n905), .A2(G860), .ZN(new_n922));
  XNOR2_X1  g497(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT102), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n922), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n921), .A2(new_n925), .ZN(G145));
  XOR2_X1   g501(.A(KEYINPUT106), .B(G37), .Z(new_n927));
  NAND2_X1  g502(.A1(new_n825), .A2(new_n827), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n782), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n778), .A2(new_n779), .A3(new_n777), .A4(new_n781), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n803), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n469), .A2(new_n471), .A3(G126), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n463), .B1(new_n933), .B2(new_n492), .ZN(new_n934));
  INV_X1    g509(.A(new_n491), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT104), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n937), .B(new_n491), .C1(new_n494), .C2(new_n463), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT103), .B1(new_n500), .B2(new_n501), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n499), .A2(new_n469), .A3(new_n471), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n496), .A3(KEYINPUT4), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n464), .A2(new_n497), .A3(new_n499), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n936), .A2(new_n938), .A3(new_n939), .A4(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n930), .A2(new_n932), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n945), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n782), .A2(new_n929), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n803), .A2(new_n931), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n928), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n477), .A2(new_n479), .A3(G130), .A4(G2105), .ZN(new_n953));
  OR2_X1    g528(.A1(G106), .A2(G2105), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n954), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n955));
  INV_X1    g530(.A(G142), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n953), .B(new_n955), .C1(new_n483), .C2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(new_n640), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n844), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n957), .A2(new_n640), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n640), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n845), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n945), .B1(new_n930), .B2(new_n932), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n948), .A2(new_n947), .A3(new_n949), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n824), .A3(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n951), .A2(new_n952), .A3(new_n963), .A4(new_n966), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n637), .A2(G160), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n637), .A2(G160), .ZN(new_n969));
  AND4_X1   g544(.A1(new_n488), .A2(new_n968), .A3(new_n482), .A4(new_n969), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n968), .A2(new_n969), .B1(new_n482), .B2(new_n488), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n963), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n964), .A2(new_n824), .A3(new_n965), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n964), .A2(new_n965), .B1(new_n825), .B2(new_n827), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n951), .A2(new_n963), .A3(new_n966), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(KEYINPUT105), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n927), .B1(new_n973), .B2(new_n979), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n977), .B(new_n978), .C1(new_n970), .C2(new_n971), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g558(.A(KEYINPUT108), .B1(new_n906), .B2(G868), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n609), .B(KEYINPUT107), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(G303), .A2(new_n868), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n515), .A2(new_n523), .A3(new_n525), .A4(new_n586), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(G305), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(G305), .B1(new_n987), .B2(new_n988), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n986), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n991), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(new_n985), .A3(new_n989), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT42), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n618), .A2(new_n617), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n581), .A2(new_n579), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n997), .A2(new_n576), .A3(new_n998), .A4(new_n615), .ZN(new_n999));
  NAND2_X1  g574(.A1(G299), .A2(new_n619), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n999), .A2(new_n1000), .A3(KEYINPUT41), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT41), .B1(new_n999), .B2(new_n1000), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n913), .B(new_n629), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n999), .A2(new_n1000), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1006), .B1(new_n1008), .B2(new_n1005), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n996), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G868), .ZN(new_n1011));
  MUX2_X1   g586(.A(KEYINPUT108), .B(new_n984), .S(new_n1011), .Z(G295));
  MUX2_X1   g587(.A(KEYINPUT108), .B(new_n984), .S(new_n1011), .Z(G331));
  OAI21_X1  g588(.A(new_n536), .B1(new_n520), .B2(new_n540), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT75), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n541), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1016), .A2(G301), .A3(new_n529), .A4(new_n535), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1015), .A2(new_n541), .B1(G89), .B2(new_n528), .ZN(new_n1019));
  AOI21_X1  g594(.A(G301), .B1(new_n1019), .B2(new_n535), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n913), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G286), .A2(G171), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1022), .A2(new_n912), .A3(new_n907), .A4(new_n1017), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(KEYINPUT109), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n913), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT109), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n1017), .A4(new_n1022), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1003), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1021), .A2(new_n1008), .A3(new_n1023), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n992), .A2(new_n994), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G37), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n995), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT43), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1004), .B1(new_n1023), .B2(new_n1021), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1007), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1031), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT43), .ZN(new_n1040));
  INV_X1    g615(.A(new_n927), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1034), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT44), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1035), .A2(KEYINPUT43), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT110), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1039), .A2(new_n1041), .A3(new_n1034), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT43), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT44), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1045), .B1(new_n1047), .B2(new_n1050), .ZN(G397));
  INV_X1    g626(.A(G1384), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n945), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n465), .A2(new_n466), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G2105), .ZN(new_n1057));
  INV_X1    g632(.A(new_n474), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(G40), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1996), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n931), .B(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n929), .B(new_n805), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n847), .B2(new_n844), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n847), .B2(new_n844), .ZN(new_n1066));
  AND2_X1   g641(.A1(G290), .A2(G1986), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G290), .A2(G1986), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1060), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G286), .A2(G8), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT117), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1966), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT45), .B1(new_n945), .B2(new_n1052), .ZN(new_n1075));
  INV_X1    g650(.A(G40), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n467), .A2(new_n1076), .A3(new_n474), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1052), .B1(new_n495), .B2(new_n502), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1077), .B1(new_n1078), .B2(new_n1054), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1074), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT114), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(new_n1074), .C1(new_n1075), .C2(new_n1079), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n945), .A2(new_n1084), .A3(new_n1052), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1059), .B1(new_n1078), .B2(KEYINPUT50), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1081), .B(new_n1083), .C1(G2084), .C2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1073), .B1(new_n1088), .B2(G8), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1088), .B2(new_n1073), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1090), .B(new_n1073), .C1(new_n1088), .C2(G8), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT62), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n945), .A2(new_n1052), .A3(new_n1077), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n868), .A2(G1976), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(G8), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n1098));
  INV_X1    g673(.A(G288), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(G1976), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1981), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n595), .A2(new_n599), .A3(new_n1102), .A4(new_n602), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n552), .B1(new_n600), .B2(new_n592), .ZN(new_n1104));
  OAI21_X1  g679(.A(G1981), .B1(new_n598), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT49), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1103), .A2(KEYINPUT49), .A3(new_n1105), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1108), .A2(G8), .A3(new_n1095), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1095), .A2(G8), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1103), .A2(KEYINPUT49), .A3(new_n1105), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT49), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1116), .A3(KEYINPUT113), .ZN(new_n1117));
  AOI221_X4 g692(.A(new_n1101), .B1(KEYINPUT52), .B2(new_n1097), .C1(new_n1112), .C2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n945), .A2(KEYINPUT45), .A3(new_n1052), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1059), .B1(new_n1078), .B2(new_n1054), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1971), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT111), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT112), .B(G2090), .Z(new_n1126));
  OR2_X1    g701(.A1(new_n1087), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(G1971), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT111), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(G303), .A2(G8), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT55), .Z(new_n1132));
  NAND3_X1  g707(.A1(new_n1130), .A2(G8), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1132), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1084), .B1(new_n945), .B2(new_n1052), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1077), .B1(new_n1078), .B2(KEYINPUT50), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1135), .A2(new_n1136), .A3(new_n1126), .ZN(new_n1137));
  OAI21_X1  g712(.A(G8), .B1(new_n1137), .B2(new_n1128), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1118), .A2(new_n1133), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1143), .A2(G2078), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1075), .A2(new_n1079), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(G1961), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1142), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1079), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1055), .A2(new_n1149), .A3(new_n1144), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1087), .A2(new_n752), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(KEYINPUT119), .ZN(new_n1152));
  INV_X1    g727(.A(G2078), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1119), .A2(new_n1120), .A3(new_n1153), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1148), .A2(new_n1152), .B1(new_n1143), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(G301), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1088), .A2(G8), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(KEYINPUT51), .A3(new_n1072), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1158), .B(new_n1159), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1094), .A2(new_n1141), .A3(new_n1156), .A4(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(G1348), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1095), .A2(G2067), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n619), .B1(new_n1164), .B2(KEYINPUT60), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n1166));
  NOR4_X1   g741(.A1(new_n1162), .A2(new_n1163), .A3(new_n1166), .A4(new_n620), .ZN(new_n1167));
  OAI22_X1  g742(.A1(new_n1165), .A2(new_n1167), .B1(KEYINPUT60), .B2(new_n1164), .ZN(new_n1168));
  OR3_X1    g743(.A1(new_n559), .A2(KEYINPUT116), .A3(new_n562), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1119), .A2(new_n1120), .A3(new_n1061), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT58), .B(G1341), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n1095), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1169), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT59), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(G1956), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1177));
  XNOR2_X1  g752(.A(KEYINPUT56), .B(G2072), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1119), .A2(new_n1120), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT57), .ZN(new_n1180));
  XNOR2_X1  g755(.A(G299), .B(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1177), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1168), .A2(new_n1175), .A3(new_n1184), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1186));
  AOI211_X1 g761(.A(new_n619), .B(new_n1164), .C1(new_n1186), .C2(new_n1181), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1186), .A2(new_n1181), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1140), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1158), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1154), .A2(new_n1143), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT120), .ZN(new_n1193));
  OAI21_X1  g768(.A(G40), .B1(new_n474), .B2(new_n1193), .ZN(new_n1194));
  AOI211_X1 g769(.A(new_n467), .B(new_n1194), .C1(new_n1193), .C2(new_n474), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1055), .A2(new_n1119), .A3(new_n1144), .A4(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1192), .A2(new_n1196), .A3(new_n1151), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(G171), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(KEYINPUT119), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1146), .A2(new_n1147), .A3(new_n1142), .ZN(new_n1202));
  OAI211_X1 g777(.A(G301), .B(new_n1192), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1197), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1200), .A2(new_n1203), .A3(KEYINPUT54), .A4(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT54), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1208), .B1(new_n1155), .B2(G301), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1209), .A2(KEYINPUT123), .A3(new_n1200), .A4(new_n1204), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n1190), .A2(new_n1191), .A3(new_n1207), .A4(new_n1210), .ZN(new_n1211));
  XOR2_X1   g786(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n1212));
  NOR2_X1   g787(.A1(new_n1197), .A2(G171), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1212), .B1(new_n1156), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT121), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g791(.A(KEYINPUT121), .B(new_n1212), .C1(new_n1156), .C2(new_n1213), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1161), .B1(new_n1211), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT115), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1088), .A2(G8), .A3(G168), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1221), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1222), .A2(new_n1133), .A3(new_n1118), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1130), .A2(G8), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n1134), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1225), .A2(KEYINPUT63), .ZN(new_n1226));
  OAI21_X1  g801(.A(new_n1220), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT63), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1228), .B1(new_n1140), .B2(new_n1221), .ZN(new_n1229));
  AND2_X1   g804(.A1(new_n1118), .A2(new_n1133), .ZN(new_n1230));
  AOI21_X1  g805(.A(new_n1228), .B1(new_n1224), .B2(new_n1134), .ZN(new_n1231));
  NAND4_X1  g806(.A1(new_n1230), .A2(KEYINPUT115), .A3(new_n1222), .A4(new_n1231), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1227), .A2(new_n1229), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g808(.A(new_n1133), .ZN(new_n1234));
  AND2_X1   g809(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1235));
  OR2_X1    g810(.A1(G288), .A2(G1976), .ZN(new_n1236));
  OAI21_X1  g811(.A(new_n1103), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  AOI22_X1  g812(.A1(new_n1234), .A2(new_n1118), .B1(new_n1237), .B2(new_n1113), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1233), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g814(.A(new_n1070), .B1(new_n1219), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g815(.A(new_n1060), .ZN(new_n1241));
  OR3_X1    g816(.A1(new_n1064), .A2(new_n847), .A3(new_n844), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n803), .A2(new_n805), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n1241), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g819(.A(KEYINPUT124), .ZN(new_n1245));
  INV_X1    g820(.A(KEYINPUT46), .ZN(new_n1246));
  OAI22_X1  g821(.A1(new_n1241), .A2(G1996), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n1063), .A2(new_n782), .ZN(new_n1248));
  AOI22_X1  g823(.A1(new_n1060), .A2(new_n1248), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1249));
  NAND4_X1  g824(.A1(new_n1060), .A2(KEYINPUT124), .A3(KEYINPUT46), .A4(new_n1061), .ZN(new_n1250));
  NAND3_X1  g825(.A1(new_n1247), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  XOR2_X1   g826(.A(new_n1251), .B(KEYINPUT47), .Z(new_n1252));
  NAND2_X1  g827(.A1(new_n1066), .A2(new_n1060), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1060), .A2(new_n1069), .ZN(new_n1254));
  XNOR2_X1  g829(.A(new_n1254), .B(KEYINPUT48), .ZN(new_n1255));
  AOI211_X1 g830(.A(new_n1244), .B(new_n1252), .C1(new_n1253), .C2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1240), .A2(new_n1256), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1259));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1260));
  NAND3_X1  g834(.A1(new_n741), .A2(new_n746), .A3(new_n701), .ZN(new_n1261));
  OAI21_X1  g835(.A(G319), .B1(new_n681), .B2(new_n685), .ZN(new_n1262));
  INV_X1    g836(.A(KEYINPUT125), .ZN(new_n1263));
  NOR3_X1   g837(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g838(.A(new_n1264), .B1(new_n980), .B2(new_n981), .ZN(new_n1265));
  OAI21_X1  g839(.A(new_n1263), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1266));
  AND4_X1   g840(.A1(new_n1260), .A2(new_n1043), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  INV_X1    g841(.A(new_n1266), .ZN(new_n1268));
  AOI21_X1  g842(.A(new_n1268), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1269));
  AOI21_X1  g843(.A(new_n1260), .B1(new_n1269), .B2(new_n1265), .ZN(new_n1270));
  OAI21_X1  g844(.A(new_n1259), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g845(.A1(new_n1043), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1272));
  NAND2_X1  g846(.A1(new_n1272), .A2(KEYINPUT126), .ZN(new_n1273));
  NAND3_X1  g847(.A1(new_n1269), .A2(new_n1260), .A3(new_n1265), .ZN(new_n1274));
  NAND3_X1  g848(.A1(new_n1273), .A2(KEYINPUT127), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g849(.A1(new_n1271), .A2(new_n1275), .ZN(G308));
  NAND2_X1  g850(.A1(new_n1273), .A2(new_n1274), .ZN(G225));
endmodule


