

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U551 ( .A1(n770), .A2(n772), .ZN(n725) );
  BUF_X1 U552 ( .A(n561), .Z(n540) );
  AND2_X1 U553 ( .A1(n772), .A2(n770), .ZN(n718) );
  NOR2_X1 U554 ( .A1(G2105), .A2(n539), .ZN(n561) );
  BUF_X1 U555 ( .A(n563), .Z(n891) );
  XOR2_X1 U556 ( .A(n698), .B(KEYINPUT28), .Z(n516) );
  OR2_X1 U557 ( .A1(n710), .A2(n709), .ZN(n517) );
  AND2_X1 U558 ( .A1(n712), .A2(n995), .ZN(n518) );
  XOR2_X1 U559 ( .A(G543), .B(KEYINPUT0), .Z(n519) );
  NOR2_X1 U560 ( .A1(n697), .A2(n696), .ZN(n712) );
  OR2_X1 U561 ( .A1(n751), .A2(n727), .ZN(n728) );
  NOR2_X1 U562 ( .A1(n713), .A2(n518), .ZN(n714) );
  INV_X1 U563 ( .A(KEYINPUT29), .ZN(n716) );
  INV_X1 U564 ( .A(KEYINPUT31), .ZN(n734) );
  INV_X1 U565 ( .A(KEYINPUT88), .ZN(n693) );
  INV_X1 U566 ( .A(n1007), .ZN(n761) );
  BUF_X1 U567 ( .A(n724), .Z(n739) );
  NOR2_X1 U568 ( .A1(n739), .A2(n764), .ZN(n765) );
  XNOR2_X1 U569 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n534) );
  NOR2_X1 U570 ( .A1(n765), .A2(KEYINPUT33), .ZN(n766) );
  XNOR2_X1 U571 ( .A(n541), .B(KEYINPUT65), .ZN(n563) );
  NOR2_X1 U572 ( .A1(n643), .A2(n525), .ZN(n659) );
  INV_X1 U573 ( .A(KEYINPUT87), .ZN(n535) );
  XNOR2_X1 U574 ( .A(n536), .B(n535), .ZN(n538) );
  NOR2_X1 U575 ( .A1(G651), .A2(G543), .ZN(n655) );
  NAND2_X1 U576 ( .A1(n655), .A2(G89), .ZN(n520) );
  XNOR2_X1 U577 ( .A(n520), .B(KEYINPUT4), .ZN(n522) );
  XNOR2_X1 U578 ( .A(KEYINPUT68), .B(n519), .ZN(n643) );
  XNOR2_X1 U579 ( .A(G651), .B(KEYINPUT69), .ZN(n525) );
  NAND2_X1 U580 ( .A1(G76), .A2(n659), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U582 ( .A(KEYINPUT5), .B(n523), .ZN(n531) );
  NOR2_X2 U583 ( .A1(G651), .A2(n643), .ZN(n656) );
  NAND2_X1 U584 ( .A1(n656), .A2(G51), .ZN(n524) );
  XOR2_X1 U585 ( .A(KEYINPUT79), .B(n524), .Z(n528) );
  NOR2_X1 U586 ( .A1(G543), .A2(n525), .ZN(n526) );
  XOR2_X2 U587 ( .A(KEYINPUT1), .B(n526), .Z(n663) );
  NAND2_X1 U588 ( .A1(G63), .A2(n663), .ZN(n527) );
  NAND2_X1 U589 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U590 ( .A(KEYINPUT6), .B(n529), .Z(n530) );
  NAND2_X1 U591 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U592 ( .A(KEYINPUT7), .B(n532), .ZN(G168) );
  XOR2_X1 U593 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U594 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  XNOR2_X2 U595 ( .A(n534), .B(n533), .ZN(n895) );
  NAND2_X1 U596 ( .A1(G138), .A2(n895), .ZN(n536) );
  AND2_X1 U597 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  NAND2_X1 U598 ( .A1(n892), .A2(G114), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n545) );
  INV_X1 U600 ( .A(G2104), .ZN(n539) );
  NAND2_X1 U601 ( .A1(G102), .A2(n540), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n539), .A2(G2105), .ZN(n541) );
  NAND2_X1 U603 ( .A1(G126), .A2(n891), .ZN(n542) );
  NAND2_X1 U604 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U605 ( .A1(n545), .A2(n544), .ZN(G164) );
  XOR2_X1 U606 ( .A(G2443), .B(G2446), .Z(n547) );
  XNOR2_X1 U607 ( .A(G2427), .B(G2451), .ZN(n546) );
  XNOR2_X1 U608 ( .A(n547), .B(n546), .ZN(n553) );
  XOR2_X1 U609 ( .A(G2430), .B(G2454), .Z(n549) );
  XNOR2_X1 U610 ( .A(G1341), .B(G1348), .ZN(n548) );
  XNOR2_X1 U611 ( .A(n549), .B(n548), .ZN(n551) );
  XOR2_X1 U612 ( .A(G2435), .B(G2438), .Z(n550) );
  XNOR2_X1 U613 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U614 ( .A(n553), .B(n552), .Z(n554) );
  AND2_X1 U615 ( .A1(G14), .A2(n554), .ZN(G401) );
  NAND2_X1 U616 ( .A1(n655), .A2(G85), .ZN(n556) );
  NAND2_X1 U617 ( .A1(G72), .A2(n659), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n656), .A2(G47), .ZN(n558) );
  NAND2_X1 U620 ( .A1(G60), .A2(n663), .ZN(n557) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  OR2_X1 U622 ( .A1(n560), .A2(n559), .ZN(G290) );
  NAND2_X1 U623 ( .A1(n561), .A2(G101), .ZN(n562) );
  XOR2_X1 U624 ( .A(KEYINPUT23), .B(n562), .Z(n565) );
  NAND2_X1 U625 ( .A1(n563), .A2(G125), .ZN(n564) );
  NAND2_X1 U626 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U627 ( .A(n566), .B(KEYINPUT66), .ZN(n570) );
  NAND2_X1 U628 ( .A1(n895), .A2(G137), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n892), .A2(G113), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U632 ( .A(n571), .B(KEYINPUT64), .ZN(n692) );
  BUF_X1 U633 ( .A(n692), .Z(G160) );
  NAND2_X1 U634 ( .A1(n656), .A2(G52), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G64), .A2(n663), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n655), .A2(G90), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G77), .A2(n659), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U640 ( .A(KEYINPUT9), .B(n577), .Z(n578) );
  NOR2_X1 U641 ( .A1(n579), .A2(n578), .ZN(G171) );
  AND2_X1 U642 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U643 ( .A(G132), .ZN(G219) );
  INV_X1 U644 ( .A(G82), .ZN(G220) );
  NAND2_X1 U645 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n580), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U647 ( .A(G223), .ZN(n837) );
  NAND2_X1 U648 ( .A1(n837), .A2(G567), .ZN(n581) );
  XOR2_X1 U649 ( .A(KEYINPUT11), .B(n581), .Z(G234) );
  NAND2_X1 U650 ( .A1(G56), .A2(n663), .ZN(n582) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(n582), .Z(n588) );
  NAND2_X1 U652 ( .A1(n655), .A2(G81), .ZN(n583) );
  XNOR2_X1 U653 ( .A(n583), .B(KEYINPUT12), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G68), .A2(n659), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U656 ( .A(KEYINPUT13), .B(n586), .Z(n587) );
  NOR2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U658 ( .A(n589), .B(KEYINPUT74), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G43), .A2(n656), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n998) );
  INV_X1 U661 ( .A(G860), .ZN(n615) );
  OR2_X1 U662 ( .A1(n998), .A2(n615), .ZN(n592) );
  XOR2_X1 U663 ( .A(KEYINPUT75), .B(n592), .Z(G153) );
  INV_X1 U664 ( .A(G171), .ZN(G301) );
  NAND2_X1 U665 ( .A1(n663), .A2(G66), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT76), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n655), .A2(G92), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G79), .A2(n659), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U670 ( .A1(G54), .A2(n656), .ZN(n596) );
  XNOR2_X1 U671 ( .A(KEYINPUT77), .B(n596), .ZN(n597) );
  NOR2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U674 ( .A(KEYINPUT15), .B(n601), .Z(n1002) );
  INV_X1 U675 ( .A(G868), .ZN(n674) );
  NAND2_X1 U676 ( .A1(n1002), .A2(n674), .ZN(n602) );
  XNOR2_X1 U677 ( .A(n602), .B(KEYINPUT78), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n604), .A2(n603), .ZN(G284) );
  NAND2_X1 U680 ( .A1(n656), .A2(G53), .ZN(n606) );
  NAND2_X1 U681 ( .A1(G65), .A2(n663), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n655), .A2(G91), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n607), .B(KEYINPUT70), .ZN(n609) );
  NAND2_X1 U685 ( .A1(G78), .A2(n659), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U687 ( .A(KEYINPUT71), .B(n610), .Z(n611) );
  NOR2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n995) );
  XOR2_X1 U689 ( .A(n995), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U690 ( .A1(G299), .A2(G868), .ZN(n614) );
  NOR2_X1 U691 ( .A1(G286), .A2(n674), .ZN(n613) );
  NOR2_X1 U692 ( .A1(n614), .A2(n613), .ZN(G297) );
  NAND2_X1 U693 ( .A1(n615), .A2(G559), .ZN(n616) );
  INV_X1 U694 ( .A(n1002), .ZN(n638) );
  NAND2_X1 U695 ( .A1(n616), .A2(n638), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n617), .B(KEYINPUT80), .ZN(n619) );
  XOR2_X1 U697 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n618) );
  XNOR2_X1 U698 ( .A(n619), .B(n618), .ZN(G148) );
  NOR2_X1 U699 ( .A1(G868), .A2(n998), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G868), .A2(n638), .ZN(n620) );
  NOR2_X1 U701 ( .A1(G559), .A2(n620), .ZN(n621) );
  NOR2_X1 U702 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U703 ( .A1(G99), .A2(n540), .ZN(n624) );
  NAND2_X1 U704 ( .A1(G111), .A2(n892), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n891), .A2(G123), .ZN(n625) );
  XNOR2_X1 U707 ( .A(n625), .B(KEYINPUT18), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G135), .A2(n895), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n977) );
  XNOR2_X1 U711 ( .A(n977), .B(G2096), .ZN(n631) );
  INV_X1 U712 ( .A(G2100), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n631), .A2(n630), .ZN(G156) );
  NAND2_X1 U714 ( .A1(n655), .A2(G93), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G80), .A2(n659), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n656), .A2(G55), .ZN(n635) );
  NAND2_X1 U718 ( .A1(G67), .A2(n663), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n636) );
  OR2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n675) );
  XNOR2_X1 U721 ( .A(n998), .B(KEYINPUT82), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n638), .A2(G559), .ZN(n639) );
  XNOR2_X1 U723 ( .A(n640), .B(n639), .ZN(n672) );
  NOR2_X1 U724 ( .A1(n672), .A2(G860), .ZN(n641) );
  XOR2_X1 U725 ( .A(KEYINPUT83), .B(n641), .Z(n642) );
  XOR2_X1 U726 ( .A(n675), .B(n642), .Z(G145) );
  NAND2_X1 U727 ( .A1(G49), .A2(n656), .ZN(n645) );
  NAND2_X1 U728 ( .A1(G87), .A2(n643), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U730 ( .A1(n663), .A2(n646), .ZN(n648) );
  NAND2_X1 U731 ( .A1(G651), .A2(G74), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n648), .A2(n647), .ZN(G288) );
  NAND2_X1 U733 ( .A1(G88), .A2(n655), .ZN(n650) );
  NAND2_X1 U734 ( .A1(G50), .A2(n656), .ZN(n649) );
  NAND2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U736 ( .A1(G75), .A2(n659), .ZN(n652) );
  NAND2_X1 U737 ( .A1(G62), .A2(n663), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U739 ( .A1(n654), .A2(n653), .ZN(G166) );
  NAND2_X1 U740 ( .A1(G86), .A2(n655), .ZN(n658) );
  NAND2_X1 U741 ( .A1(G48), .A2(n656), .ZN(n657) );
  NAND2_X1 U742 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n659), .A2(G73), .ZN(n660) );
  XOR2_X1 U744 ( .A(KEYINPUT2), .B(n660), .Z(n661) );
  NOR2_X1 U745 ( .A1(n662), .A2(n661), .ZN(n665) );
  NAND2_X1 U746 ( .A1(G61), .A2(n663), .ZN(n664) );
  NAND2_X1 U747 ( .A1(n665), .A2(n664), .ZN(G305) );
  XNOR2_X1 U748 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n666) );
  XOR2_X1 U749 ( .A(n666), .B(n675), .Z(n667) );
  XNOR2_X1 U750 ( .A(n667), .B(G288), .ZN(n670) );
  XNOR2_X1 U751 ( .A(G166), .B(G299), .ZN(n668) );
  XNOR2_X1 U752 ( .A(n668), .B(G290), .ZN(n669) );
  XNOR2_X1 U753 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U754 ( .A(n671), .B(G305), .ZN(n906) );
  XOR2_X1 U755 ( .A(n906), .B(n672), .Z(n673) );
  NOR2_X1 U756 ( .A1(n674), .A2(n673), .ZN(n677) );
  NOR2_X1 U757 ( .A1(G868), .A2(n675), .ZN(n676) );
  NOR2_X1 U758 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U759 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XOR2_X1 U760 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U761 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U762 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U763 ( .A1(n681), .A2(G2072), .ZN(n682) );
  XOR2_X1 U764 ( .A(KEYINPUT85), .B(n682), .Z(G158) );
  XNOR2_X1 U765 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  XNOR2_X1 U766 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n690) );
  NAND2_X1 U768 ( .A1(G108), .A2(G120), .ZN(n683) );
  NOR2_X1 U769 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U770 ( .A1(G69), .A2(n684), .ZN(n842) );
  NAND2_X1 U771 ( .A1(n842), .A2(G567), .ZN(n689) );
  NOR2_X1 U772 ( .A1(G220), .A2(G219), .ZN(n685) );
  XOR2_X1 U773 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U774 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U775 ( .A1(G96), .A2(n687), .ZN(n843) );
  NAND2_X1 U776 ( .A1(n843), .A2(G2106), .ZN(n688) );
  NAND2_X1 U777 ( .A1(n689), .A2(n688), .ZN(n844) );
  NOR2_X1 U778 ( .A1(n690), .A2(n844), .ZN(n691) );
  XNOR2_X1 U779 ( .A(n691), .B(KEYINPUT86), .ZN(n840) );
  NAND2_X1 U780 ( .A1(G36), .A2(n840), .ZN(G176) );
  INV_X1 U781 ( .A(G166), .ZN(G303) );
  NAND2_X1 U782 ( .A1(n692), .A2(G40), .ZN(n694) );
  XNOR2_X2 U783 ( .A(n694), .B(n693), .ZN(n770) );
  NOR2_X1 U784 ( .A1(G164), .A2(G1384), .ZN(n772) );
  NAND2_X1 U785 ( .A1(G8), .A2(n725), .ZN(n724) );
  NAND2_X1 U786 ( .A1(n718), .A2(G2072), .ZN(n695) );
  XNOR2_X1 U787 ( .A(n695), .B(KEYINPUT27), .ZN(n697) );
  XOR2_X1 U788 ( .A(G1956), .B(KEYINPUT96), .Z(n927) );
  NOR2_X1 U789 ( .A1(n718), .A2(n927), .ZN(n696) );
  NOR2_X1 U790 ( .A1(n712), .A2(n995), .ZN(n698) );
  NAND2_X1 U791 ( .A1(G1348), .A2(n725), .ZN(n700) );
  NAND2_X1 U792 ( .A1(G2067), .A2(n718), .ZN(n699) );
  NAND2_X1 U793 ( .A1(n700), .A2(n699), .ZN(n711) );
  NAND2_X1 U794 ( .A1(n1002), .A2(n711), .ZN(n703) );
  XOR2_X1 U795 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n705) );
  NOR2_X1 U796 ( .A1(G1996), .A2(n705), .ZN(n701) );
  NOR2_X1 U797 ( .A1(n998), .A2(n701), .ZN(n702) );
  NAND2_X1 U798 ( .A1(n703), .A2(n702), .ZN(n710) );
  INV_X1 U799 ( .A(G1341), .ZN(n999) );
  NAND2_X1 U800 ( .A1(n999), .A2(n705), .ZN(n704) );
  NAND2_X1 U801 ( .A1(n704), .A2(n725), .ZN(n708) );
  AND2_X1 U802 ( .A1(G1996), .A2(n718), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U804 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U805 ( .A1(n711), .A2(n1002), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n517), .A2(n714), .ZN(n715) );
  NAND2_X1 U807 ( .A1(n516), .A2(n715), .ZN(n717) );
  XNOR2_X1 U808 ( .A(n717), .B(n716), .ZN(n723) );
  XOR2_X1 U809 ( .A(G2078), .B(KEYINPUT25), .Z(n952) );
  NOR2_X1 U810 ( .A1(n952), .A2(n725), .ZN(n720) );
  NOR2_X1 U811 ( .A1(n718), .A2(G1961), .ZN(n719) );
  NOR2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U813 ( .A(KEYINPUT95), .B(n721), .ZN(n731) );
  NAND2_X1 U814 ( .A1(n731), .A2(G171), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n737) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n724), .ZN(n751) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n725), .ZN(n748) );
  INV_X1 U818 ( .A(n748), .ZN(n726) );
  NAND2_X1 U819 ( .A1(n726), .A2(G8), .ZN(n727) );
  XNOR2_X1 U820 ( .A(n728), .B(KEYINPUT30), .ZN(n729) );
  NOR2_X1 U821 ( .A1(n729), .A2(G168), .ZN(n730) );
  XNOR2_X1 U822 ( .A(n730), .B(KEYINPUT98), .ZN(n733) );
  NOR2_X1 U823 ( .A1(n731), .A2(G171), .ZN(n732) );
  NOR2_X1 U824 ( .A1(n733), .A2(n732), .ZN(n735) );
  XNOR2_X1 U825 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n749) );
  NAND2_X1 U827 ( .A1(n749), .A2(G286), .ZN(n744) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n725), .ZN(n738) );
  XOR2_X1 U829 ( .A(KEYINPUT99), .B(n738), .Z(n741) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n739), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U834 ( .A(n745), .B(KEYINPUT100), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n746), .A2(G8), .ZN(n747) );
  XNOR2_X1 U836 ( .A(n747), .B(KEYINPUT32), .ZN(n755) );
  NAND2_X1 U837 ( .A1(G8), .A2(n748), .ZN(n753) );
  INV_X1 U838 ( .A(n749), .ZN(n750) );
  NOR2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n811) );
  NOR2_X1 U842 ( .A1(G288), .A2(G1976), .ZN(n756) );
  XNOR2_X1 U843 ( .A(n756), .B(KEYINPUT101), .ZN(n767) );
  INV_X1 U844 ( .A(n767), .ZN(n758) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n757) );
  NOR2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n1006) );
  NAND2_X1 U847 ( .A1(n811), .A2(n1006), .ZN(n759) );
  XNOR2_X1 U848 ( .A(n759), .B(KEYINPUT102), .ZN(n762) );
  NAND2_X1 U849 ( .A1(G288), .A2(G1976), .ZN(n760) );
  XNOR2_X1 U850 ( .A(n760), .B(KEYINPUT103), .ZN(n1007) );
  NAND2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U852 ( .A(n763), .B(KEYINPUT104), .ZN(n764) );
  XNOR2_X1 U853 ( .A(n766), .B(KEYINPUT105), .ZN(n808) );
  XOR2_X1 U854 ( .A(G1981), .B(G305), .Z(n1014) );
  NOR2_X1 U855 ( .A1(n739), .A2(n767), .ZN(n768) );
  NAND2_X1 U856 ( .A1(KEYINPUT33), .A2(n768), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n1014), .A2(n769), .ZN(n806) );
  INV_X1 U858 ( .A(n770), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n771), .A2(n772), .ZN(n829) );
  XOR2_X1 U860 ( .A(KEYINPUT37), .B(G2067), .Z(n827) );
  XNOR2_X1 U861 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n783) );
  NAND2_X1 U862 ( .A1(G104), .A2(n540), .ZN(n774) );
  NAND2_X1 U863 ( .A1(G140), .A2(n895), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U865 ( .A(KEYINPUT34), .B(n775), .ZN(n780) );
  NAND2_X1 U866 ( .A1(G128), .A2(n891), .ZN(n777) );
  NAND2_X1 U867 ( .A1(G116), .A2(n892), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U869 ( .A(n778), .B(KEYINPUT35), .Z(n779) );
  NOR2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U871 ( .A(KEYINPUT36), .B(n781), .Z(n782) );
  XOR2_X1 U872 ( .A(n783), .B(n782), .Z(n888) );
  NAND2_X1 U873 ( .A1(n827), .A2(n888), .ZN(n784) );
  XNOR2_X1 U874 ( .A(KEYINPUT91), .B(n784), .ZN(n986) );
  NAND2_X1 U875 ( .A1(n829), .A2(n986), .ZN(n825) );
  XNOR2_X1 U876 ( .A(G1986), .B(G290), .ZN(n1004) );
  NAND2_X1 U877 ( .A1(n1004), .A2(n829), .ZN(n785) );
  AND2_X1 U878 ( .A1(n825), .A2(n785), .ZN(n805) );
  NAND2_X1 U879 ( .A1(G105), .A2(n540), .ZN(n786) );
  XNOR2_X1 U880 ( .A(n786), .B(KEYINPUT38), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G129), .A2(n891), .ZN(n788) );
  NAND2_X1 U882 ( .A1(G117), .A2(n892), .ZN(n787) );
  NAND2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U884 ( .A1(G141), .A2(n895), .ZN(n789) );
  XNOR2_X1 U885 ( .A(KEYINPUT93), .B(n789), .ZN(n790) );
  NOR2_X1 U886 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n878) );
  NAND2_X1 U888 ( .A1(G1996), .A2(n878), .ZN(n794) );
  XOR2_X1 U889 ( .A(KEYINPUT94), .B(n794), .Z(n803) );
  NAND2_X1 U890 ( .A1(G95), .A2(n540), .ZN(n796) );
  NAND2_X1 U891 ( .A1(G107), .A2(n892), .ZN(n795) );
  NAND2_X1 U892 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n891), .A2(G119), .ZN(n797) );
  XOR2_X1 U894 ( .A(KEYINPUT92), .B(n797), .Z(n798) );
  NOR2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U896 ( .A1(n895), .A2(G131), .ZN(n800) );
  NAND2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n883) );
  AND2_X1 U898 ( .A1(G1991), .A2(n883), .ZN(n802) );
  NOR2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n983) );
  INV_X1 U900 ( .A(n983), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n804), .A2(n829), .ZN(n819) );
  NAND2_X1 U902 ( .A1(n805), .A2(n819), .ZN(n818) );
  NOR2_X1 U903 ( .A1(n806), .A2(n818), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n834) );
  NOR2_X1 U905 ( .A1(G1981), .A2(G305), .ZN(n809) );
  XOR2_X1 U906 ( .A(n809), .B(KEYINPUT24), .Z(n810) );
  NOR2_X1 U907 ( .A1(n739), .A2(n810), .ZN(n816) );
  NOR2_X1 U908 ( .A1(G2090), .A2(G303), .ZN(n812) );
  NAND2_X1 U909 ( .A1(G8), .A2(n812), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n811), .A2(n813), .ZN(n814) );
  AND2_X1 U911 ( .A1(n814), .A2(n739), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n817) );
  OR2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n832) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n878), .ZN(n968) );
  INV_X1 U915 ( .A(n819), .ZN(n822) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U917 ( .A1(G1991), .A2(n883), .ZN(n978) );
  NOR2_X1 U918 ( .A1(n820), .A2(n978), .ZN(n821) );
  NOR2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U920 ( .A1(n968), .A2(n823), .ZN(n824) );
  XNOR2_X1 U921 ( .A(KEYINPUT39), .B(n824), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n828) );
  OR2_X1 U923 ( .A1(n888), .A2(n827), .ZN(n979) );
  NAND2_X1 U924 ( .A1(n828), .A2(n979), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  AND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(n836) );
  XNOR2_X1 U928 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n836), .B(n835), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U932 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U935 ( .A(KEYINPUT107), .B(n841), .Z(G188) );
  NOR2_X1 U936 ( .A1(n843), .A2(n842), .ZN(G325) );
  XOR2_X1 U937 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G108), .ZN(G238) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  INV_X1 U942 ( .A(G69), .ZN(G235) );
  INV_X1 U943 ( .A(n844), .ZN(G319) );
  XOR2_X1 U944 ( .A(G2100), .B(G2096), .Z(n846) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U950 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U951 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U953 ( .A(G1976), .B(G1981), .Z(n854) );
  XNOR2_X1 U954 ( .A(G1966), .B(G1956), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(n855), .B(G2474), .Z(n857) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1971), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U959 ( .A(KEYINPUT41), .B(G1961), .Z(n859) );
  XNOR2_X1 U960 ( .A(G1996), .B(G1991), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(G229) );
  NAND2_X1 U963 ( .A1(G100), .A2(n540), .ZN(n863) );
  NAND2_X1 U964 ( .A1(G112), .A2(n892), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U966 ( .A1(G124), .A2(n891), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n864), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G136), .A2(n895), .ZN(n865) );
  XOR2_X1 U969 ( .A(KEYINPUT109), .B(n865), .Z(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U971 ( .A1(n869), .A2(n868), .ZN(G162) );
  NAND2_X1 U972 ( .A1(G103), .A2(n540), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G139), .A2(n895), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G127), .A2(n891), .ZN(n873) );
  NAND2_X1 U976 ( .A1(G115), .A2(n892), .ZN(n872) );
  NAND2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U978 ( .A(KEYINPUT47), .B(n874), .ZN(n875) );
  XNOR2_X1 U979 ( .A(KEYINPUT111), .B(n875), .ZN(n876) );
  NOR2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n970) );
  XNOR2_X1 U981 ( .A(n970), .B(G160), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n879), .B(n878), .ZN(n887) );
  XOR2_X1 U983 ( .A(KEYINPUT113), .B(KEYINPUT48), .Z(n881) );
  XNOR2_X1 U984 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U985 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U986 ( .A(n882), .B(KEYINPUT112), .Z(n885) );
  XOR2_X1 U987 ( .A(n883), .B(n977), .Z(n884) );
  XNOR2_X1 U988 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U989 ( .A(n887), .B(n886), .Z(n890) );
  XOR2_X1 U990 ( .A(G164), .B(n888), .Z(n889) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n904) );
  NAND2_X1 U992 ( .A1(G130), .A2(n891), .ZN(n894) );
  NAND2_X1 U993 ( .A1(G118), .A2(n892), .ZN(n893) );
  NAND2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n901) );
  NAND2_X1 U995 ( .A1(G106), .A2(n540), .ZN(n897) );
  NAND2_X1 U996 ( .A1(G142), .A2(n895), .ZN(n896) );
  NAND2_X1 U997 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U998 ( .A(KEYINPUT110), .B(n898), .Z(n899) );
  XNOR2_X1 U999 ( .A(KEYINPUT45), .B(n899), .ZN(n900) );
  NOR2_X1 U1000 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1001 ( .A(G162), .B(n902), .Z(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(G286), .B(n906), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(KEYINPUT115), .B(G301), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n907), .B(n1002), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1008 ( .A(n910), .B(n998), .Z(n911) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n911), .ZN(G397) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n913), .B(n912), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(KEYINPUT117), .B(n914), .ZN(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n917), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(n918), .A2(G401), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(n919), .B(KEYINPUT118), .ZN(G308) );
  INV_X1 U1019 ( .A(G308), .ZN(G225) );
  XNOR2_X1 U1020 ( .A(G1966), .B(G21), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(G5), .B(G1961), .ZN(n920) );
  NOR2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n934) );
  XOR2_X1 U1023 ( .A(G1981), .B(G6), .Z(n926) );
  XOR2_X1 U1024 ( .A(KEYINPUT126), .B(G4), .Z(n923) );
  XNOR2_X1 U1025 ( .A(G1348), .B(KEYINPUT59), .ZN(n922) );
  XNOR2_X1 U1026 ( .A(n923), .B(n922), .ZN(n924) );
  XNOR2_X1 U1027 ( .A(KEYINPUT125), .B(n924), .ZN(n925) );
  NAND2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n927), .B(G20), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n999), .B(G19), .ZN(n928) );
  NAND2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(n932), .B(KEYINPUT60), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n942) );
  XNOR2_X1 U1035 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n940) );
  XOR2_X1 U1036 ( .A(G1986), .B(G24), .Z(n938) );
  XNOR2_X1 U1037 ( .A(G1971), .B(G22), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(G23), .B(G1976), .ZN(n935) );
  NOR2_X1 U1039 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1040 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1041 ( .A(n940), .B(n939), .Z(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(KEYINPUT61), .B(n943), .ZN(n945) );
  INV_X1 U1044 ( .A(G16), .ZN(n944) );
  NAND2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n946), .A2(G11), .ZN(n994) );
  XNOR2_X1 U1047 ( .A(G2067), .B(G26), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(G2072), .B(G33), .ZN(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1050 ( .A(n949), .B(KEYINPUT120), .ZN(n951) );
  XOR2_X1 U1051 ( .A(G1991), .B(G25), .Z(n950) );
  NAND2_X1 U1052 ( .A1(n951), .A2(n950), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(G1996), .B(G32), .ZN(n954) );
  XNOR2_X1 U1054 ( .A(n952), .B(G27), .ZN(n953) );
  NOR2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1056 ( .A(n955), .B(KEYINPUT121), .ZN(n956) );
  NOR2_X1 U1057 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1058 ( .A1(G28), .A2(n958), .ZN(n959) );
  XNOR2_X1 U1059 ( .A(n959), .B(KEYINPUT53), .ZN(n962) );
  XOR2_X1 U1060 ( .A(G2084), .B(KEYINPUT54), .Z(n960) );
  XNOR2_X1 U1061 ( .A(G34), .B(n960), .ZN(n961) );
  NAND2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n964) );
  XNOR2_X1 U1063 ( .A(G35), .B(G2090), .ZN(n963) );
  NOR2_X1 U1064 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1065 ( .A1(G29), .A2(n965), .ZN(n966) );
  XNOR2_X1 U1066 ( .A(n966), .B(KEYINPUT55), .ZN(n992) );
  XOR2_X1 U1067 ( .A(G2090), .B(G162), .Z(n967) );
  NOR2_X1 U1068 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1069 ( .A(KEYINPUT51), .B(n969), .Z(n976) );
  XNOR2_X1 U1070 ( .A(KEYINPUT50), .B(KEYINPUT119), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(G2072), .B(n970), .ZN(n972) );
  XNOR2_X1 U1072 ( .A(G164), .B(G2078), .ZN(n971) );
  NAND2_X1 U1073 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1074 ( .A(n974), .B(n973), .ZN(n975) );
  NAND2_X1 U1075 ( .A1(n976), .A2(n975), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n980) );
  NAND2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(G2084), .B(G160), .ZN(n984) );
  NAND2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(KEYINPUT52), .B(n989), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(G29), .A2(n990), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n1024) );
  XNOR2_X1 U1087 ( .A(n995), .B(G1956), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(G171), .B(G1961), .ZN(n996) );
  NAND2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n1001) );
  XOR2_X1 U1090 ( .A(n999), .B(n998), .Z(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1019) );
  XNOR2_X1 U1092 ( .A(G1348), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1011) );
  NAND2_X1 U1094 ( .A1(G1971), .A2(G303), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(KEYINPUT123), .B(n1009), .Z(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(G1966), .B(G168), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(n1012), .B(KEYINPUT122), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT57), .B(n1015), .Z(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(KEYINPUT56), .B(G16), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(n1022), .B(KEYINPUT124), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

