//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n450, new_n452, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n635, new_n636, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT69), .Z(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n460), .A2(KEYINPUT70), .B1(new_n449), .B2(new_n456), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(KEYINPUT70), .B2(new_n460), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT71), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT74), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT73), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT73), .B1(new_n470), .B2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(KEYINPUT74), .A3(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n469), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n466), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n470), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT72), .ZN(new_n484));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G125), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n472), .B1(new_n486), .B2(new_n477), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n476), .B1(new_n484), .B2(new_n489), .ZN(G160));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT74), .A2(G2104), .ZN(new_n493));
  AOI22_X1  g068(.A1(KEYINPUT73), .A2(new_n478), .B1(new_n493), .B2(new_n470), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(G2105), .A3(new_n469), .ZN(new_n495));
  INV_X1    g070(.A(G124), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n474), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(G136), .B2(new_n498), .ZN(G162));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n474), .B2(new_n500), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n500), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n485), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT77), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n485), .A2(KEYINPUT77), .A3(new_n502), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n501), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(G114), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G2105), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(G126), .A2(G2105), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n469), .A2(new_n471), .A3(new_n473), .A4(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n514), .A2(KEYINPUT75), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(KEYINPUT75), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT76), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n494), .A2(new_n520), .A3(new_n469), .A4(new_n513), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n514), .A2(KEYINPUT75), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n511), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT76), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n508), .B1(new_n519), .B2(new_n524), .ZN(G164));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT79), .B1(new_n526), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT79), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT5), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n527), .A2(new_n530), .B1(new_n526), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT78), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT6), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(G651), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(KEYINPUT78), .A3(KEYINPUT6), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n534), .A2(new_n536), .B1(new_n533), .B2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G88), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G50), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n538), .A2(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n531), .A2(G62), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT80), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n543), .A2(new_n544), .B1(G75), .B2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n545), .B1(new_n544), .B2(new_n543), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n542), .B1(new_n546), .B2(G651), .ZN(G166));
  NAND3_X1  g122(.A1(new_n531), .A2(G63), .A3(G651), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT81), .ZN(new_n549));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT7), .ZN(new_n551));
  INV_X1    g126(.A(G51), .ZN(new_n552));
  INV_X1    g127(.A(G89), .ZN(new_n553));
  OAI221_X1 g128(.A(new_n551), .B1(new_n540), .B2(new_n552), .C1(new_n553), .C2(new_n538), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n549), .A2(new_n554), .ZN(G168));
  AOI22_X1  g130(.A1(new_n531), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n535), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  INV_X1    g133(.A(G52), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n538), .A2(new_n558), .B1(new_n540), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(G171));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n527), .A2(new_n530), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n526), .A2(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G56), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT82), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n535), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n569), .B1(new_n568), .B2(new_n567), .ZN(new_n570));
  INV_X1    g145(.A(new_n538), .ZN(new_n571));
  INV_X1    g146(.A(new_n540), .ZN(new_n572));
  AOI22_X1  g147(.A1(G81), .A2(new_n571), .B1(new_n572), .B2(G43), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(G860), .A3(new_n573), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n574), .B(KEYINPUT83), .Z(G153));
  NAND4_X1  g150(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g151(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n577));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(G319), .A2(G483), .A3(G661), .A4(new_n579), .ZN(G188));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n572), .A2(new_n581), .A3(G53), .ZN(new_n582));
  INV_X1    g157(.A(G53), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT9), .B1(new_n540), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT85), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n582), .A2(new_n587), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G78), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G65), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n565), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT86), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT86), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n594), .B(new_n590), .C1(new_n565), .C2(new_n591), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n593), .A2(new_n595), .A3(KEYINPUT87), .A4(G651), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n571), .A2(G91), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n593), .A2(new_n595), .A3(G651), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n589), .A2(new_n596), .A3(new_n597), .A4(new_n600), .ZN(G299));
  NOR2_X1   g176(.A1(G171), .A2(KEYINPUT88), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n603));
  NOR3_X1   g178(.A1(new_n557), .A2(new_n560), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n602), .A2(new_n604), .ZN(G301));
  INV_X1    g180(.A(G168), .ZN(G286));
  INV_X1    g181(.A(G166), .ZN(G303));
  NAND2_X1  g182(.A1(new_n571), .A2(G87), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n572), .A2(G49), .ZN(new_n609));
  OAI21_X1  g184(.A(G651), .B1(new_n531), .B2(G74), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(G288));
  NAND3_X1  g186(.A1(new_n537), .A2(G48), .A3(G543), .ZN(new_n612));
  INV_X1    g187(.A(G86), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n538), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n531), .A2(G61), .ZN(new_n616));
  NAND2_X1  g191(.A1(G73), .A2(G543), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n535), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n619), .ZN(G305));
  AOI22_X1  g195(.A1(G85), .A2(new_n571), .B1(new_n572), .B2(G47), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n531), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n535), .B2(new_n622), .ZN(G290));
  NAND2_X1  g198(.A1(new_n571), .A2(G92), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(G79), .A2(G543), .ZN(new_n627));
  INV_X1    g202(.A(G66), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n565), .B2(new_n628), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n629), .A2(G651), .B1(new_n572), .B2(G54), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  MUX2_X1   g206(.A(new_n631), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g207(.A(new_n631), .B(G301), .S(G868), .Z(G321));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NOR2_X1   g209(.A1(G286), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G299), .B(KEYINPUT89), .Z(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n634), .ZN(G280));
  XOR2_X1   g212(.A(G280), .B(KEYINPUT90), .Z(G297));
  INV_X1    g213(.A(new_n631), .ZN(new_n639));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G860), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT91), .Z(G148));
  NAND2_X1  g217(.A1(new_n570), .A2(new_n573), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(new_n634), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n631), .A2(G559), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(new_n634), .ZN(G323));
  XNOR2_X1  g221(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n647));
  XNOR2_X1  g222(.A(G323), .B(new_n647), .ZN(G282));
  NAND2_X1  g223(.A1(new_n485), .A2(new_n465), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT12), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT13), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(new_n652));
  OR2_X1    g227(.A1(G99), .A2(G2105), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n653), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n654));
  INV_X1    g229(.A(G123), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n495), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(G135), .B2(new_n498), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n658), .A2(G2096), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(G2096), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n652), .A2(new_n659), .A3(new_n660), .ZN(G156));
  INV_X1    g236(.A(KEYINPUT14), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2427), .B(G2438), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2430), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2451), .B(G2454), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1341), .B(G1348), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n667), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2443), .B(G2446), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  AND3_X1   g250(.A1(new_n674), .A2(G14), .A3(new_n675), .ZN(G401));
  XOR2_X1   g251(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(KEYINPUT17), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2072), .B(G2078), .Z(new_n684));
  INV_X1    g259(.A(new_n677), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2096), .B(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1961), .B(G1966), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(new_n694), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT20), .Z(new_n698));
  AOI211_X1 g273(.A(new_n696), .B(new_n698), .C1(new_n691), .C2(new_n695), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(G229));
  MUX2_X1   g280(.A(G6), .B(G305), .S(G16), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT32), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1981), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G22), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G166), .B2(G16), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(G1971), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n710), .A2(G1971), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G23), .ZN(new_n714));
  INV_X1    g289(.A(G288), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n716), .B(new_n717), .Z(new_n718));
  NOR4_X1   g293(.A1(new_n708), .A2(new_n711), .A3(new_n712), .A4(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  MUX2_X1   g297(.A(G24), .B(G290), .S(G16), .Z(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G1986), .Z(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G25), .ZN(new_n726));
  INV_X1    g301(.A(G119), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n472), .A2(G107), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n495), .A2(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n498), .A2(G131), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n726), .B1(new_n732), .B2(new_n725), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT95), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT94), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n733), .B(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n724), .B1(KEYINPUT96), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(KEYINPUT96), .B2(new_n737), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n721), .A2(new_n722), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT36), .ZN(new_n741));
  INV_X1    g316(.A(G34), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(KEYINPUT24), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n742), .B2(KEYINPUT24), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(KEYINPUT98), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(KEYINPUT98), .B2(new_n744), .ZN(new_n746));
  INV_X1    g321(.A(G160), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(new_n725), .ZN(new_n748));
  INV_X1    g323(.A(G2084), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n725), .A2(G32), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT26), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n754), .A2(new_n755), .B1(G105), .B2(new_n465), .ZN(new_n756));
  INV_X1    g331(.A(G129), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n495), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G141), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n474), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n751), .B1(new_n762), .B2(new_n725), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT27), .B(G1996), .Z(new_n764));
  AND2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G1961), .ZN(new_n766));
  NOR2_X1   g341(.A1(G171), .A2(new_n713), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G5), .B2(new_n713), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n750), .B(new_n765), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT102), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n713), .A2(G20), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT23), .ZN(new_n772));
  INV_X1    g347(.A(G299), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n713), .ZN(new_n774));
  INV_X1    g349(.A(G1956), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G29), .A2(G35), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G162), .B2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT29), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2090), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT25), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n782), .B1(new_n784), .B2(G2105), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n498), .A2(G139), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(new_n725), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n725), .B2(G33), .ZN(new_n789));
  INV_X1    g364(.A(G2072), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT31), .B(G11), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(G28), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT101), .Z(new_n795));
  OAI211_X1 g370(.A(new_n795), .B(new_n725), .C1(new_n793), .C2(G28), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n792), .B(new_n796), .C1(new_n658), .C2(new_n725), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n789), .B2(new_n790), .ZN(new_n798));
  NOR2_X1   g373(.A1(G16), .A2(G21), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G168), .B2(G16), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT100), .B(G1966), .Z(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n800), .A2(new_n802), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n791), .A2(new_n798), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n748), .A2(new_n749), .ZN(new_n806));
  OAI221_X1 g381(.A(new_n806), .B1(new_n768), .B2(new_n766), .C1(new_n763), .C2(new_n764), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n780), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n725), .A2(G27), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G164), .B2(new_n725), .ZN(new_n810));
  INV_X1    g385(.A(G2078), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n770), .A2(new_n776), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n713), .A2(G4), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n639), .B2(new_n713), .ZN(new_n815));
  INV_X1    g390(.A(G1348), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  MUX2_X1   g392(.A(G19), .B(new_n643), .S(G16), .Z(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(G1341), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n725), .A2(G26), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT28), .ZN(new_n821));
  INV_X1    g396(.A(G128), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n472), .A2(G116), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n495), .A2(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G140), .B2(new_n498), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n821), .B1(new_n826), .B2(new_n725), .ZN(new_n827));
  INV_X1    g402(.A(G2067), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n817), .A2(new_n819), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT97), .Z(new_n831));
  NOR2_X1   g406(.A1(new_n813), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n741), .A2(new_n832), .ZN(G150));
  INV_X1    g408(.A(G150), .ZN(G311));
  AOI22_X1  g409(.A1(new_n531), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(new_n535), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n571), .A2(G93), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n572), .A2(G55), .ZN(new_n838));
  AOI21_X1  g413(.A(KEYINPUT103), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  INV_X1    g415(.A(G55), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n538), .A2(new_n840), .B1(new_n540), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n836), .B1(new_n839), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT104), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n847), .B(new_n836), .C1(new_n839), .C2(new_n844), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n848), .A3(new_n643), .ZN(new_n849));
  INV_X1    g424(.A(new_n845), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n850), .A2(new_n847), .A3(new_n570), .A4(new_n573), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT38), .Z(new_n853));
  NOR2_X1   g428(.A1(new_n631), .A2(new_n640), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n856), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n845), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT37), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(G145));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n761), .B(new_n826), .ZN(new_n863));
  OR2_X1    g438(.A1(G106), .A2(G2105), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n864), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n865));
  INV_X1    g440(.A(G130), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n498), .A2(new_n867), .A3(G142), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n498), .B2(G142), .ZN(new_n869));
  OAI221_X1 g444(.A(new_n865), .B1(new_n866), .B2(new_n495), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n863), .B(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n732), .B(new_n650), .Z(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n507), .A2(new_n523), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n873), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n875), .B1(new_n874), .B2(new_n876), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n787), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT105), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(G162), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n747), .ZN(new_n884));
  INV_X1    g459(.A(new_n787), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n878), .B2(new_n879), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n884), .B1(new_n881), .B2(new_n886), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n862), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n892), .A2(KEYINPUT40), .A3(new_n888), .A4(new_n887), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n891), .A2(new_n893), .ZN(G395));
  XOR2_X1   g469(.A(new_n852), .B(new_n645), .Z(new_n895));
  NAND2_X1  g470(.A1(G299), .A2(new_n639), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n600), .A2(new_n596), .A3(new_n597), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n589), .A3(new_n631), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(KEYINPUT107), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n897), .A2(new_n902), .A3(new_n589), .A4(new_n631), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n896), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(G299), .B2(new_n639), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n904), .A2(new_n905), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n900), .B1(new_n907), .B2(new_n895), .ZN(new_n908));
  XOR2_X1   g483(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NAND2_X1  g486(.A1(G290), .A2(KEYINPUT108), .ZN(new_n912));
  OR2_X1    g487(.A1(G290), .A2(KEYINPUT108), .ZN(new_n913));
  NAND2_X1  g488(.A1(G166), .A2(KEYINPUT109), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(G166), .A2(KEYINPUT109), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n912), .B(new_n913), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(G290), .B(KEYINPUT108), .ZN(new_n918));
  INV_X1    g493(.A(new_n916), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n914), .ZN(new_n920));
  XNOR2_X1  g495(.A(G305), .B(G288), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n917), .B2(new_n920), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n910), .A2(new_n911), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n910), .B2(new_n911), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(G868), .B2(new_n850), .ZN(G295));
  OAI21_X1  g503(.A(new_n927), .B1(G868), .B2(new_n850), .ZN(G331));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n930));
  OAI21_X1  g505(.A(G168), .B1(new_n602), .B2(new_n604), .ZN(new_n931));
  OAI22_X1  g506(.A1(new_n549), .A2(new_n554), .B1(new_n557), .B2(new_n560), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n849), .A2(new_n851), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n851), .B2(new_n849), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n899), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n933), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n852), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n849), .A2(new_n851), .A3(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n924), .B(new_n936), .C1(new_n907), .C2(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n941), .A2(new_n888), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n899), .A2(new_n905), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n901), .A2(new_n903), .A3(new_n906), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n936), .B(new_n943), .C1(new_n940), .C2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n924), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(KEYINPUT112), .A3(new_n946), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n942), .A2(new_n949), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n904), .A2(new_n905), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n906), .A2(new_n898), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n939), .A3(new_n938), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n924), .B1(new_n956), .B2(new_n936), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n941), .A2(new_n888), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n930), .B1(new_n952), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n907), .A2(new_n940), .ZN(new_n961));
  INV_X1    g536(.A(new_n936), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n946), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n942), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT111), .B1(new_n964), .B2(KEYINPUT43), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n960), .A2(new_n965), .A3(KEYINPUT44), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n942), .A2(new_n949), .A3(new_n951), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT113), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n970), .A3(KEYINPUT43), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n942), .A2(new_n950), .A3(new_n963), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n966), .B1(KEYINPUT44), .B2(new_n973), .ZN(G397));
  AND2_X1   g549(.A1(KEYINPUT124), .A2(G8), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n484), .A2(new_n489), .ZN(new_n976));
  INV_X1    g551(.A(new_n476), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(G40), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n521), .A2(new_n522), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT76), .B1(new_n979), .B2(new_n512), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n518), .B(new_n511), .C1(new_n521), .C2(new_n522), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n507), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1384), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n978), .B1(new_n984), .B2(KEYINPUT50), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n875), .A2(new_n986), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT116), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n507), .B2(new_n523), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n990), .A3(new_n986), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n985), .A2(new_n749), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n982), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n994));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  AOI211_X1 g570(.A(new_n995), .B(new_n476), .C1(new_n484), .C2(new_n489), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n875), .A2(new_n983), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n994), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n801), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n993), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n975), .B1(new_n1002), .B2(G286), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT51), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1005), .B(new_n975), .C1(new_n1002), .C2(G286), .ZN(new_n1006));
  INV_X1    g581(.A(G8), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n993), .B2(new_n1001), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G286), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1004), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n992), .A2(new_n1012), .A3(new_n996), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n766), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n998), .B1(G164), .B2(G1384), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n978), .B1(KEYINPUT45), .B2(new_n989), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n811), .A3(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n875), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n811), .A2(KEYINPUT53), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n487), .A2(new_n995), .A3(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n999), .A2(new_n977), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1014), .A2(new_n1019), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G301), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n766), .A2(new_n1013), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1000), .A2(new_n1021), .ZN(new_n1028));
  AOI21_X1  g603(.A(G301), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1011), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G2090), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n985), .A2(new_n1031), .A3(new_n992), .ZN(new_n1032));
  INV_X1    g607(.A(G1971), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT45), .B1(new_n982), .B2(new_n983), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1020), .A2(new_n996), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1007), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(G166), .A2(new_n1007), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT55), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n982), .A2(new_n986), .A3(new_n983), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n978), .B1(new_n997), .B2(KEYINPUT50), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1042), .A3(new_n1031), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1007), .B1(new_n1036), .B2(new_n1043), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1044), .A2(new_n1039), .ZN(new_n1045));
  INV_X1    g620(.A(G1981), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n615), .A2(new_n619), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(G1981), .B1(new_n614), .B2(new_n618), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(KEYINPUT49), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT117), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1047), .A2(new_n1048), .A3(new_n1051), .A4(KEYINPUT49), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(G8), .B1(new_n997), .B2(new_n978), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT49), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1054), .ZN(new_n1058));
  INV_X1    g633(.A(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1058), .B(new_n1060), .C1(new_n1059), .C2(G288), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G288), .A2(new_n1059), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT52), .B1(new_n1054), .B2(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1057), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1040), .A2(new_n1045), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1024), .A2(G171), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1027), .A2(G301), .A3(new_n1028), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(KEYINPUT54), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1010), .A2(new_n1030), .A3(new_n1065), .A4(new_n1068), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT56), .B(G2072), .Z(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1015), .A2(new_n1016), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT120), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT57), .B1(new_n582), .B2(new_n584), .ZN(new_n1074));
  AOI22_X1  g649(.A1(G299), .A2(KEYINPUT57), .B1(new_n897), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n775), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1015), .A2(new_n1078), .A3(new_n1016), .A4(new_n1071), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT122), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1956), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1034), .A2(new_n1035), .A3(new_n1070), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(new_n1078), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n1075), .A4(new_n1073), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1075), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1035), .B1(new_n984), .B2(new_n998), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1078), .B1(new_n1089), .B2(new_n1071), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1087), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1081), .A2(KEYINPUT61), .A3(new_n1086), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1080), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT61), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n997), .A2(new_n978), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT58), .B(G1341), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1996), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n1089), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT59), .B1(new_n1099), .B2(new_n643), .ZN(new_n1100));
  OR3_X1    g675(.A1(new_n1099), .A2(KEYINPUT59), .A3(new_n643), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1093), .A2(new_n1094), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n639), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n639), .A2(new_n1104), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1013), .A2(new_n816), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n997), .A2(new_n978), .A3(G2067), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT121), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n1112), .B(new_n1109), .C1(new_n1013), .C2(new_n816), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1105), .B(new_n1107), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(G1348), .B1(new_n985), .B2(new_n992), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1112), .B1(new_n1115), .B2(new_n1109), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1108), .A2(KEYINPUT121), .A3(new_n1110), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n1103), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1107), .B1(new_n1120), .B2(new_n1105), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1092), .B(new_n1102), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1116), .A2(new_n1080), .A3(new_n1117), .A4(new_n639), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1091), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1069), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1064), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G288), .A2(G1976), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n1128), .B(KEYINPUT118), .Z(new_n1129));
  NAND2_X1  g704(.A1(new_n1057), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1054), .B1(new_n1130), .B2(new_n1047), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1040), .A2(new_n1045), .A3(new_n1064), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1008), .A2(G168), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1040), .A2(KEYINPUT63), .A3(G168), .A4(new_n1008), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1064), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT119), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1064), .B(new_n1141), .C1(new_n1037), .C2(new_n1039), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1138), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1132), .B1(new_n1137), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT126), .B1(new_n1126), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1132), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1138), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1146), .B1(new_n1149), .B2(new_n1136), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1101), .A2(new_n1100), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1092), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1105), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1106), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1156), .A2(new_n1118), .A3(new_n1114), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1124), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1150), .B(new_n1151), .C1(new_n1158), .C2(new_n1069), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1160), .A2(new_n1029), .A3(new_n1065), .A4(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1145), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n999), .A2(new_n978), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT114), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1165), .A2(new_n1098), .A3(new_n762), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT115), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1164), .A2(new_n1098), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1168), .A2(new_n761), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1165), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n826), .B(new_n828), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n732), .B(new_n735), .Z(new_n1174));
  AOI21_X1  g749(.A(new_n1173), .B1(new_n1174), .B2(new_n1170), .ZN(new_n1175));
  NOR2_X1   g750(.A1(G290), .A2(G1986), .ZN(new_n1176));
  AND2_X1   g751(.A1(G290), .A2(G1986), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1164), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1163), .A2(new_n1179), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n730), .A2(new_n731), .A3(new_n735), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1167), .A2(new_n1181), .A3(new_n1172), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n826), .A2(new_n828), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1165), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT46), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1168), .A2(new_n1185), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT127), .Z(new_n1187));
  NAND2_X1  g762(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1170), .A2(new_n761), .B1(new_n1185), .B2(new_n1168), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1190), .B(KEYINPUT47), .Z(new_n1191));
  NAND2_X1  g766(.A1(new_n1164), .A2(new_n1176), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT48), .ZN(new_n1193));
  AOI211_X1 g768(.A(new_n1184), .B(new_n1191), .C1(new_n1175), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1180), .A2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g770(.A1(new_n892), .A2(new_n888), .A3(new_n887), .ZN(new_n1197));
  INV_X1    g771(.A(G227), .ZN(new_n1198));
  NAND2_X1  g772(.A1(G319), .A2(new_n1198), .ZN(new_n1199));
  NOR3_X1   g773(.A1(G229), .A2(G401), .A3(new_n1199), .ZN(new_n1200));
  OAI211_X1 g774(.A(new_n1197), .B(new_n1200), .C1(new_n960), .C2(new_n965), .ZN(G225));
  INV_X1    g775(.A(G225), .ZN(G308));
endmodule


