//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G125), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G125), .B(G140), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(KEYINPUT16), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G125), .ZN(new_n194));
  INV_X1    g008(.A(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n189), .B1(new_n197), .B2(new_n187), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n193), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G128), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n204), .B(new_n206), .C1(G119), .C2(new_n205), .ZN(new_n207));
  XNOR2_X1  g021(.A(G119), .B(G128), .ZN(new_n208));
  XOR2_X1   g022(.A(KEYINPUT24), .B(G110), .Z(new_n209));
  AOI22_X1  g023(.A1(new_n207), .A2(G110), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n201), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n197), .A2(G146), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n212), .B1(new_n192), .B2(G146), .ZN(new_n213));
  XOR2_X1   g027(.A(KEYINPUT72), .B(G110), .Z(new_n214));
  OAI22_X1  g028(.A1(new_n207), .A2(new_n214), .B1(new_n208), .B2(new_n209), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT73), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT73), .B1(new_n213), .B2(new_n215), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n211), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(KEYINPUT74), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n225), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n211), .B(new_n227), .C1(new_n218), .C2(new_n219), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G217), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT69), .B(G902), .Z(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G234), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(G902), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n226), .A2(new_n231), .A3(new_n228), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT25), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n226), .A2(new_n238), .A3(new_n231), .A4(new_n228), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n232), .B(KEYINPUT71), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n234), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G237), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n221), .A3(G210), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(KEYINPUT27), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G101), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n199), .A2(G143), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT0), .B(G128), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT11), .B1(new_n259), .B2(G134), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(G134), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(KEYINPUT11), .A3(G134), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G137), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(G137), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n267), .A2(new_n263), .A3(new_n258), .A4(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n257), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(KEYINPUT2), .B2(G113), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n274));
  INV_X1    g088(.A(G113), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT64), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT2), .A2(G113), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT65), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(KEYINPUT2), .A3(G113), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n273), .A2(new_n276), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n203), .A2(G116), .ZN(new_n283));
  INV_X1    g097(.A(G116), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G119), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n283), .B2(new_n285), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n283), .A2(new_n285), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n276), .A2(new_n273), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n278), .A2(new_n280), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n252), .A2(new_n295), .A3(G128), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n249), .B(new_n251), .C1(KEYINPUT1), .C2(new_n205), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n266), .A2(G137), .ZN(new_n298));
  OAI21_X1  g112(.A(G131), .B1(new_n298), .B2(new_n261), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n296), .A2(new_n269), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n271), .A2(new_n290), .A3(new_n294), .A4(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n284), .A2(G119), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n203), .A2(G116), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT66), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n294), .B1(new_n306), .B2(new_n281), .ZN(new_n307));
  INV_X1    g121(.A(new_n300), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n267), .A2(new_n263), .A3(new_n268), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G131), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n310), .A2(new_n269), .B1(new_n254), .B2(new_n256), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n307), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n248), .B1(new_n301), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n301), .A2(new_n248), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n247), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n307), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT30), .B1(new_n308), .B2(new_n311), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n271), .A2(new_n320), .A3(new_n300), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n318), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n247), .ZN(new_n323));
  INV_X1    g137(.A(new_n301), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT67), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT31), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n308), .A2(new_n311), .A3(KEYINPUT30), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n320), .B1(new_n271), .B2(new_n300), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n307), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n330), .A2(new_n326), .A3(new_n247), .A4(new_n301), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT31), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n317), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(G472), .A2(G902), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(KEYINPUT32), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT32), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n332), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n319), .A2(new_n321), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n324), .B1(new_n339), .B2(new_n307), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n340), .A2(new_n326), .A3(KEYINPUT31), .A4(new_n247), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n316), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n335), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n337), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n336), .A2(KEYINPUT70), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n338), .A2(new_n341), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n343), .B1(new_n346), .B2(new_n317), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT32), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n231), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT68), .B1(new_n301), .B2(new_n248), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n313), .A2(new_n352), .ZN(new_n353));
  AOI211_X1 g167(.A(KEYINPUT68), .B(new_n248), .C1(new_n301), .C2(new_n312), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n323), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n351), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n323), .B1(new_n322), .B2(new_n324), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n314), .A2(new_n315), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n356), .B(new_n359), .C1(new_n360), .C2(new_n323), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G472), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n242), .B1(new_n350), .B2(new_n363), .ZN(new_n364));
  XOR2_X1   g178(.A(KEYINPUT88), .B(G475), .Z(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n243), .A2(new_n221), .A3(G214), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n250), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n243), .A2(new_n221), .A3(G143), .A4(G214), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(KEYINPUT17), .A3(G131), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n193), .A2(new_n200), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n368), .A2(new_n373), .A3(new_n258), .A4(new_n369), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT86), .B1(new_n370), .B2(G131), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n370), .A2(G131), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n372), .B1(new_n377), .B2(KEYINPUT17), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n197), .A2(KEYINPUT84), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n191), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n381), .A3(G146), .ZN(new_n382));
  INV_X1    g196(.A(new_n212), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT85), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT18), .A2(G131), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n370), .B(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n382), .A2(new_n388), .A3(new_n383), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n378), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G113), .B(G122), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n378), .A2(new_n394), .A3(new_n390), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G902), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n366), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(G475), .A2(G902), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT19), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n379), .B2(new_n381), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n191), .A2(KEYINPUT19), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n199), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n377), .A2(new_n405), .A3(new_n193), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n394), .B1(new_n390), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n397), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI211_X1 g223(.A(KEYINPUT87), .B(new_n394), .C1(new_n390), .C2(new_n406), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n401), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT20), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n413), .B(new_n401), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n400), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G116), .B(G122), .ZN(new_n416));
  INV_X1    g230(.A(G107), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT89), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n416), .B(G107), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n250), .A2(G128), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n205), .A2(G143), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT90), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT90), .B1(new_n423), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n266), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(KEYINPUT13), .ZN(new_n429));
  MUX2_X1   g243(.A(KEYINPUT13), .B(new_n429), .S(new_n423), .Z(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G134), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n419), .A2(new_n422), .A3(new_n428), .A4(new_n431), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n284), .A2(G122), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n417), .B1(new_n433), .B2(KEYINPUT14), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(new_n416), .ZN(new_n435));
  INV_X1    g249(.A(new_n428), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n426), .A2(new_n266), .A3(new_n427), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT9), .B(G234), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n440), .A2(new_n230), .A3(G953), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n432), .A2(new_n438), .A3(new_n441), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n231), .ZN(new_n446));
  INV_X1    g260(.A(G478), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(KEYINPUT15), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n446), .B(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n415), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(G234), .A2(G237), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n452), .A2(G952), .A3(new_n221), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n351), .A2(G953), .A3(new_n452), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(G898), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G469), .ZN(new_n457));
  XOR2_X1   g271(.A(G110), .B(G140), .Z(new_n458));
  INV_X1    g272(.A(G227), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(G953), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n458), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n310), .A2(new_n269), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n462), .A2(KEYINPUT77), .ZN(new_n463));
  INV_X1    g277(.A(G101), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT3), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n465), .A2(new_n417), .A3(KEYINPUT76), .A4(G104), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n417), .A2(KEYINPUT76), .A3(G104), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT3), .B1(new_n393), .B2(G107), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n464), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n417), .A2(G104), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n393), .A2(G107), .ZN(new_n471));
  OAI21_X1  g285(.A(G101), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n296), .A2(new_n297), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n463), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT12), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(KEYINPUT10), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G101), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(KEYINPUT4), .A3(new_n469), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT4), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n483), .A3(G101), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n257), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n462), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT10), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n473), .B2(new_n474), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n479), .A2(new_n485), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT12), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n463), .B(new_n490), .C1(new_n475), .C2(new_n476), .ZN(new_n491));
  AND4_X1   g305(.A1(new_n461), .A2(new_n478), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n479), .A2(new_n485), .A3(new_n488), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n462), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n461), .B1(new_n494), .B2(new_n489), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n457), .B(new_n231), .C1(new_n492), .C2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n478), .A2(new_n489), .A3(new_n491), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n461), .B(KEYINPUT75), .Z(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(new_n461), .A3(new_n489), .ZN(new_n500));
  AOI21_X1  g314(.A(G902), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n496), .B1(new_n501), .B2(new_n457), .ZN(new_n502));
  OAI21_X1  g316(.A(G221), .B1(new_n440), .B2(G902), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n451), .A2(new_n456), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n482), .A2(new_n307), .A3(new_n484), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT5), .B1(new_n287), .B2(new_n288), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT5), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n275), .B1(new_n302), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n469), .A2(new_n472), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n294), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G110), .B(G122), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n506), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n257), .A2(G125), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n296), .A2(new_n195), .A3(new_n297), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G224), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(G953), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT7), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n517), .B1(new_n518), .B2(G953), .ZN(new_n522));
  OAI221_X1 g336(.A(new_n514), .B1(new_n517), .B2(new_n521), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n513), .B(KEYINPUT8), .Z(new_n524));
  NAND2_X1  g338(.A1(new_n291), .A2(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n509), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n511), .A2(new_n294), .A3(new_n526), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n507), .A2(new_n509), .B1(new_n281), .B2(new_n291), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(new_n511), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT81), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT81), .B1(new_n528), .B2(new_n511), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n524), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n399), .B1(new_n523), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n506), .A2(new_n512), .ZN(new_n535));
  INV_X1    g349(.A(new_n513), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(KEYINPUT6), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT80), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n513), .B1(new_n506), .B2(new_n512), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT79), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT6), .B(new_n514), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  AOI211_X1 g356(.A(KEYINPUT79), .B(new_n513), .C1(new_n506), .C2(new_n512), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n537), .A2(KEYINPUT79), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n540), .A2(new_n541), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT80), .A4(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n538), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n515), .A2(new_n519), .A3(new_n516), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n522), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n534), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G210), .B1(G237), .B2(G902), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT82), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT82), .ZN(new_n555));
  INV_X1    g369(.A(new_n553), .ZN(new_n556));
  INV_X1    g370(.A(new_n551), .ZN(new_n557));
  AOI211_X1 g371(.A(new_n557), .B(new_n538), .C1(new_n544), .C2(new_n548), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n555), .B(new_n556), .C1(new_n558), .C2(new_n534), .ZN(new_n559));
  INV_X1    g373(.A(new_n538), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n541), .B1(new_n535), .B2(new_n536), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT80), .B1(new_n563), .B2(new_n547), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n542), .A2(new_n539), .A3(new_n543), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n551), .B(new_n560), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n534), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n553), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n554), .A2(new_n559), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT83), .ZN(new_n570));
  OAI21_X1  g384(.A(G214), .B1(G237), .B2(G902), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT78), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n569), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n570), .B1(new_n569), .B2(new_n573), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n364), .B(new_n505), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G101), .ZN(G3));
  INV_X1    g391(.A(new_n347), .ZN(new_n578));
  OAI21_X1  g392(.A(G472), .B1(new_n342), .B2(new_n351), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n504), .A2(new_n242), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT91), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n584));
  NOR4_X1   g398(.A1(new_n580), .A2(new_n504), .A3(new_n584), .A4(new_n242), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n571), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n556), .B1(new_n558), .B2(new_n534), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n587), .B1(new_n588), .B2(new_n568), .ZN(new_n589));
  INV_X1    g403(.A(new_n400), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n390), .A2(new_n406), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT87), .B1(new_n591), .B2(new_n394), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n407), .A2(new_n408), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n397), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n413), .B1(new_n594), .B2(new_n401), .ZN(new_n595));
  INV_X1    g409(.A(new_n414), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n445), .A2(new_n447), .A3(new_n231), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT92), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n444), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n445), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n443), .B(new_n444), .C1(new_n600), .C2(new_n599), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n351), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n598), .B1(new_n604), .B2(new_n447), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n597), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n456), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n586), .A2(new_n589), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT34), .B(G104), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  OAI211_X1 g425(.A(new_n449), .B(new_n590), .C1(new_n595), .C2(new_n596), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT93), .B1(new_n612), .B2(new_n456), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT93), .ZN(new_n614));
  INV_X1    g428(.A(new_n456), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n415), .A2(new_n614), .A3(new_n615), .A4(new_n449), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n586), .A2(new_n589), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT35), .B(G107), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G9));
  NOR2_X1   g434(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n216), .B(new_n217), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT94), .B1(new_n622), .B2(new_n211), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT94), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n220), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n621), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n622), .A2(KEYINPUT94), .A3(new_n211), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n220), .A2(new_n624), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n627), .B(new_n628), .C1(KEYINPUT36), .C2(new_n225), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n626), .A2(new_n629), .A3(new_n233), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n237), .B2(new_n241), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n580), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n505), .B(new_n633), .C1(new_n574), .C2(new_n575), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT37), .B(G110), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n453), .B1(new_n454), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n612), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n589), .A2(new_n631), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n504), .B1(new_n350), .B2(new_n363), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n205), .ZN(G30));
  INV_X1    g457(.A(new_n504), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n638), .B(KEYINPUT39), .Z(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n646), .A2(KEYINPUT40), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n415), .A2(new_n450), .ZN(new_n648));
  AND4_X1   g462(.A1(new_n571), .A2(new_n647), .A3(new_n632), .A4(new_n648), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n569), .A2(KEYINPUT38), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n569), .A2(KEYINPUT38), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n247), .B1(new_n301), .B2(new_n312), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n399), .B1(new_n325), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G472), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n350), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n646), .A2(KEYINPUT40), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n649), .A2(new_n652), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G143), .ZN(G45));
  NOR4_X1   g473(.A1(new_n342), .A2(KEYINPUT70), .A3(new_n337), .A4(new_n343), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n348), .B1(new_n347), .B2(KEYINPUT32), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n660), .B1(new_n661), .B2(new_n344), .ZN(new_n662));
  INV_X1    g476(.A(new_n363), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n644), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n415), .A2(new_n605), .A3(new_n638), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n588), .A2(new_n568), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n571), .A4(new_n631), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT95), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  AOI211_X1 g482(.A(new_n556), .B(new_n534), .C1(new_n549), .C2(new_n551), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n553), .B1(new_n566), .B2(new_n567), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n571), .B(new_n631), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n638), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n597), .A2(new_n606), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT95), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n641), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  OAI21_X1  g492(.A(new_n571), .B1(new_n669), .B2(new_n670), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n231), .B1(new_n492), .B2(new_n495), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(G469), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n503), .A3(new_n496), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT96), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n681), .A2(KEYINPUT96), .A3(new_n503), .A4(new_n496), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n364), .A2(new_n687), .A3(new_n608), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT97), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT41), .B(G113), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND3_X1  g505(.A1(new_n364), .A2(new_n687), .A3(new_n617), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  NAND2_X1  g507(.A1(new_n350), .A2(new_n363), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n415), .A2(new_n631), .A3(new_n450), .A4(new_n615), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n687), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  NOR2_X1   g512(.A1(new_n686), .A2(new_n456), .ZN(new_n699));
  INV_X1    g513(.A(new_n346), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT98), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n353), .B2(new_n354), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT68), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n313), .A2(new_n703), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n704), .B(KEYINPUT98), .C1(new_n313), .C2(new_n352), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n247), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n335), .B1(new_n700), .B2(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n239), .A2(new_n240), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n708), .A2(new_n236), .B1(new_n233), .B2(new_n229), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n707), .A2(new_n709), .A3(new_n579), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n699), .A2(new_n589), .A3(new_n648), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  INV_X1    g527(.A(KEYINPUT99), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n666), .A2(new_n571), .A3(new_n684), .A4(new_n685), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n707), .A2(new_n631), .A3(new_n579), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n665), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n714), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n707), .A2(new_n631), .A3(new_n579), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n673), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n686), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT99), .A4(new_n589), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  NAND3_X1  g538(.A1(new_n363), .A2(new_n336), .A3(new_n344), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n709), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(KEYINPUT42), .A3(new_n665), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n669), .B1(KEYINPUT82), .B2(new_n588), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n559), .A3(new_n571), .A4(new_n644), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT100), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n726), .A2(new_n732), .A3(new_n673), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT100), .ZN(new_n734));
  AND4_X1   g548(.A1(new_n559), .A2(new_n554), .A3(new_n568), .A4(new_n571), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(new_n734), .A3(new_n644), .A4(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n364), .A2(new_n735), .A3(new_n644), .A4(new_n665), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n731), .A2(new_n736), .B1(new_n737), .B2(new_n732), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n258), .ZN(G33));
  NAND4_X1  g553(.A1(new_n364), .A2(new_n735), .A3(new_n644), .A4(new_n639), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  NAND2_X1  g555(.A1(new_n606), .A2(new_n415), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT101), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n581), .B2(new_n632), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n580), .A2(KEYINPUT101), .A3(new_n631), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n748), .A2(KEYINPUT44), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(KEYINPUT44), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n499), .A2(new_n500), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT45), .ZN(new_n752));
  OAI21_X1  g566(.A(G469), .B1(new_n752), .B2(G902), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n496), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n503), .A3(new_n645), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n749), .A2(new_n735), .A3(new_n750), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  NAND2_X1  g574(.A1(new_n756), .A2(new_n503), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n762));
  OR3_X1    g576(.A1(new_n761), .A2(KEYINPUT102), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(KEYINPUT102), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n762), .A2(KEYINPUT102), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n761), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n735), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n769), .A2(new_n709), .A3(new_n694), .A4(new_n673), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  AND2_X1   g586(.A1(new_n681), .A2(new_n496), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT49), .Z(new_n774));
  NAND3_X1  g588(.A1(new_n709), .A2(new_n573), .A3(new_n503), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n775), .A2(new_n742), .ZN(new_n776));
  OR4_X1    g590(.A1(new_n652), .A2(new_n656), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n650), .A2(new_n587), .A3(new_n651), .A4(new_n721), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n744), .A2(new_n453), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT110), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(KEYINPUT110), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n710), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT113), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(KEYINPUT50), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n735), .A2(new_n721), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT114), .Z(new_n788));
  INV_X1    g602(.A(new_n453), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n656), .A2(new_n242), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n415), .A2(new_n605), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n785), .A2(KEYINPUT50), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n786), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n782), .A2(new_n783), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n788), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n799), .B1(new_n788), .B2(new_n798), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n716), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n773), .B(KEYINPUT111), .Z(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n503), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n735), .B(new_n784), .C1(new_n768), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT109), .B1(new_n797), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT51), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  OAI211_X1 g623(.A(KEYINPUT109), .B(new_n809), .C1(new_n797), .C2(new_n806), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n727), .B1(new_n800), .B2(new_n801), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT48), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT48), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n813), .B(new_n727), .C1(new_n800), .C2(new_n801), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n788), .A2(new_n597), .A3(new_n606), .A4(new_n790), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n784), .A2(new_n687), .ZN(new_n818));
  AND4_X1   g632(.A1(G952), .A2(new_n817), .A3(new_n221), .A4(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n816), .B1(new_n815), .B2(new_n819), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n808), .B(new_n810), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n451), .A2(new_n632), .A3(new_n638), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n641), .A2(new_n735), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n735), .A2(new_n644), .A3(new_n720), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n740), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n731), .A2(new_n736), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n737), .A2(new_n732), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT104), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n612), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n415), .A2(KEYINPUT104), .A3(new_n449), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n456), .B1(new_n833), .B2(new_n607), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n586), .B(new_n834), .C1(new_n574), .C2(new_n575), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n576), .A2(new_n634), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n688), .A2(new_n692), .A3(new_n697), .A4(new_n712), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n829), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n718), .A2(new_n722), .B1(new_n641), .B2(new_n640), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n589), .A2(new_n648), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n504), .A2(new_n631), .A3(new_n638), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n656), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n842), .A2(new_n677), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT105), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n842), .A2(new_n677), .A3(KEYINPUT52), .A4(new_n846), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n847), .A2(KEYINPUT105), .A3(new_n848), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n841), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(KEYINPUT106), .B(KEYINPUT53), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n849), .A2(new_n851), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT103), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n838), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n715), .A2(new_n695), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n686), .A2(new_n710), .A3(new_n456), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n860), .A2(new_n694), .B1(new_n844), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(KEYINPUT103), .A3(new_n688), .A4(new_n692), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n837), .A3(new_n829), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n856), .B1(new_n857), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT108), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n849), .A2(new_n851), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n836), .B1(new_n859), .B2(new_n863), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n829), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT108), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n871), .A3(new_n856), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n855), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OR3_X1    g689(.A1(new_n870), .A2(KEYINPUT107), .A3(new_n856), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT107), .B1(new_n870), .B2(new_n856), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n852), .A2(new_n869), .A3(new_n829), .A4(new_n853), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n876), .A2(new_n877), .B1(new_n839), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n875), .B1(new_n879), .B2(new_n874), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n822), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(G952), .A2(G953), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n777), .B1(new_n881), .B2(new_n882), .ZN(G75));
  AND3_X1   g697(.A1(new_n870), .A2(new_n871), .A3(new_n856), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n871), .B1(new_n870), .B2(new_n856), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n854), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n351), .A3(new_n556), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n549), .A2(new_n551), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n558), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT55), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n221), .A2(G952), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n887), .A2(new_n889), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n887), .A2(KEYINPUT118), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n892), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n896), .B1(new_n897), .B2(new_n899), .ZN(G51));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n873), .A2(new_n231), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n752), .A2(G469), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n901), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n886), .A2(new_n351), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n906), .A2(KEYINPUT119), .A3(new_n903), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(G469), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT57), .Z(new_n910));
  NOR2_X1   g724(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n873), .A2(new_n874), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n492), .A2(new_n495), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n894), .B1(new_n908), .B2(new_n915), .ZN(G54));
  NAND4_X1  g730(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .A4(new_n594), .ZN(new_n917));
  INV_X1    g731(.A(new_n594), .ZN(new_n918));
  NAND2_X1  g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n906), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n917), .A2(new_n895), .A3(new_n920), .ZN(G60));
  NOR2_X1   g735(.A1(new_n911), .A2(new_n912), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n602), .A2(new_n603), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT120), .ZN(new_n924));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT59), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n895), .B1(new_n922), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n924), .B1(new_n880), .B2(new_n926), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT121), .Z(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT60), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n867), .A2(new_n872), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(new_n854), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n626), .A2(new_n629), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n894), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n229), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n873), .B2(new_n934), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n938), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n886), .A2(new_n937), .A3(new_n933), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n940), .A2(new_n895), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n941), .A3(new_n895), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n945), .A2(KEYINPUT61), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n943), .A2(new_n947), .ZN(G66));
  NOR3_X1   g762(.A1(new_n455), .A2(new_n518), .A3(new_n221), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n869), .B2(new_n221), .ZN(new_n950));
  INV_X1    g764(.A(new_n549), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(G898), .B2(new_n221), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n950), .B(new_n952), .ZN(G69));
  AND2_X1   g767(.A1(new_n842), .A2(new_n677), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n658), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT62), .Z(new_n956));
  AOI21_X1  g770(.A(new_n646), .B1(new_n833), .B2(new_n607), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(new_n364), .A3(new_n735), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n759), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n959), .A2(KEYINPUT123), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n959), .A2(KEYINPUT123), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n956), .B(new_n771), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n221), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n403), .A2(new_n404), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n339), .B(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n221), .A2(G900), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n758), .A2(new_n844), .A3(new_n727), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n771), .A2(new_n759), .A3(new_n740), .A4(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n738), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n954), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n968), .B1(new_n975), .B2(new_n221), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n967), .B1(new_n976), .B2(new_n966), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n459), .B2(new_n637), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT124), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n979), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n981), .B(new_n967), .C1(new_n976), .C2(new_n966), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT126), .ZN(new_n986));
  INV_X1    g800(.A(new_n869), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n975), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n323), .A3(new_n340), .ZN(new_n989));
  INV_X1    g803(.A(new_n985), .ZN(new_n990));
  INV_X1    g804(.A(new_n325), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n359), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT127), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n879), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n986), .B1(new_n962), .B2(new_n987), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n340), .A2(new_n323), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n894), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n989), .A2(new_n994), .A3(new_n997), .ZN(G57));
endmodule


