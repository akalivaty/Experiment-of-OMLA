

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U547 ( .A1(n516), .A2(n623), .ZN(n1049) );
  INV_X1 U548 ( .A(n571), .ZN(n1024) );
  AND2_X2 U549 ( .A1(n559), .A2(n520), .ZN(n689) );
  NAND2_X1 U550 ( .A1(n689), .A2(G81), .ZN(n617) );
  INV_X1 U551 ( .A(KEYINPUT40), .ZN(n551) );
  XOR2_X1 U552 ( .A(n753), .B(KEYINPUT28), .Z(n754) );
  NAND2_X1 U553 ( .A1(n526), .A2(KEYINPUT29), .ZN(n525) );
  INV_X1 U554 ( .A(n754), .ZN(n526) );
  NAND2_X1 U555 ( .A1(n540), .A2(G8), .ZN(n539) );
  INV_X1 U556 ( .A(KEYINPUT32), .ZN(n540) );
  NOR2_X1 U557 ( .A1(G1966), .A2(n815), .ZN(n764) );
  NOR2_X1 U558 ( .A1(n834), .A2(n836), .ZN(n736) );
  XNOR2_X1 U559 ( .A(n519), .B(n518), .ZN(n517) );
  INV_X1 U560 ( .A(KEYINPUT13), .ZN(n518) );
  XOR2_X1 U561 ( .A(KEYINPUT107), .B(n865), .Z(n866) );
  NOR2_X1 U562 ( .A1(n552), .A2(n551), .ZN(n550) );
  NAND2_X1 U563 ( .A1(n547), .A2(n546), .ZN(n545) );
  NAND2_X1 U564 ( .A1(n548), .A2(n551), .ZN(n547) );
  NAND2_X1 U565 ( .A1(n866), .A2(n514), .ZN(n546) );
  INV_X1 U566 ( .A(n866), .ZN(n548) );
  AND2_X1 U567 ( .A1(n527), .A2(n524), .ZN(n523) );
  AND2_X1 U568 ( .A1(n525), .A2(n760), .ZN(n524) );
  NAND2_X1 U569 ( .A1(n522), .A2(KEYINPUT29), .ZN(n521) );
  BUF_X1 U570 ( .A(n761), .Z(n780) );
  INV_X1 U571 ( .A(G8), .ZN(n534) );
  NAND2_X1 U572 ( .A1(n537), .A2(n536), .ZN(n535) );
  INV_X1 U573 ( .A(n786), .ZN(n537) );
  INV_X1 U574 ( .A(KEYINPUT99), .ZN(n778) );
  NOR2_X1 U575 ( .A1(n538), .A2(n532), .ZN(n531) );
  NAND2_X1 U576 ( .A1(n535), .A2(n533), .ZN(n532) );
  NOR2_X1 U577 ( .A1(n541), .A2(n539), .ZN(n538) );
  NAND2_X1 U578 ( .A1(n534), .A2(KEYINPUT32), .ZN(n533) );
  XNOR2_X1 U579 ( .A(n728), .B(n727), .ZN(n834) );
  NOR2_X1 U580 ( .A1(n726), .A2(G1384), .ZN(n728) );
  NAND2_X1 U581 ( .A1(n761), .A2(G8), .ZN(n762) );
  XNOR2_X1 U582 ( .A(n570), .B(n569), .ZN(n584) );
  NOR2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n569) );
  XNOR2_X1 U584 ( .A(n568), .B(KEYINPUT17), .ZN(n570) );
  INV_X1 U585 ( .A(KEYINPUT68), .ZN(n568) );
  NOR2_X1 U586 ( .A1(n622), .A2(n517), .ZN(n516) );
  INV_X1 U587 ( .A(G543), .ZN(n520) );
  NAND2_X1 U588 ( .A1(n866), .A2(n551), .ZN(n543) );
  XOR2_X1 U589 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U590 ( .A(n736), .ZN(n761) );
  XNOR2_X2 U591 ( .A(n576), .B(KEYINPUT67), .ZN(n585) );
  AND2_X1 U592 ( .A1(n786), .A2(KEYINPUT32), .ZN(n512) );
  AND2_X1 U593 ( .A1(n847), .A2(n859), .ZN(n513) );
  OR2_X1 U594 ( .A1(n851), .A2(KEYINPUT40), .ZN(n514) );
  NOR2_X1 U595 ( .A1(n815), .A2(n803), .ZN(n515) );
  NAND2_X1 U596 ( .A1(n621), .A2(n620), .ZN(n519) );
  NAND2_X1 U597 ( .A1(n523), .A2(n521), .ZN(n777) );
  INV_X1 U598 ( .A(n529), .ZN(n522) );
  NAND2_X1 U599 ( .A1(n529), .A2(n528), .ZN(n527) );
  AND2_X1 U600 ( .A1(n754), .A2(n755), .ZN(n528) );
  NAND2_X1 U601 ( .A1(n751), .A2(n750), .ZN(n529) );
  NAND2_X1 U602 ( .A1(n531), .A2(n530), .ZN(n794) );
  NAND2_X1 U603 ( .A1(n541), .A2(n512), .ZN(n530) );
  INV_X1 U604 ( .A(n539), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n779), .B(n778), .ZN(n541) );
  OR2_X1 U606 ( .A1(n544), .A2(n542), .ZN(G329) );
  NOR2_X1 U607 ( .A1(n553), .A2(n543), .ZN(n542) );
  NAND2_X1 U608 ( .A1(n549), .A2(n545), .ZN(n544) );
  NAND2_X1 U609 ( .A1(n553), .A2(n550), .ZN(n549) );
  INV_X1 U610 ( .A(n851), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n850), .B(n849), .ZN(n553) );
  OR2_X1 U612 ( .A1(n815), .A2(n814), .ZN(n554) );
  INV_X1 U613 ( .A(KEYINPUT26), .ZN(n729) );
  INV_X1 U614 ( .A(KEYINPUT97), .ZN(n741) );
  BUF_X1 U615 ( .A(n736), .Z(n756) );
  INV_X1 U616 ( .A(G168), .ZN(n769) );
  INV_X1 U617 ( .A(KEYINPUT29), .ZN(n755) );
  INV_X1 U618 ( .A(KEYINPUT31), .ZN(n774) );
  INV_X1 U619 ( .A(KEYINPUT95), .ZN(n763) );
  INV_X1 U620 ( .A(KEYINPUT104), .ZN(n849) );
  NAND2_X1 U621 ( .A1(n694), .A2(G56), .ZN(n616) );
  INV_X1 U622 ( .A(KEYINPUT1), .ZN(n560) );
  NOR2_X1 U623 ( .A1(G651), .A2(n678), .ZN(n695) );
  NAND2_X1 U624 ( .A1(n689), .A2(G89), .ZN(n555) );
  XNOR2_X1 U625 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  XOR2_X1 U626 ( .A(G543), .B(KEYINPUT0), .Z(n678) );
  INV_X1 U627 ( .A(G651), .ZN(n559) );
  NOR2_X2 U628 ( .A1(n678), .A2(n559), .ZN(n690) );
  NAND2_X1 U629 ( .A1(G76), .A2(n690), .ZN(n556) );
  NAND2_X1 U630 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U631 ( .A(n558), .B(KEYINPUT5), .ZN(n566) );
  NOR2_X1 U632 ( .A1(G543), .A2(n559), .ZN(n561) );
  XNOR2_X2 U633 ( .A(n561), .B(n560), .ZN(n694) );
  NAND2_X1 U634 ( .A1(G63), .A2(n694), .ZN(n563) );
  NAND2_X1 U635 ( .A1(G51), .A2(n695), .ZN(n562) );
  NAND2_X1 U636 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U637 ( .A(KEYINPUT6), .B(n564), .Z(n565) );
  NAND2_X1 U638 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U639 ( .A(n567), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 U640 ( .A(n584), .ZN(n571) );
  NAND2_X1 U641 ( .A1(G137), .A2(n1024), .ZN(n575) );
  INV_X1 U642 ( .A(G2104), .ZN(n577) );
  NOR2_X1 U643 ( .A1(n577), .A2(G2105), .ZN(n572) );
  XNOR2_X1 U644 ( .A(n572), .B(KEYINPUT66), .ZN(n604) );
  NAND2_X1 U645 ( .A1(n604), .A2(G101), .ZN(n573) );
  XOR2_X1 U646 ( .A(KEYINPUT23), .B(n573), .Z(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G2105), .A2(G2104), .ZN(n576) );
  NAND2_X1 U649 ( .A1(G113), .A2(n585), .ZN(n579) );
  AND2_X1 U650 ( .A1(n577), .A2(G2105), .ZN(n1019) );
  NAND2_X1 U651 ( .A1(G125), .A2(n1019), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X2 U653 ( .A1(n581), .A2(n580), .ZN(G160) );
  NAND2_X1 U654 ( .A1(n1019), .A2(G126), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G102), .A2(n604), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n584), .A2(G138), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n585), .A2(G114), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n591) );
  INV_X1 U661 ( .A(KEYINPUT87), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n591), .B(n590), .ZN(n726) );
  BUF_X1 U663 ( .A(n726), .Z(G164) );
  XOR2_X1 U664 ( .A(G2427), .B(G2446), .Z(n594) );
  XNOR2_X1 U665 ( .A(G1348), .B(G2430), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n594), .B(n593), .ZN(n595) );
  XOR2_X1 U667 ( .A(n595), .B(G2435), .Z(n597) );
  XNOR2_X1 U668 ( .A(G1341), .B(G2438), .ZN(n596) );
  XNOR2_X1 U669 ( .A(n597), .B(n596), .ZN(n601) );
  XOR2_X1 U670 ( .A(G2454), .B(G2451), .Z(n599) );
  XNOR2_X1 U671 ( .A(KEYINPUT108), .B(G2443), .ZN(n598) );
  XNOR2_X1 U672 ( .A(n599), .B(n598), .ZN(n600) );
  XOR2_X1 U673 ( .A(n601), .B(n600), .Z(n602) );
  AND2_X1 U674 ( .A1(G14), .A2(n602), .ZN(G401) );
  AND2_X1 U675 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U676 ( .A1(G123), .A2(n1019), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT18), .ZN(n611) );
  BUF_X1 U678 ( .A(n604), .Z(n1022) );
  NAND2_X1 U679 ( .A1(G99), .A2(n1022), .ZN(n606) );
  NAND2_X1 U680 ( .A1(G135), .A2(n1024), .ZN(n605) );
  NAND2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U682 ( .A1(G111), .A2(n585), .ZN(n607) );
  XNOR2_X1 U683 ( .A(KEYINPUT79), .B(n607), .ZN(n608) );
  NOR2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U686 ( .A(KEYINPUT80), .B(n612), .ZN(n1041) );
  XNOR2_X1 U687 ( .A(n1041), .B(G2096), .ZN(n613) );
  OR2_X1 U688 ( .A1(G2100), .A2(n613), .ZN(G156) );
  INV_X1 U689 ( .A(G57), .ZN(G237) );
  INV_X1 U690 ( .A(G132), .ZN(G219) );
  NAND2_X1 U691 ( .A1(G7), .A2(G661), .ZN(n614) );
  XOR2_X1 U692 ( .A(n614), .B(KEYINPUT10), .Z(n867) );
  NAND2_X1 U693 ( .A1(n867), .A2(G567), .ZN(n615) );
  XOR2_X1 U694 ( .A(KEYINPUT11), .B(n615), .Z(G234) );
  XOR2_X1 U695 ( .A(KEYINPUT14), .B(n616), .Z(n622) );
  XOR2_X1 U696 ( .A(KEYINPUT12), .B(KEYINPUT75), .Z(n618) );
  XNOR2_X1 U697 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U698 ( .A(KEYINPUT74), .B(n619), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n690), .A2(G68), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n695), .A2(G43), .ZN(n623) );
  INV_X1 U701 ( .A(G860), .ZN(n665) );
  OR2_X1 U702 ( .A1(n1049), .A2(n665), .ZN(G153) );
  NAND2_X1 U703 ( .A1(G64), .A2(n694), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G52), .A2(n695), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G90), .A2(n689), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G77), .A2(n690), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U709 ( .A(KEYINPUT70), .B(n628), .Z(n629) );
  XNOR2_X1 U710 ( .A(KEYINPUT9), .B(n629), .ZN(n630) );
  NOR2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U712 ( .A(KEYINPUT71), .B(n632), .ZN(G301) );
  NAND2_X1 U713 ( .A1(G868), .A2(G301), .ZN(n642) );
  NAND2_X1 U714 ( .A1(G54), .A2(n695), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G92), .A2(n689), .ZN(n634) );
  NAND2_X1 U716 ( .A1(G79), .A2(n690), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n694), .A2(G66), .ZN(n635) );
  XOR2_X1 U719 ( .A(KEYINPUT76), .B(n635), .Z(n636) );
  NOR2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U722 ( .A(n640), .B(KEYINPUT15), .Z(n954) );
  INV_X1 U723 ( .A(G868), .ZN(n709) );
  NAND2_X1 U724 ( .A1(n954), .A2(n709), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(G284) );
  NAND2_X1 U726 ( .A1(G65), .A2(n694), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G53), .A2(n695), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U729 ( .A1(G91), .A2(n689), .ZN(n646) );
  NAND2_X1 U730 ( .A1(G78), .A2(n690), .ZN(n645) );
  NAND2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U732 ( .A1(n648), .A2(n647), .ZN(n955) );
  XOR2_X1 U733 ( .A(n955), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U734 ( .A1(G299), .A2(G868), .ZN(n649) );
  XOR2_X1 U735 ( .A(KEYINPUT77), .B(n649), .Z(n651) );
  NOR2_X1 U736 ( .A1(G286), .A2(n709), .ZN(n650) );
  NOR2_X1 U737 ( .A1(n651), .A2(n650), .ZN(G297) );
  NAND2_X1 U738 ( .A1(G559), .A2(n665), .ZN(n652) );
  XNOR2_X1 U739 ( .A(KEYINPUT78), .B(n652), .ZN(n653) );
  INV_X1 U740 ( .A(n954), .ZN(n1050) );
  NAND2_X1 U741 ( .A1(n653), .A2(n1050), .ZN(n654) );
  XNOR2_X1 U742 ( .A(KEYINPUT16), .B(n654), .ZN(G148) );
  NOR2_X1 U743 ( .A1(G868), .A2(n1049), .ZN(n657) );
  NAND2_X1 U744 ( .A1(G868), .A2(n1050), .ZN(n655) );
  NOR2_X1 U745 ( .A1(G559), .A2(n655), .ZN(n656) );
  NOR2_X1 U746 ( .A1(n657), .A2(n656), .ZN(G282) );
  NAND2_X1 U747 ( .A1(G93), .A2(n689), .ZN(n659) );
  NAND2_X1 U748 ( .A1(G67), .A2(n694), .ZN(n658) );
  NAND2_X1 U749 ( .A1(n659), .A2(n658), .ZN(n663) );
  NAND2_X1 U750 ( .A1(G80), .A2(n690), .ZN(n661) );
  NAND2_X1 U751 ( .A1(G55), .A2(n695), .ZN(n660) );
  NAND2_X1 U752 ( .A1(n661), .A2(n660), .ZN(n662) );
  OR2_X1 U753 ( .A1(n663), .A2(n662), .ZN(n708) );
  NAND2_X1 U754 ( .A1(G559), .A2(n1050), .ZN(n664) );
  XOR2_X1 U755 ( .A(n1049), .B(n664), .Z(n706) );
  NAND2_X1 U756 ( .A1(n665), .A2(n706), .ZN(n666) );
  XNOR2_X1 U757 ( .A(n666), .B(KEYINPUT81), .ZN(n667) );
  XOR2_X1 U758 ( .A(n708), .B(n667), .Z(G145) );
  NAND2_X1 U759 ( .A1(G60), .A2(n694), .ZN(n669) );
  NAND2_X1 U760 ( .A1(G47), .A2(n695), .ZN(n668) );
  NAND2_X1 U761 ( .A1(n669), .A2(n668), .ZN(n672) );
  NAND2_X1 U762 ( .A1(G85), .A2(n689), .ZN(n670) );
  XNOR2_X1 U763 ( .A(KEYINPUT69), .B(n670), .ZN(n671) );
  NOR2_X1 U764 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U765 ( .A1(n690), .A2(G72), .ZN(n673) );
  NAND2_X1 U766 ( .A1(n674), .A2(n673), .ZN(G290) );
  NAND2_X1 U767 ( .A1(G49), .A2(n695), .ZN(n676) );
  NAND2_X1 U768 ( .A1(G74), .A2(G651), .ZN(n675) );
  NAND2_X1 U769 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U770 ( .A1(n694), .A2(n677), .ZN(n680) );
  NAND2_X1 U771 ( .A1(n678), .A2(G87), .ZN(n679) );
  NAND2_X1 U772 ( .A1(n680), .A2(n679), .ZN(G288) );
  NAND2_X1 U773 ( .A1(G73), .A2(n690), .ZN(n681) );
  XNOR2_X1 U774 ( .A(n681), .B(KEYINPUT2), .ZN(n688) );
  NAND2_X1 U775 ( .A1(G61), .A2(n694), .ZN(n683) );
  NAND2_X1 U776 ( .A1(G48), .A2(n695), .ZN(n682) );
  NAND2_X1 U777 ( .A1(n683), .A2(n682), .ZN(n686) );
  NAND2_X1 U778 ( .A1(n689), .A2(G86), .ZN(n684) );
  XOR2_X1 U779 ( .A(KEYINPUT82), .B(n684), .Z(n685) );
  NOR2_X1 U780 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U781 ( .A1(n688), .A2(n687), .ZN(G305) );
  NAND2_X1 U782 ( .A1(n689), .A2(G88), .ZN(n693) );
  NAND2_X1 U783 ( .A1(G75), .A2(n690), .ZN(n691) );
  XOR2_X1 U784 ( .A(KEYINPUT83), .B(n691), .Z(n692) );
  NAND2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n699) );
  NAND2_X1 U786 ( .A1(G62), .A2(n694), .ZN(n697) );
  NAND2_X1 U787 ( .A1(G50), .A2(n695), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U789 ( .A1(n699), .A2(n698), .ZN(G166) );
  XNOR2_X1 U790 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n700) );
  XOR2_X1 U791 ( .A(n700), .B(n708), .Z(n703) );
  XNOR2_X1 U792 ( .A(G299), .B(G290), .ZN(n701) );
  XNOR2_X1 U793 ( .A(n701), .B(G288), .ZN(n702) );
  XNOR2_X1 U794 ( .A(n703), .B(n702), .ZN(n705) );
  XNOR2_X1 U795 ( .A(G305), .B(G166), .ZN(n704) );
  XNOR2_X1 U796 ( .A(n705), .B(n704), .ZN(n1048) );
  XNOR2_X1 U797 ( .A(n706), .B(n1048), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n707), .A2(G868), .ZN(n711) );
  NAND2_X1 U799 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n711), .A2(n710), .ZN(G295) );
  NAND2_X1 U801 ( .A1(G2078), .A2(G2084), .ZN(n712) );
  XOR2_X1 U802 ( .A(KEYINPUT20), .B(n712), .Z(n713) );
  NAND2_X1 U803 ( .A1(G2090), .A2(n713), .ZN(n714) );
  XNOR2_X1 U804 ( .A(KEYINPUT21), .B(n714), .ZN(n715) );
  NAND2_X1 U805 ( .A1(n715), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U806 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  XNOR2_X1 U807 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U808 ( .A1(G219), .A2(G220), .ZN(n717) );
  XNOR2_X1 U809 ( .A(KEYINPUT22), .B(KEYINPUT85), .ZN(n716) );
  XNOR2_X1 U810 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U811 ( .A1(n718), .A2(G218), .ZN(n719) );
  NAND2_X1 U812 ( .A1(G96), .A2(n719), .ZN(n995) );
  NAND2_X1 U813 ( .A1(G2106), .A2(n995), .ZN(n723) );
  NAND2_X1 U814 ( .A1(G120), .A2(G69), .ZN(n720) );
  NOR2_X1 U815 ( .A1(G237), .A2(n720), .ZN(n721) );
  NAND2_X1 U816 ( .A1(G108), .A2(n721), .ZN(n994) );
  NAND2_X1 U817 ( .A1(G567), .A2(n994), .ZN(n722) );
  NAND2_X1 U818 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U819 ( .A(KEYINPUT86), .B(n724), .ZN(n871) );
  NAND2_X1 U820 ( .A1(G661), .A2(G483), .ZN(n725) );
  NOR2_X1 U821 ( .A1(n871), .A2(n725), .ZN(n870) );
  NAND2_X1 U822 ( .A1(n870), .A2(G36), .ZN(G176) );
  XOR2_X1 U823 ( .A(G166), .B(KEYINPUT88), .Z(G303) );
  INV_X1 U824 ( .A(G301), .ZN(G171) );
  INV_X1 U825 ( .A(KEYINPUT64), .ZN(n727) );
  NAND2_X1 U826 ( .A1(G160), .A2(G40), .ZN(n836) );
  NAND2_X1 U827 ( .A1(n736), .A2(G1996), .ZN(n730) );
  XNOR2_X1 U828 ( .A(n730), .B(n729), .ZN(n734) );
  NAND2_X1 U829 ( .A1(n761), .A2(G1341), .ZN(n732) );
  INV_X1 U830 ( .A(n1049), .ZN(n731) );
  NAND2_X1 U831 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U832 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U833 ( .A(n735), .B(KEYINPUT65), .ZN(n743) );
  OR2_X1 U834 ( .A1(n743), .A2(n954), .ZN(n740) );
  NOR2_X1 U835 ( .A1(n756), .A2(G1348), .ZN(n738) );
  NOR2_X1 U836 ( .A1(G2067), .A2(n780), .ZN(n737) );
  NOR2_X1 U837 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U838 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X1 U839 ( .A(n742), .B(n741), .ZN(n745) );
  NAND2_X1 U840 ( .A1(n954), .A2(n743), .ZN(n744) );
  NAND2_X1 U841 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U842 ( .A(n746), .B(KEYINPUT98), .ZN(n751) );
  NAND2_X1 U843 ( .A1(n756), .A2(G2072), .ZN(n747) );
  XNOR2_X1 U844 ( .A(n747), .B(KEYINPUT27), .ZN(n749) );
  INV_X1 U845 ( .A(G1956), .ZN(n1007) );
  NOR2_X1 U846 ( .A1(n1007), .A2(n756), .ZN(n748) );
  NOR2_X1 U847 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U848 ( .A1(n752), .A2(n955), .ZN(n750) );
  NOR2_X1 U849 ( .A1(n752), .A2(n955), .ZN(n753) );
  XOR2_X1 U850 ( .A(G2078), .B(KEYINPUT25), .Z(n887) );
  NAND2_X1 U851 ( .A1(n756), .A2(n887), .ZN(n758) );
  NAND2_X1 U852 ( .A1(G1961), .A2(n780), .ZN(n757) );
  NAND2_X1 U853 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U854 ( .A(KEYINPUT96), .B(n759), .Z(n771) );
  NAND2_X1 U855 ( .A1(n771), .A2(G171), .ZN(n760) );
  XOR2_X2 U856 ( .A(KEYINPUT93), .B(n762), .Z(n815) );
  XNOR2_X1 U857 ( .A(n764), .B(n763), .ZN(n790) );
  NOR2_X1 U858 ( .A1(G2084), .A2(n780), .ZN(n765) );
  XNOR2_X1 U859 ( .A(KEYINPUT94), .B(n765), .ZN(n787) );
  INV_X1 U860 ( .A(n787), .ZN(n766) );
  NAND2_X1 U861 ( .A1(G8), .A2(n766), .ZN(n767) );
  NOR2_X1 U862 ( .A1(n790), .A2(n767), .ZN(n768) );
  XNOR2_X1 U863 ( .A(n768), .B(KEYINPUT30), .ZN(n770) );
  AND2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n773) );
  NOR2_X1 U865 ( .A1(G171), .A2(n771), .ZN(n772) );
  NOR2_X1 U866 ( .A1(n773), .A2(n772), .ZN(n775) );
  XNOR2_X1 U867 ( .A(n775), .B(n774), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n788) );
  NAND2_X1 U869 ( .A1(n788), .A2(G286), .ZN(n779) );
  NOR2_X1 U870 ( .A1(G2090), .A2(n780), .ZN(n781) );
  XOR2_X1 U871 ( .A(KEYINPUT101), .B(n781), .Z(n784) );
  NOR2_X1 U872 ( .A1(G1971), .A2(n815), .ZN(n782) );
  XNOR2_X1 U873 ( .A(n782), .B(KEYINPUT100), .ZN(n783) );
  NOR2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n785), .A2(G303), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n787), .A2(G8), .ZN(n792) );
  INV_X1 U877 ( .A(n788), .ZN(n789) );
  NOR2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n802) );
  NOR2_X1 U881 ( .A1(G303), .A2(G2090), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G8), .A2(n795), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n802), .A2(n796), .ZN(n797) );
  NAND2_X1 U884 ( .A1(n797), .A2(n815), .ZN(n811) );
  NOR2_X1 U885 ( .A1(G1976), .A2(G288), .ZN(n969) );
  NOR2_X1 U886 ( .A1(G303), .A2(G1971), .ZN(n978) );
  NOR2_X1 U887 ( .A1(n969), .A2(n978), .ZN(n798) );
  XNOR2_X1 U888 ( .A(n798), .B(KEYINPUT102), .ZN(n800) );
  INV_X1 U889 ( .A(KEYINPUT33), .ZN(n799) );
  AND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n809) );
  NAND2_X1 U892 ( .A1(G1976), .A2(G288), .ZN(n970) );
  INV_X1 U893 ( .A(n970), .ZN(n803) );
  OR2_X1 U894 ( .A1(KEYINPUT33), .A2(n515), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n969), .A2(KEYINPUT33), .ZN(n804) );
  OR2_X1 U896 ( .A1(n804), .A2(n815), .ZN(n805) );
  AND2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U898 ( .A(G1981), .B(G305), .Z(n962) );
  AND2_X1 U899 ( .A1(n807), .A2(n962), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U901 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U902 ( .A(n812), .B(KEYINPUT103), .ZN(n816) );
  NOR2_X1 U903 ( .A1(G1981), .A2(G305), .ZN(n813) );
  XOR2_X1 U904 ( .A(n813), .B(KEYINPUT24), .Z(n814) );
  NAND2_X1 U905 ( .A1(n816), .A2(n554), .ZN(n848) );
  NAND2_X1 U906 ( .A1(G117), .A2(n585), .ZN(n818) );
  NAND2_X1 U907 ( .A1(G129), .A2(n1019), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U909 ( .A(KEYINPUT90), .B(n819), .ZN(n823) );
  NAND2_X1 U910 ( .A1(n1022), .A2(G105), .ZN(n820) );
  XNOR2_X1 U911 ( .A(n820), .B(KEYINPUT38), .ZN(n821) );
  XNOR2_X1 U912 ( .A(n821), .B(KEYINPUT91), .ZN(n822) );
  NOR2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U914 ( .A1(G141), .A2(n1024), .ZN(n824) );
  NAND2_X1 U915 ( .A1(n825), .A2(n824), .ZN(n1038) );
  AND2_X1 U916 ( .A1(n1038), .A2(G1996), .ZN(n833) );
  NAND2_X1 U917 ( .A1(G95), .A2(n1022), .ZN(n827) );
  NAND2_X1 U918 ( .A1(G131), .A2(n1024), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n831) );
  NAND2_X1 U920 ( .A1(G107), .A2(n585), .ZN(n829) );
  NAND2_X1 U921 ( .A1(G119), .A2(n1019), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n1033) );
  XNOR2_X1 U924 ( .A(G1991), .B(KEYINPUT89), .ZN(n886) );
  NOR2_X1 U925 ( .A1(n1033), .A2(n886), .ZN(n832) );
  NOR2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n909) );
  INV_X1 U927 ( .A(n834), .ZN(n835) );
  NOR2_X1 U928 ( .A1(n836), .A2(n835), .ZN(n864) );
  XOR2_X1 U929 ( .A(n864), .B(KEYINPUT92), .Z(n837) );
  NOR2_X1 U930 ( .A1(n909), .A2(n837), .ZN(n855) );
  INV_X1 U931 ( .A(n855), .ZN(n847) );
  NAND2_X1 U932 ( .A1(G104), .A2(n1022), .ZN(n839) );
  NAND2_X1 U933 ( .A1(G140), .A2(n1024), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U935 ( .A(KEYINPUT34), .B(n840), .ZN(n845) );
  NAND2_X1 U936 ( .A1(G116), .A2(n585), .ZN(n842) );
  NAND2_X1 U937 ( .A1(G128), .A2(n1019), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n842), .A2(n841), .ZN(n843) );
  XOR2_X1 U939 ( .A(KEYINPUT35), .B(n843), .Z(n844) );
  NOR2_X1 U940 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U941 ( .A(KEYINPUT36), .B(n846), .ZN(n1045) );
  XNOR2_X1 U942 ( .A(G2067), .B(KEYINPUT37), .ZN(n861) );
  NOR2_X1 U943 ( .A1(n1045), .A2(n861), .ZN(n911) );
  NAND2_X1 U944 ( .A1(n864), .A2(n911), .ZN(n859) );
  NAND2_X1 U945 ( .A1(n848), .A2(n513), .ZN(n850) );
  XNOR2_X1 U946 ( .A(G1986), .B(G290), .ZN(n959) );
  NAND2_X1 U947 ( .A1(n864), .A2(n959), .ZN(n851) );
  NOR2_X1 U948 ( .A1(G1996), .A2(n1038), .ZN(n903) );
  NOR2_X1 U949 ( .A1(G1986), .A2(G290), .ZN(n852) );
  AND2_X1 U950 ( .A1(n886), .A2(n1033), .ZN(n900) );
  NOR2_X1 U951 ( .A1(n852), .A2(n900), .ZN(n853) );
  XOR2_X1 U952 ( .A(KEYINPUT105), .B(n853), .Z(n854) );
  NOR2_X1 U953 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n856), .B(KEYINPUT106), .ZN(n857) );
  NOR2_X1 U955 ( .A1(n903), .A2(n857), .ZN(n858) );
  XNOR2_X1 U956 ( .A(KEYINPUT39), .B(n858), .ZN(n860) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n862) );
  NAND2_X1 U958 ( .A1(n1045), .A2(n861), .ZN(n913) );
  NAND2_X1 U959 ( .A1(n862), .A2(n913), .ZN(n863) );
  NAND2_X1 U960 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G2106), .A2(n867), .ZN(G217) );
  INV_X1 U962 ( .A(n867), .ZN(G223) );
  AND2_X1 U963 ( .A1(G15), .A2(G2), .ZN(n868) );
  NAND2_X1 U964 ( .A1(G661), .A2(n868), .ZN(G259) );
  NAND2_X1 U965 ( .A1(G3), .A2(G1), .ZN(n869) );
  NAND2_X1 U966 ( .A1(n870), .A2(n869), .ZN(G188) );
  INV_X1 U967 ( .A(n871), .ZN(G319) );
  XNOR2_X1 U968 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  XOR2_X1 U969 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  NAND2_X1 U971 ( .A1(G124), .A2(n1019), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n872), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U973 ( .A1(n1024), .A2(G136), .ZN(n873) );
  XOR2_X1 U974 ( .A(KEYINPUT115), .B(n873), .Z(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U976 ( .A1(n585), .A2(G112), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G100), .A2(n1022), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(G162) );
  XOR2_X1 U980 ( .A(G32), .B(G1996), .Z(n880) );
  NAND2_X1 U981 ( .A1(n880), .A2(G28), .ZN(n885) );
  XNOR2_X1 U982 ( .A(G2067), .B(G26), .ZN(n882) );
  XNOR2_X1 U983 ( .A(G33), .B(G2072), .ZN(n881) );
  NOR2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n883), .B(KEYINPUT123), .ZN(n884) );
  NOR2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n891) );
  XOR2_X1 U987 ( .A(n886), .B(G25), .Z(n889) );
  XNOR2_X1 U988 ( .A(G27), .B(n887), .ZN(n888) );
  NOR2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n892), .B(KEYINPUT53), .ZN(n895) );
  XOR2_X1 U992 ( .A(G2084), .B(G34), .Z(n893) );
  XNOR2_X1 U993 ( .A(KEYINPUT54), .B(n893), .ZN(n894) );
  NAND2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n897) );
  XNOR2_X1 U995 ( .A(G35), .B(G2090), .ZN(n896) );
  NOR2_X1 U996 ( .A1(n897), .A2(n896), .ZN(n988) );
  NAND2_X1 U997 ( .A1(KEYINPUT55), .A2(n988), .ZN(n898) );
  NAND2_X1 U998 ( .A1(G11), .A2(n898), .ZN(n987) );
  XOR2_X1 U999 ( .A(G2084), .B(G160), .Z(n899) );
  NOR2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(n1041), .A2(n901), .ZN(n907) );
  XOR2_X1 U1002 ( .A(G2090), .B(G162), .Z(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(KEYINPUT51), .B(n904), .Z(n905) );
  XNOR2_X1 U1005 ( .A(n905), .B(KEYINPUT121), .ZN(n906) );
  NOR2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n912), .B(KEYINPUT122), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(n927) );
  NAND2_X1 U1011 ( .A1(G103), .A2(n1022), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(G139), .A2(n1024), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n922) );
  NAND2_X1 U1014 ( .A1(n1019), .A2(G127), .ZN(n917) );
  XOR2_X1 U1015 ( .A(KEYINPUT119), .B(n917), .Z(n919) );
  NAND2_X1 U1016 ( .A1(n585), .A2(G115), .ZN(n918) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1018 ( .A(KEYINPUT47), .B(n920), .Z(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n1032) );
  XOR2_X1 U1020 ( .A(G2072), .B(n1032), .Z(n924) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1023 ( .A(KEYINPUT50), .B(n925), .Z(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(KEYINPUT52), .B(n928), .ZN(n930) );
  INV_X1 U1026 ( .A(KEYINPUT55), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1028 ( .A1(n931), .A2(G29), .ZN(n985) );
  XOR2_X1 U1029 ( .A(G20), .B(G1956), .Z(n935) );
  XNOR2_X1 U1030 ( .A(G1981), .B(G6), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(G1341), .B(G19), .ZN(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1034 ( .A(KEYINPUT59), .B(G1348), .Z(n936) );
  XNOR2_X1 U1035 ( .A(G4), .B(n936), .ZN(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(KEYINPUT60), .B(n939), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(G1966), .B(G21), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(G5), .B(G1961), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G1971), .B(G22), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(G23), .B(G1976), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n947) );
  XOR2_X1 U1045 ( .A(G1986), .B(G24), .Z(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(KEYINPUT58), .B(n948), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1049 ( .A(KEYINPUT61), .B(n951), .Z(n953) );
  XOR2_X1 U1050 ( .A(G16), .B(KEYINPUT125), .Z(n952) );
  NOR2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n982) );
  XOR2_X1 U1052 ( .A(G16), .B(KEYINPUT56), .Z(n980) );
  XOR2_X1 U1053 ( .A(n954), .B(G1348), .Z(n961) );
  XOR2_X1 U1054 ( .A(n1007), .B(n955), .Z(n957) );
  NAND2_X1 U1055 ( .A1(G1971), .A2(G303), .ZN(n956) );
  NAND2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n968) );
  XOR2_X1 U1059 ( .A(G301), .B(G1961), .Z(n966) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G168), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1062 ( .A(n964), .B(KEYINPUT57), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(G1341), .B(n1049), .ZN(n974) );
  INV_X1 U1066 ( .A(n969), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(KEYINPUT124), .B(n972), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(n983), .B(KEYINPUT126), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n992) );
  INV_X1 U1077 ( .A(n988), .ZN(n990) );
  NOR2_X1 U1078 ( .A1(G29), .A2(KEYINPUT55), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1081 ( .A(KEYINPUT62), .B(n993), .Z(G311) );
  XNOR2_X1 U1082 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1083 ( .A(G120), .ZN(G236) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1085 ( .A(n996), .B(KEYINPUT111), .Z(G325) );
  INV_X1 U1086 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1087 ( .A(KEYINPUT112), .B(G2678), .Z(n998) );
  XNOR2_X1 U1088 ( .A(G2090), .B(G2072), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(n998), .B(n997), .ZN(n1002) );
  XOR2_X1 U1090 ( .A(KEYINPUT43), .B(KEYINPUT42), .Z(n1000) );
  XNOR2_X1 U1091 ( .A(G2067), .B(KEYINPUT113), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(n1000), .B(n999), .ZN(n1001) );
  XOR2_X1 U1093 ( .A(n1002), .B(n1001), .Z(n1004) );
  XNOR2_X1 U1094 ( .A(G2096), .B(G2100), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(n1004), .B(n1003), .ZN(n1006) );
  XOR2_X1 U1096 ( .A(G2078), .B(G2084), .Z(n1005) );
  XNOR2_X1 U1097 ( .A(n1006), .B(n1005), .ZN(G227) );
  XOR2_X1 U1098 ( .A(G1986), .B(n1007), .Z(n1018) );
  XOR2_X1 U1099 ( .A(G1976), .B(G1971), .Z(n1009) );
  XNOR2_X1 U1100 ( .A(G1981), .B(G1961), .ZN(n1008) );
  XNOR2_X1 U1101 ( .A(n1009), .B(n1008), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(G2474), .B(KEYINPUT114), .Z(n1012) );
  INV_X1 U1103 ( .A(G1996), .ZN(n1010) );
  XOR2_X1 U1104 ( .A(n1010), .B(G1966), .Z(n1011) );
  XNOR2_X1 U1105 ( .A(n1012), .B(n1011), .ZN(n1013) );
  XOR2_X1 U1106 ( .A(n1014), .B(n1013), .Z(n1016) );
  XNOR2_X1 U1107 ( .A(G1991), .B(KEYINPUT41), .ZN(n1015) );
  XNOR2_X1 U1108 ( .A(n1016), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1109 ( .A(n1018), .B(n1017), .ZN(G229) );
  NAND2_X1 U1110 ( .A1(G118), .A2(n585), .ZN(n1021) );
  NAND2_X1 U1111 ( .A1(G130), .A2(n1019), .ZN(n1020) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(G106), .A2(n1022), .ZN(n1023) );
  XNOR2_X1 U1114 ( .A(n1023), .B(KEYINPUT116), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(G142), .A2(n1024), .ZN(n1025) );
  NAND2_X1 U1116 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1117 ( .A(KEYINPUT117), .B(n1027), .ZN(n1028) );
  XNOR2_X1 U1118 ( .A(KEYINPUT45), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1119 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1120 ( .A(n1032), .B(n1031), .Z(n1037) );
  XOR2_X1 U1121 ( .A(KEYINPUT118), .B(KEYINPUT46), .Z(n1035) );
  XNOR2_X1 U1122 ( .A(n1033), .B(KEYINPUT48), .ZN(n1034) );
  XNOR2_X1 U1123 ( .A(n1035), .B(n1034), .ZN(n1036) );
  XOR2_X1 U1124 ( .A(n1037), .B(n1036), .Z(n1040) );
  XOR2_X1 U1125 ( .A(G164), .B(n1038), .Z(n1039) );
  XNOR2_X1 U1126 ( .A(n1040), .B(n1039), .ZN(n1042) );
  XOR2_X1 U1127 ( .A(n1042), .B(n1041), .Z(n1044) );
  XNOR2_X1 U1128 ( .A(G160), .B(G162), .ZN(n1043) );
  XNOR2_X1 U1129 ( .A(n1044), .B(n1043), .ZN(n1046) );
  XOR2_X1 U1130 ( .A(n1046), .B(n1045), .Z(n1047) );
  NOR2_X1 U1131 ( .A1(G37), .A2(n1047), .ZN(G395) );
  XNOR2_X1 U1132 ( .A(n1049), .B(n1048), .ZN(n1052) );
  XOR2_X1 U1133 ( .A(G301), .B(n1050), .Z(n1051) );
  XNOR2_X1 U1134 ( .A(n1052), .B(n1051), .ZN(n1053) );
  XNOR2_X1 U1135 ( .A(n1053), .B(G286), .ZN(n1054) );
  NOR2_X1 U1136 ( .A1(G37), .A2(n1054), .ZN(G397) );
  NOR2_X1 U1137 ( .A1(G227), .A2(G229), .ZN(n1055) );
  XOR2_X1 U1138 ( .A(KEYINPUT49), .B(n1055), .Z(n1056) );
  NAND2_X1 U1139 ( .A1(G319), .A2(n1056), .ZN(n1057) );
  NOR2_X1 U1140 ( .A1(G401), .A2(n1057), .ZN(n1060) );
  NOR2_X1 U1141 ( .A1(G395), .A2(G397), .ZN(n1058) );
  XNOR2_X1 U1142 ( .A(n1058), .B(KEYINPUT120), .ZN(n1059) );
  NAND2_X1 U1143 ( .A1(n1060), .A2(n1059), .ZN(G225) );
  INV_X1 U1144 ( .A(G225), .ZN(G308) );
  INV_X1 U1145 ( .A(G108), .ZN(G238) );
endmodule

