//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n220), .A2(KEYINPUT66), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(KEYINPUT66), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n212), .B1(new_n215), .B2(new_n218), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G226), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n237), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT71), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(new_n213), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n252), .B1(new_n208), .B2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G1), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT72), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT72), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n206), .A2(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(G68), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n253), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G68), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G77), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n207), .A2(G33), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n272), .A2(KEYINPUT11), .ZN(new_n273));
  INV_X1    g0073(.A(new_n256), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n267), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n275), .A2(KEYINPUT12), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(KEYINPUT12), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n276), .A2(new_n277), .B1(new_n272), .B2(KEYINPUT11), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n264), .A2(new_n273), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT76), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT76), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n264), .A2(new_n281), .A3(new_n278), .A4(new_n273), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G232), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(G226), .B2(G1698), .ZN(new_n291));
  INV_X1    g0091(.A(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT3), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT3), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n291), .A2(new_n296), .B1(new_n292), .B2(new_n202), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n288), .B1(new_n297), .B2(new_n285), .ZN(new_n298));
  INV_X1    g0098(.A(new_n287), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n285), .A2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n300), .A2(KEYINPUT75), .ZN(new_n301));
  OAI21_X1  g0101(.A(G238), .B1(new_n300), .B2(KEYINPUT75), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT13), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT14), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(G169), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n304), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n305), .B1(new_n304), .B2(G169), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n284), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(G200), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n283), .B(new_n311), .C1(new_n312), .C2(new_n304), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT8), .B(G58), .ZN(new_n316));
  INV_X1    g0116(.A(G150), .ZN(new_n317));
  INV_X1    g0117(.A(new_n266), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n316), .A2(new_n270), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(G50), .A2(G58), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n207), .B1(new_n320), .B2(new_n267), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n265), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n263), .A2(G50), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n257), .A2(new_n324), .B1(G50), .B2(new_n256), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT3), .B(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G222), .A2(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(G1698), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G223), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(new_n285), .C1(G77), .C2(new_n328), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G41), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n286), .B1(new_n252), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n299), .ZN(new_n336));
  INV_X1    g0136(.A(G226), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n252), .A2(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n287), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n333), .B(new_n336), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n326), .B1(new_n327), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(G179), .B2(new_n340), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(G200), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT74), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n344), .B(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(KEYINPUT9), .B2(new_n326), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n326), .A2(KEYINPUT9), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n312), .B2(new_n340), .ZN(new_n349));
  OR3_X1    g0149(.A1(new_n347), .A2(KEYINPUT10), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT10), .B1(new_n347), .B2(new_n349), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n343), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n300), .A2(G232), .B1(new_n335), .B2(new_n299), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT77), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n293), .A2(new_n295), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n292), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(G223), .A2(G1698), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n337), .B2(G1698), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n357), .A2(new_n359), .B1(G33), .B2(G87), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n353), .B(new_n312), .C1(new_n360), .C2(new_n338), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n336), .B1(new_n339), .B2(new_n289), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n292), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n328), .B2(new_n354), .ZN(new_n364));
  INV_X1    g0164(.A(new_n359), .ZN(new_n365));
  INV_X1    g0165(.A(G87), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n364), .A2(new_n365), .B1(new_n292), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n362), .B1(new_n367), .B2(new_n285), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n361), .B1(new_n368), .B2(G200), .ZN(new_n369));
  INV_X1    g0169(.A(G58), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(new_n267), .ZN(new_n371));
  NOR2_X1   g0171(.A1(G58), .A2(G68), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n266), .A2(G159), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n364), .B2(new_n207), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n355), .A2(new_n377), .A3(new_n207), .A4(new_n356), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G68), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT16), .B(new_n376), .C1(new_n378), .C2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n377), .B1(new_n328), .B2(G20), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n296), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n267), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n382), .B1(new_n385), .B2(new_n375), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n386), .A3(new_n265), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n316), .B1(new_n206), .B2(G20), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n258), .A2(new_n388), .B1(new_n274), .B2(new_n316), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n369), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT79), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT79), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n369), .A2(new_n387), .A3(new_n392), .A4(new_n389), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(KEYINPUT17), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT17), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n369), .A2(new_n387), .A3(new_n395), .A4(new_n389), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n396), .A2(KEYINPUT80), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n387), .A2(new_n389), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n353), .B(G179), .C1(new_n360), .C2(new_n338), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n368), .B2(new_n327), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(KEYINPUT18), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT78), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT78), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n399), .A2(new_n404), .A3(KEYINPUT18), .A4(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n399), .A2(new_n401), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT18), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT80), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n391), .A2(new_n410), .A3(KEYINPUT17), .A4(new_n393), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n398), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n262), .A2(G77), .A3(new_n263), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G20), .A2(G77), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT15), .B(G87), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n415), .B1(new_n316), .B2(new_n318), .C1(new_n270), .C2(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n265), .B1(new_n269), .B2(new_n274), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n328), .A2(G238), .A3(G1698), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n328), .A2(G232), .A3(new_n330), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(new_n203), .C2(new_n328), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n285), .ZN(new_n423));
  INV_X1    g0223(.A(G244), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n423), .B(new_n336), .C1(new_n424), .C2(new_n339), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n419), .B1(G200), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n312), .B2(new_n425), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT73), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n425), .B2(new_n327), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n425), .A2(G179), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n430), .A2(KEYINPUT73), .B1(new_n414), .B2(new_n418), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n315), .A2(new_n352), .A3(new_n413), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT86), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT19), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(new_n207), .A3(G33), .ZN(new_n440));
  OR2_X1    g0240(.A1(KEYINPUT81), .A2(G97), .ZN(new_n441));
  NAND2_X1  g0241(.A1(KEYINPUT81), .A2(G97), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(G87), .A2(G107), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n207), .B1(new_n292), .B2(new_n202), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n443), .B1(new_n447), .B2(KEYINPUT19), .ZN(new_n448));
  AOI211_X1 g0248(.A(G20), .B(new_n267), .C1(new_n355), .C2(new_n356), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n438), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n357), .A2(new_n207), .A3(G68), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n439), .B1(new_n445), .B2(new_n446), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n451), .B(KEYINPUT86), .C1(new_n452), .C2(new_n443), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n453), .A3(new_n265), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n274), .A2(new_n416), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT87), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(KEYINPUT87), .A3(new_n455), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n206), .A2(G33), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n258), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(new_n366), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n463), .B(KEYINPUT89), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT90), .ZN(new_n465));
  INV_X1    g0265(.A(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G1), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n467), .A2(G250), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n286), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n338), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(G238), .A2(G1698), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n424), .B2(G1698), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G116), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n364), .A2(new_n474), .B1(new_n292), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n471), .B1(new_n476), .B2(new_n285), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n465), .B1(new_n477), .B2(G190), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n357), .A2(new_n473), .B1(G33), .B2(G116), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n470), .B1(new_n479), .B2(new_n338), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G200), .ZN(new_n481));
  OAI211_X1 g0281(.A(G190), .B(new_n470), .C1(new_n479), .C2(new_n338), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n478), .B1(new_n483), .B2(new_n465), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n460), .A2(new_n464), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n462), .A2(new_n416), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n454), .A2(KEYINPUT87), .A3(new_n455), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT87), .B1(new_n454), .B2(new_n455), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT88), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT88), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n492), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n477), .A2(new_n307), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n480), .A2(new_n327), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n486), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n441), .A2(new_n442), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(KEYINPUT6), .A3(new_n203), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT82), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G97), .A2(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n204), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n502), .B1(new_n204), .B2(new_n503), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n508), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n328), .A2(new_n377), .A3(G20), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT7), .B1(new_n296), .B2(new_n207), .ZN(new_n511));
  OAI21_X1  g0311(.A(G107), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT83), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT83), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n514), .B(G107), .C1(new_n510), .C2(new_n511), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n509), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n265), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n256), .A2(G97), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n462), .B2(new_n202), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(G41), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n206), .B(G45), .C1(new_n523), .C2(KEYINPUT5), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT85), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n524), .A2(new_n525), .B1(KEYINPUT5), .B2(new_n523), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n525), .B2(new_n524), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n527), .A2(new_n338), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G257), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G283), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n328), .A2(KEYINPUT4), .A3(G244), .A4(new_n330), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n330), .A2(G244), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n355), .B2(new_n356), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n530), .B(new_n531), .C1(new_n533), .C2(KEYINPUT4), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n293), .A2(new_n295), .A3(G250), .A4(G1698), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n535), .B(KEYINPUT84), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n285), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n526), .B(new_n335), .C1(new_n525), .C2(new_n524), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n529), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n327), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n529), .A2(new_n537), .A3(new_n307), .A4(new_n538), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n522), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(G200), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n520), .B1(new_n516), .B2(new_n265), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n529), .A2(new_n537), .A3(G190), .A4(new_n538), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT91), .B1(new_n499), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n497), .B1(new_n491), .B2(new_n493), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT91), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n542), .A2(new_n546), .ZN(new_n551));
  NOR4_X1   g0351(.A1(new_n549), .A2(new_n486), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  OR2_X1    g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT23), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n554), .A2(KEYINPUT93), .B1(new_n555), .B2(new_n203), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n203), .A3(G20), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT93), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n557), .A2(new_n558), .B1(new_n559), .B2(G20), .ZN(new_n560));
  OR3_X1    g0360(.A1(new_n556), .A2(new_n560), .A3(KEYINPUT94), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT94), .B1(new_n556), .B2(new_n560), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(KEYINPUT22), .A2(G87), .ZN(new_n564));
  AOI211_X1 g0364(.A(G20), .B(new_n564), .C1(new_n355), .C2(new_n356), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT92), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n366), .A2(G20), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT22), .B1(new_n328), .B2(new_n567), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n357), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n570));
  INV_X1    g0370(.A(new_n568), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT92), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n563), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT24), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n566), .B1(new_n565), .B2(new_n568), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n570), .A2(KEYINPUT92), .A3(new_n571), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(new_n563), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n253), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n274), .A2(new_n203), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT95), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT25), .ZN(new_n583));
  XOR2_X1   g0383(.A(KEYINPUT95), .B(KEYINPUT25), .Z(new_n584));
  OAI221_X1 g0384(.A(new_n583), .B1(new_n581), .B2(new_n584), .C1(new_n462), .C2(new_n203), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G257), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G1698), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(G250), .B2(G1698), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n364), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(G294), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n292), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n285), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n527), .A2(G264), .A3(new_n338), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n538), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n327), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G179), .B2(new_n595), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n586), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n330), .A2(G264), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n600), .B(new_n364), .C1(new_n587), .C2(new_n330), .ZN(new_n601));
  INV_X1    g0401(.A(G303), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n328), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n285), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n528), .A2(G270), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n604), .A2(new_n538), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n327), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n259), .A2(G116), .A3(new_n261), .A4(new_n461), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n255), .A2(G20), .A3(new_n475), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n253), .B1(G20), .B2(new_n475), .ZN(new_n610));
  INV_X1    g0410(.A(new_n500), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n207), .B(new_n530), .C1(new_n611), .C2(G33), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n612), .A3(KEYINPUT20), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT20), .B1(new_n610), .B2(new_n612), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n608), .B(new_n609), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT21), .B1(new_n607), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n606), .A2(G179), .A3(new_n616), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n604), .A2(new_n538), .A3(new_n605), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n619), .A2(KEYINPUT21), .A3(G169), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n577), .A2(new_n578), .A3(new_n563), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n578), .B1(new_n577), .B2(new_n563), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n265), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n585), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n595), .A2(G200), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n593), .A2(G190), .A3(new_n594), .A4(new_n538), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n625), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n616), .B1(new_n619), .B2(G200), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n312), .B2(new_n619), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n599), .A2(new_n622), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n437), .A2(new_n553), .A3(new_n634), .ZN(G372));
  INV_X1    g0435(.A(KEYINPUT97), .ZN(new_n636));
  INV_X1    g0436(.A(new_n483), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n464), .B(new_n637), .C1(new_n488), .C2(new_n489), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n496), .A2(KEYINPUT96), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n495), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n496), .A2(KEYINPUT96), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n639), .B1(new_n494), .B2(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n580), .A2(new_n585), .A3(new_n629), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(new_n551), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n636), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n643), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n491), .B2(new_n493), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n631), .A2(new_n542), .A3(new_n546), .ZN(new_n650));
  NOR4_X1   g0450(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT97), .A4(new_n639), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n598), .A2(new_n617), .A3(new_n621), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n647), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n492), .B1(new_n460), .B2(new_n487), .ZN(new_n654));
  INV_X1    g0454(.A(new_n493), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n643), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  INV_X1    g0457(.A(new_n542), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .A4(new_n638), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n549), .A2(new_n486), .A3(new_n542), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n659), .B(new_n656), .C1(new_n660), .C2(new_n657), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n437), .B1(new_n653), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n310), .A2(new_n433), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n663), .A2(new_n398), .A3(new_n411), .A4(new_n313), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n408), .A2(new_n402), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n350), .A2(new_n351), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n343), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n662), .A2(new_n668), .ZN(G369));
  NAND2_X1  g0469(.A1(new_n255), .A2(new_n207), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(G213), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n616), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n622), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n633), .ZN(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n675), .B1(new_n580), .B2(new_n585), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n645), .B1(KEYINPUT98), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n681), .A2(KEYINPUT98), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n598), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n599), .A2(new_n675), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n599), .ZN(new_n689));
  INV_X1    g0489(.A(new_n675), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n617), .B2(new_n621), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n685), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n687), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n210), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G1), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n445), .A2(G116), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n698), .A2(new_n699), .B1(new_n216), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT99), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n690), .B1(new_n653), .B2(new_n661), .ZN(new_n703));
  XNOR2_X1  g0503(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n656), .A2(KEYINPUT26), .A3(new_n658), .A4(new_n638), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n660), .B2(KEYINPUT26), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n649), .A2(new_n650), .A3(new_n639), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n599), .A2(new_n622), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n649), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n675), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT101), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT29), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n711), .B2(KEYINPUT29), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n705), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n634), .B(new_n690), .C1(new_n548), .C2(new_n552), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n619), .A2(new_n307), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n529), .A2(new_n537), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n595), .A2(new_n480), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  AND4_X1   g0521(.A1(new_n307), .A2(new_n619), .A3(new_n480), .A4(new_n595), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n720), .A2(new_n721), .B1(new_n722), .B2(new_n539), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n718), .A4(new_n719), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n690), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n716), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n715), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n702), .B1(new_n730), .B2(G1), .ZN(G364));
  NOR2_X1   g0531(.A1(new_n254), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n206), .B1(new_n732), .B2(G45), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n697), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n680), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(G330), .B1(new_n677), .B2(new_n633), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n678), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n695), .A2(new_n296), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G355), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G116), .B2(new_n210), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n247), .A2(G45), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n364), .A2(new_n210), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n466), .B2(new_n217), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n213), .B1(G20), .B2(new_n327), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n741), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n735), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G200), .ZN(new_n754));
  NOR4_X1   g0554(.A1(new_n207), .A2(new_n312), .A3(new_n754), .A4(G179), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR4_X1   g0556(.A1(new_n207), .A2(new_n754), .A3(G179), .A4(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n756), .A2(new_n602), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n207), .A2(new_n307), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G311), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n762), .A2(new_n312), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n296), .B1(new_n764), .B2(new_n765), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G179), .A2(G200), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT103), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n207), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n760), .B(new_n769), .C1(G329), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT102), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n762), .B2(new_n754), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n761), .A2(KEYINPUT102), .A3(G200), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n777), .A2(G190), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n207), .B1(new_n771), .B2(G190), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G326), .A2(new_n780), .B1(new_n782), .B2(G294), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n777), .A2(new_n312), .A3(new_n778), .ZN(new_n784));
  XOR2_X1   g0584(.A(KEYINPUT33), .B(G317), .Z(new_n785));
  OAI211_X1 g0585(.A(new_n775), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n756), .A2(new_n366), .B1(new_n758), .B2(new_n203), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n328), .B1(new_n764), .B2(new_n269), .C1(new_n370), .C2(new_n768), .ZN(new_n788));
  INV_X1    g0588(.A(new_n784), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n787), .B(new_n788), .C1(new_n789), .C2(G68), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n781), .A2(KEYINPUT104), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n781), .A2(KEYINPUT104), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G97), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n774), .A2(G159), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT32), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n796), .A2(KEYINPUT32), .B1(new_n780), .B2(G50), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n790), .A2(new_n795), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n786), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n753), .B1(new_n800), .B2(new_n750), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n736), .A2(new_n738), .B1(new_n742), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n419), .A2(new_n675), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n433), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n804), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n434), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n703), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n434), .A2(new_n675), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n653), .B2(new_n661), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n735), .B1(new_n813), .B2(new_n729), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n729), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n750), .A2(new_n739), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n735), .B1(G77), .B2(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n756), .A2(new_n203), .B1(new_n758), .B2(new_n366), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n296), .B1(new_n764), .B2(new_n475), .C1(new_n591), .C2(new_n768), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n819), .B(new_n820), .C1(G311), .C2(new_n774), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G283), .A2(new_n789), .B1(new_n780), .B2(G303), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n821), .A2(new_n795), .A3(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G143), .A2(new_n767), .B1(new_n763), .B2(G159), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n784), .B2(new_n317), .C1(new_n825), .C2(new_n779), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT34), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n357), .B1(new_n773), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT105), .ZN(new_n832));
  INV_X1    g0632(.A(G50), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n756), .A2(new_n833), .B1(new_n758), .B2(new_n267), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n782), .B2(G58), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n829), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n823), .B1(new_n828), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n818), .B1(new_n837), .B2(new_n750), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n808), .B2(new_n740), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n815), .A2(new_n839), .ZN(G384));
  AND2_X1   g0640(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n842));
  NOR4_X1   g0642(.A1(new_n841), .A2(new_n842), .A3(new_n475), .A4(new_n215), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT36), .ZN(new_n844));
  OR3_X1    g0644(.A1(new_n371), .A2(new_n216), .A3(new_n269), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n833), .A2(G68), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n206), .B(G13), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n376), .B1(new_n378), .B2(new_n380), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n382), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n850), .A2(new_n265), .A3(new_n381), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n673), .B1(new_n851), .B2(new_n389), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n412), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n673), .B1(new_n387), .B2(new_n389), .ZN(new_n854));
  AOI211_X1 g0654(.A(KEYINPUT37), .B(new_n854), .C1(new_n399), .C2(new_n401), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(new_n391), .A3(new_n393), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n391), .A2(new_n393), .ZN(new_n857));
  INV_X1    g0657(.A(new_n401), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n858), .A2(new_n673), .B1(new_n851), .B2(new_n389), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT37), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n853), .A2(KEYINPUT38), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n284), .A2(new_n675), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n310), .A2(new_n313), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(new_n310), .B2(new_n313), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n811), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n659), .A2(new_n656), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n657), .B1(new_n499), .B2(new_n658), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n656), .A2(new_n646), .A3(new_n638), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT97), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n644), .A2(new_n636), .A3(new_n646), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n709), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n872), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n433), .A2(new_n675), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n866), .B(new_n871), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n408), .A2(new_n402), .A3(new_n673), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT106), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n310), .A2(new_n675), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n865), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n853), .B2(new_n861), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT39), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n398), .A2(new_n665), .A3(new_n411), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n854), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n406), .A2(new_n390), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n894), .B2(new_n854), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n856), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n863), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n899), .A3(new_n865), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT107), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n891), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(new_n891), .B2(new_n900), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n888), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n882), .A2(KEYINPUT106), .A3(new_n883), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n886), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n705), .B(new_n437), .C1(new_n713), .C2(new_n714), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n668), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n906), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n808), .B1(new_n868), .B2(new_n869), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n728), .A2(new_n866), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n910), .B1(new_n716), .B2(new_n727), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n913), .B1(new_n898), .B2(new_n865), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n912), .A2(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n916), .A2(new_n437), .A3(new_n728), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n437), .B2(new_n728), .ZN(new_n918));
  OR3_X1    g0718(.A1(new_n917), .A2(new_n918), .A3(new_n679), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n909), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n206), .B2(new_n732), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n909), .A2(new_n919), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n848), .B1(new_n921), .B2(new_n922), .ZN(G367));
  AND3_X1   g0723(.A1(new_n237), .A2(new_n210), .A3(new_n364), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n751), .B1(new_n210), .B2(new_n416), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n735), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n756), .A2(new_n370), .B1(new_n758), .B2(new_n269), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n328), .B1(new_n764), .B2(new_n833), .C1(new_n317), .C2(new_n768), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n927), .B(new_n928), .C1(G137), .C2(new_n774), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n794), .A2(G68), .ZN(new_n930));
  AOI22_X1  g0730(.A1(G143), .A2(new_n780), .B1(new_n789), .B2(G159), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n758), .A2(new_n611), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n364), .B1(new_n764), .B2(new_n759), .C1(new_n602), .C2(new_n768), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n933), .B(new_n934), .C1(G317), .C2(new_n774), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT46), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n756), .B2(new_n475), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n755), .A2(KEYINPUT46), .A3(G116), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n937), .B(new_n938), .C1(new_n784), .C2(new_n591), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT110), .ZN(new_n940));
  AOI22_X1  g0740(.A1(G311), .A2(new_n780), .B1(new_n782), .B2(G107), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n935), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n939), .A2(KEYINPUT110), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n932), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT111), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT47), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n926), .B1(new_n946), .B2(new_n750), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n690), .B1(new_n460), .B2(new_n464), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n649), .A2(new_n639), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n649), .B2(new_n948), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n741), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n733), .B(KEYINPUT109), .Z(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n686), .B(new_n692), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(new_n680), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n729), .A3(new_n715), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n522), .A2(new_n675), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n547), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT108), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n658), .A2(new_n675), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n547), .A2(KEYINPUT108), .A3(new_n958), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n685), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(new_n684), .C2(new_n691), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT45), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT44), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n693), .B2(new_n964), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n965), .B1(new_n684), .B2(new_n691), .ZN(new_n971));
  INV_X1    g0771(.A(new_n964), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(KEYINPUT44), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n968), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n687), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n968), .A2(new_n974), .A3(new_n687), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n730), .B1(new_n957), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n696), .B(KEYINPUT41), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n954), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n689), .A2(new_n965), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n691), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n964), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n961), .A2(new_n963), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n542), .B1(new_n986), .B2(new_n599), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n985), .A2(KEYINPUT42), .B1(new_n690), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT42), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n984), .A2(new_n989), .A3(new_n964), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT43), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n950), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n950), .A2(new_n992), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n988), .A2(new_n992), .A3(new_n950), .A4(new_n990), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n687), .A2(new_n972), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n995), .A2(new_n998), .A3(new_n996), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n952), .B1(new_n982), .B2(new_n1002), .ZN(G387));
  OAI21_X1  g0803(.A(new_n364), .B1(new_n758), .B2(new_n475), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G303), .A2(new_n763), .B1(new_n767), .B2(G317), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n784), .B2(new_n765), .C1(new_n766), .C2(new_n779), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT48), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n782), .A2(G283), .B1(G294), .B2(new_n755), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT49), .Z(new_n1012));
  AOI211_X1 g0812(.A(new_n1004), .B(new_n1012), .C1(G326), .C2(new_n774), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n793), .A2(new_n416), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n774), .A2(G150), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G50), .A2(new_n767), .B1(new_n763), .B2(G68), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n755), .A2(G77), .B1(new_n757), .B2(G97), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n357), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(G159), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1019), .A2(new_n779), .B1(new_n784), .B2(new_n316), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1014), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n750), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n743), .A2(new_n699), .B1(new_n203), .B2(new_n695), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n242), .A2(G45), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT112), .Z(new_n1025));
  AOI211_X1 g0825(.A(G45), .B(new_n699), .C1(G68), .C2(G77), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n316), .A2(G50), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n747), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT113), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1023), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n734), .B1(new_n1031), .B2(new_n751), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1022), .A2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT114), .Z(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n983), .B2(new_n741), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n956), .B2(new_n954), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n957), .A2(new_n696), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n730), .B2(new_n956), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1038), .ZN(G393));
  INV_X1    g0839(.A(new_n979), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n972), .A2(new_n741), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n751), .B1(new_n210), .B2(new_n611), .C1(new_n250), .C2(new_n747), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n735), .A2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n780), .A2(G317), .B1(G311), .B2(new_n767), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT52), .Z(new_n1045));
  AOI21_X1  g0845(.A(new_n328), .B1(new_n763), .B2(G294), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n203), .B2(new_n758), .C1(new_n759), .C2(new_n756), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G322), .B2(new_n774), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G303), .A2(new_n789), .B1(new_n782), .B2(G116), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1045), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n779), .A2(new_n317), .B1(new_n768), .B2(new_n1019), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT51), .Z(new_n1052));
  NAND2_X1  g0852(.A1(new_n794), .A2(G77), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n784), .A2(new_n833), .B1(new_n764), .B2(new_n316), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT115), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n357), .B1(new_n758), .B2(new_n366), .C1(new_n756), .C2(new_n267), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G143), .B2(new_n774), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1050), .B1(new_n1052), .B2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT116), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1043), .B1(new_n1060), .B2(new_n750), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1040), .A2(new_n954), .B1(new_n1041), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n957), .A2(new_n979), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n696), .B1(new_n957), .B2(new_n979), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT117), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT117), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1062), .B(new_n1068), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(G390));
  AND3_X1   g0870(.A1(new_n898), .A2(new_n899), .A3(new_n865), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n899), .B1(new_n864), .B2(new_n865), .ZN(new_n1072));
  OAI21_X1  g0872(.A(KEYINPUT107), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n891), .A2(new_n900), .A3(new_n901), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(new_n740), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n734), .B1(new_n316), .B2(new_n816), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(KEYINPUT54), .B(G143), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n296), .B1(new_n763), .B2(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n833), .B2(new_n758), .C1(new_n830), .C2(new_n768), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n780), .A2(G128), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n755), .A2(G150), .ZN(new_n1083));
  XOR2_X1   g0883(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1084));
  XNOR2_X1  g0884(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1082), .B(new_n1085), .C1(new_n825), .C2(new_n784), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1081), .B(new_n1086), .C1(G125), .C2(new_n774), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n794), .A2(G159), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n296), .B1(new_n764), .B2(new_n611), .C1(new_n475), .C2(new_n768), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n203), .A2(new_n784), .B1(new_n779), .B2(new_n759), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n773), .A2(new_n591), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n756), .A2(new_n366), .B1(new_n758), .B2(new_n267), .ZN(new_n1092));
  NOR4_X1   g0892(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1087), .A2(new_n1088), .B1(new_n1053), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n750), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1077), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1076), .A2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n675), .B(new_n809), .C1(new_n707), .C2(new_n710), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n871), .B1(new_n1098), .B2(new_n881), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n888), .B1(new_n898), .B2(new_n865), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n881), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n812), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n888), .B1(new_n1103), .B2(new_n871), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1101), .B1(new_n1104), .B2(new_n1075), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n679), .B1(new_n716), .B2(new_n727), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1106), .A2(new_n808), .A3(new_n871), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n880), .A2(new_n881), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n887), .B1(new_n1109), .B2(new_n870), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n902), .A2(new_n903), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n679), .B(new_n809), .C1(new_n716), .C2(new_n727), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1099), .A2(new_n1100), .B1(new_n871), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n953), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  AOI211_X1 g0915(.A(KEYINPUT119), .B(new_n1097), .C1(new_n1108), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT119), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1106), .A2(new_n808), .A3(new_n871), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n1101), .C1(new_n1104), .C2(new_n1075), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1110), .A2(new_n1111), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1119), .B(new_n954), .C1(new_n1120), .C2(new_n1118), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1097), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1117), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1116), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1119), .B1(new_n1120), .B2(new_n1118), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1106), .A2(new_n437), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n907), .A2(new_n668), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n871), .B1(new_n1106), .B2(new_n808), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1103), .B1(new_n1107), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n870), .B1(new_n729), .B2(new_n809), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1098), .A2(new_n881), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1118), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1127), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1125), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1108), .A2(new_n1127), .A3(new_n1133), .A4(new_n1119), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n1136), .A3(new_n696), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT120), .B1(new_n1124), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1119), .A2(new_n954), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1118), .B1(new_n1112), .B2(new_n1101), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1122), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT119), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1121), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1143));
  AND4_X1   g0943(.A1(KEYINPUT120), .A2(new_n1137), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1138), .A2(new_n1144), .ZN(G378));
  NAND2_X1  g0945(.A1(new_n914), .A2(new_n915), .ZN(new_n1146));
  AOI221_X4 g0946(.A(new_n910), .B1(new_n864), .B2(new_n865), .C1(new_n716), .C2(new_n727), .ZN(new_n1147));
  OAI211_X1 g0947(.A(G330), .B(new_n1146), .C1(new_n1147), .C2(KEYINPUT40), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n326), .A2(new_n673), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT55), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n352), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n352), .A2(new_n1153), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1150), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1156), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n1149), .A3(new_n1154), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1148), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n916), .A2(G330), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1164), .A2(new_n906), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n905), .A2(new_n904), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1166), .A2(new_n886), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n954), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n735), .B1(G50), .B2(new_n817), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n357), .A2(G41), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G50), .B(new_n1170), .C1(new_n292), .C2(new_n523), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n773), .B2(new_n759), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n767), .A2(G107), .B1(G77), .B2(new_n755), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n370), .B2(new_n758), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(G116), .C2(new_n780), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n784), .A2(new_n202), .B1(new_n764), .B2(new_n416), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT121), .Z(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1177), .A3(new_n930), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT58), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1171), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n784), .A2(new_n830), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G128), .A2(new_n767), .B1(new_n763), .B2(G137), .ZN(new_n1182));
  INV_X1    g0982(.A(G125), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1182), .B1(new_n756), .B2(new_n1078), .C1(new_n779), .C2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1181), .B(new_n1184), .C1(G150), .C2(new_n794), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n292), .B(new_n523), .C1(new_n758), .C2(new_n1019), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G124), .B2(new_n774), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT59), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1180), .B1(new_n1179), .B2(new_n1178), .C1(new_n1187), .C2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1169), .B1(new_n1192), .B2(new_n750), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1162), .B2(new_n740), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1168), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT57), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1166), .A2(new_n886), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT40), .B1(new_n914), .B2(new_n866), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n728), .A2(new_n915), .A3(new_n911), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1198), .A2(new_n1199), .A3(new_n1160), .A4(new_n679), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1162), .B1(new_n916), .B2(G330), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n905), .A2(new_n904), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT106), .B1(new_n882), .B2(new_n883), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n1200), .A2(new_n1201), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1196), .B1(new_n1197), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1127), .B1(new_n1125), .B2(new_n1134), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n697), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1197), .A2(new_n1204), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n907), .A2(new_n668), .A3(new_n1126), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1105), .A2(new_n1107), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1210), .B2(new_n1133), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1196), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1195), .B1(new_n1207), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(G375));
  NAND2_X1  g1014(.A1(new_n870), .A2(new_n739), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n735), .B1(G68), .B2(new_n817), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n794), .A2(G50), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n774), .A2(G128), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n768), .A2(new_n825), .B1(new_n764), .B2(new_n317), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n756), .A2(new_n1019), .B1(new_n758), .B2(new_n370), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1219), .A2(new_n364), .A3(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G132), .A2(new_n780), .B1(new_n789), .B2(new_n1079), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1217), .A2(new_n1218), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n756), .A2(new_n202), .B1(new_n758), .B2(new_n269), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n296), .B1(new_n764), .B2(new_n203), .C1(new_n759), .C2(new_n768), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(G303), .C2(new_n774), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n475), .B2(new_n784), .C1(new_n591), .C2(new_n779), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1223), .B1(new_n1227), .B2(new_n1014), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1216), .B1(new_n1228), .B2(new_n750), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1133), .A2(new_n954), .B1(new_n1215), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1209), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1134), .A2(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n981), .B(KEYINPUT123), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1230), .B1(new_n1232), .B2(new_n1233), .ZN(G381));
  NAND3_X1  g1034(.A1(new_n1036), .A2(new_n802), .A3(new_n1038), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1235), .A2(G381), .A3(G384), .ZN(new_n1236));
  INV_X1    g1036(.A(G387), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G390), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1137), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1213), .A4(new_n1240), .ZN(G407));
  NAND2_X1  g1041(.A1(new_n674), .A2(G213), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1213), .A2(new_n1240), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(G407), .A2(G213), .A3(new_n1244), .ZN(G409));
  AOI21_X1  g1045(.A(new_n802), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1235), .ZN(new_n1248));
  AND3_X1   g1048(.A1(G387), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G387), .B1(new_n1069), .B2(new_n1067), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G390), .A2(new_n1237), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1235), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(new_n1246), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(G387), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1252), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1251), .A2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1213), .B1(new_n1138), .B2(new_n1144), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1208), .A2(new_n1211), .A3(new_n1233), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1240), .B1(new_n1259), .B2(new_n1195), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1243), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1232), .A2(KEYINPUT60), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n697), .B1(new_n1231), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G384), .B1(new_n1265), .B2(new_n1230), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1231), .A2(new_n1263), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n696), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1263), .B1(new_n1134), .B2(new_n1231), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G384), .B(new_n1230), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1266), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1261), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT62), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1242), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1243), .A2(G2897), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1230), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1279));
  INV_X1    g1079(.A(G384), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT124), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n1270), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1281), .B2(new_n1270), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1278), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT124), .B1(new_n1266), .B2(new_n1271), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1277), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1276), .A2(new_n1285), .A3(new_n1287), .ZN(new_n1288));
  XOR2_X1   g1088(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1289));
  NAND3_X1  g1089(.A1(new_n1274), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1273), .A2(KEYINPUT62), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1257), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT126), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1281), .A2(new_n1282), .A3(new_n1270), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1277), .B1(new_n1286), .B2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1284), .A2(new_n1278), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1285), .A2(KEYINPUT125), .A3(new_n1287), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1276), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1281), .A2(KEYINPUT63), .A3(new_n1270), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1275), .A2(new_n1242), .A3(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT61), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1251), .A2(new_n1303), .A3(new_n1256), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT63), .B1(new_n1261), .B2(new_n1272), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  AND4_X1   g1107(.A1(new_n1293), .A2(new_n1300), .A3(new_n1305), .A4(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1309), .A2(new_n1306), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1293), .B1(new_n1310), .B2(new_n1300), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1292), .B1(new_n1308), .B2(new_n1311), .ZN(G405));
  INV_X1    g1112(.A(new_n1240), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1258), .B1(new_n1213), .B2(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1314), .B(new_n1272), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1315), .B(new_n1257), .ZN(G402));
endmodule


