//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n800,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917;
  XOR2_X1   g000(.A(G71gat), .B(G78gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204));
  INV_X1    g003(.A(G71gat), .ZN(new_n205));
  INV_X1    g004(.A(G78gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G57gat), .B(G64gat), .Z(new_n208));
  NAND3_X1  g007(.A1(new_n203), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n207), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(new_n202), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT94), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n215));
  AOI21_X1  g014(.A(G1gat), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G8gat), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n214), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(KEYINPUT88), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n216), .A2(new_n217), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n216), .A2(new_n217), .ZN(new_n223));
  AOI211_X1 g022(.A(G1gat), .B(G8gat), .C1(new_n214), .C2(new_n215), .ZN(new_n224));
  OAI22_X1  g023(.A1(new_n223), .A2(new_n224), .B1(KEYINPUT88), .B2(new_n219), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n213), .A2(KEYINPUT21), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(G231gat), .A2(G233gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G127gat), .B(G155gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(G211gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n229), .A2(new_n231), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n212), .A2(KEYINPUT21), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n236), .B(new_n237), .Z(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n235), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G232gat), .A2(G233gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT41), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G85gat), .A2(G92gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT95), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT7), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G99gat), .A2(G106gat), .ZN(new_n248));
  INV_X1    g047(.A(G85gat), .ZN(new_n249));
  INV_X1    g048(.A(G92gat), .ZN(new_n250));
  AOI22_X1  g049(.A1(KEYINPUT8), .A2(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n244), .A2(KEYINPUT95), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n244), .A2(KEYINPUT95), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n247), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G99gat), .B(G106gat), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n247), .A2(new_n256), .A3(new_n251), .A4(new_n254), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G43gat), .B(G50gat), .Z(new_n261));
  INV_X1    g060(.A(KEYINPUT87), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(G29gat), .A2(G36gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT14), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT14), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(G29gat), .B2(G36gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(G29gat), .A2(G36gat), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n263), .A2(new_n269), .A3(KEYINPUT15), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(new_n262), .B2(new_n261), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT15), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n271), .B2(new_n261), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n243), .B1(new_n260), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT96), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n275), .A2(KEYINPUT17), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT17), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n270), .B(new_n280), .C1(new_n272), .C2(new_n274), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n279), .A2(new_n258), .A3(new_n259), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(new_n242), .A3(new_n241), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n241), .A2(new_n242), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n278), .A2(new_n285), .A3(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n287), .A2(KEYINPUT97), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(KEYINPUT97), .ZN(new_n289));
  XOR2_X1   g088(.A(G134gat), .B(G162gat), .Z(new_n290));
  XNOR2_X1  g089(.A(G190gat), .B(G218gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OR3_X1    g092(.A1(new_n288), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n288), .B2(new_n289), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n240), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n222), .A2(new_n225), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(new_n281), .A3(new_n279), .ZN(new_n299));
  NAND2_X1  g098(.A1(G229gat), .A2(G233gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n276), .A2(new_n222), .A3(new_n225), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n299), .A2(KEYINPUT18), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n300), .B(KEYINPUT13), .Z(new_n303));
  NOR2_X1   g102(.A1(new_n298), .A2(new_n275), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n272), .A2(new_n274), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n222), .A2(new_n225), .B1(new_n305), .B2(new_n270), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT91), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n302), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n308), .B1(new_n302), .B2(new_n307), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT89), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT18), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT89), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n299), .A2(new_n315), .A3(new_n300), .A4(new_n301), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT90), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT90), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n313), .A2(new_n319), .A3(new_n314), .A4(new_n316), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n311), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G113gat), .B(G141gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G169gat), .B(G197gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n321), .A2(KEYINPUT92), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT92), .B1(new_n321), .B2(new_n329), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n302), .A2(new_n307), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT93), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n330), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G230gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n209), .A2(new_n211), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n258), .A2(new_n338), .A3(new_n259), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT98), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n258), .A2(KEYINPUT98), .A3(new_n338), .A4(new_n259), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT100), .B(KEYINPUT10), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n257), .A2(KEYINPUT99), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n255), .B(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n212), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n213), .A2(KEYINPUT10), .A3(new_n260), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n337), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n336), .B1(new_n343), .B2(new_n347), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G120gat), .B(G148gat), .ZN(new_n353));
  INV_X1    g152(.A(G176gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G204gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n352), .B(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n335), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n361));
  INV_X1    g160(.A(G120gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G113gat), .ZN(new_n363));
  INV_X1    g162(.A(G113gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G120gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G113gat), .B(G120gat), .ZN(new_n370));
  INV_X1    g169(.A(G134gat), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n371), .A2(G127gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(G127gat), .ZN(new_n373));
  OAI22_X1  g172(.A1(new_n370), .A2(KEYINPUT1), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G141gat), .B(G148gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT2), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(G155gat), .B2(G162gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n377), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G141gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G148gat), .ZN(new_n383));
  INV_X1    g182(.A(G148gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G141gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G155gat), .B(G162gat), .ZN(new_n387));
  INV_X1    g186(.A(G155gat), .ZN(new_n388));
  INV_X1    g187(.A(G162gat), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT2), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  AND4_X1   g190(.A1(new_n369), .A2(new_n374), .A3(new_n381), .A4(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n361), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n369), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT67), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n381), .A2(new_n391), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n374), .A2(new_n369), .A3(KEYINPUT67), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n397), .A2(new_n393), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n374), .A2(new_n381), .A3(new_n369), .A4(new_n391), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n394), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n381), .A2(new_n391), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT3), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n381), .A2(new_n391), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n395), .A3(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n403), .A2(new_n404), .A3(new_n405), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n405), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT75), .B1(new_n401), .B2(KEYINPUT4), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n374), .A2(new_n369), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n414), .A2(new_n398), .A3(new_n415), .A4(new_n393), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n397), .A2(new_n399), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT4), .B1(new_n418), .B2(new_n406), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n412), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n395), .A2(new_n406), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n405), .B1(new_n421), .B2(new_n401), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT76), .B1(new_n422), .B2(new_n404), .ZN(new_n423));
  INV_X1    g222(.A(new_n405), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n369), .A2(new_n374), .B1(new_n381), .B2(new_n391), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n392), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT76), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(KEYINPUT5), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n411), .B1(new_n420), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT0), .B(G57gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(G85gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(G1gat), .B(G29gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n432), .B(new_n433), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n411), .B(new_n434), .C1(new_n420), .C2(new_n429), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT80), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n430), .A2(KEYINPUT6), .A3(new_n435), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n436), .A2(KEYINPUT80), .A3(new_n437), .A4(new_n438), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT81), .ZN(new_n446));
  NAND2_X1  g245(.A1(G183gat), .A2(G190gat), .ZN(new_n447));
  NOR2_X1   g246(.A1(G169gat), .A2(G176gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT26), .ZN(new_n450));
  NAND2_X1  g249(.A1(G169gat), .A2(G176gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT26), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT27), .B(G183gat), .ZN(new_n455));
  INV_X1    g254(.A(G190gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(KEYINPUT28), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT28), .B1(new_n455), .B2(new_n456), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n447), .B(new_n454), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT24), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n447), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(G183gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n456), .ZN(new_n464));
  NAND3_X1  g263(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT23), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT25), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n469), .B1(new_n448), .B2(KEYINPUT23), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT66), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT66), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n466), .A2(new_n468), .A3(new_n473), .A4(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n477));
  AOI21_X1  g276(.A(G176gat), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n478), .A2(KEYINPUT23), .B1(new_n449), .B2(new_n467), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT64), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n465), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n480), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n464), .B(new_n462), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT25), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n460), .B1(new_n475), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT29), .ZN(new_n486));
  NAND2_X1  g285(.A1(G226gat), .A2(G233gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(G211gat), .B(G218gat), .Z(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G197gat), .B(G204gat), .Z(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT71), .B(G211gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G218gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT22), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n495), .A2(new_n496), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n490), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n495), .A2(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n495), .A2(new_n496), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n489), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n487), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n504), .B(new_n460), .C1(new_n475), .C2(new_n484), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT73), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n503), .B1(new_n488), .B2(new_n505), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI211_X1 g308(.A(KEYINPUT73), .B(new_n503), .C1(new_n488), .C2(new_n505), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(G8gat), .B(G36gat), .Z(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G64gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(G92gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n488), .A2(new_n503), .A3(new_n505), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT37), .B1(new_n516), .B2(new_n508), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT38), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n514), .B(KEYINPUT74), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT37), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n509), .B2(new_n510), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n445), .A2(new_n446), .A3(new_n515), .A4(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n511), .A2(new_n521), .ZN(new_n525));
  INV_X1    g324(.A(new_n514), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT38), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n442), .B1(new_n439), .B2(new_n440), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n529), .A2(new_n515), .A3(new_n523), .A4(new_n444), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT81), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n524), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n503), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n486), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n398), .B1(new_n534), .B2(new_n408), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n486), .B2(new_n409), .ZN(new_n536));
  NAND2_X1  g335(.A1(G228gat), .A2(G233gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n537), .B(G22gat), .Z(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OR3_X1    g338(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G78gat), .B(G106gat), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT31), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(G50gat), .Z(new_n543));
  OR2_X1    g342(.A1(new_n543), .A2(KEYINPUT78), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n539), .B1(new_n535), .B2(new_n536), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(KEYINPUT78), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n547), .B(KEYINPUT79), .Z(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n540), .A2(new_n544), .A3(new_n545), .A4(new_n548), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n515), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n511), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n519), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n511), .A2(KEYINPUT30), .A3(new_n514), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n403), .A2(new_n410), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n424), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(KEYINPUT39), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(new_n435), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n421), .A2(new_n405), .A3(new_n401), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(KEYINPUT39), .A3(new_n563), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n562), .A2(KEYINPUT40), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT40), .B1(new_n562), .B2(new_n564), .ZN(new_n566));
  INV_X1    g365(.A(new_n436), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n552), .B1(new_n558), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n532), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT82), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n485), .B(new_n418), .ZN(new_n573));
  NAND2_X1  g372(.A1(G227gat), .A2(G233gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT68), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(KEYINPUT68), .A3(new_n575), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT33), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n573), .A2(new_n575), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT34), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(KEYINPUT70), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G71gat), .B(G99gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT69), .ZN(new_n588));
  XOR2_X1   g387(.A(G15gat), .B(G43gat), .Z(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  NAND3_X1  g389(.A1(new_n582), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT33), .B1(new_n578), .B2(new_n579), .ZN(new_n592));
  INV_X1    g391(.A(new_n590), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n585), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT32), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n584), .A2(KEYINPUT70), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n580), .B(KEYINPUT32), .C1(KEYINPUT70), .C2(new_n584), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n591), .A2(new_n598), .A3(new_n594), .A4(new_n599), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n443), .A2(new_n439), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n552), .B1(new_n558), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT36), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n532), .A2(KEYINPUT82), .A3(new_n569), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n572), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT84), .ZN(new_n612));
  INV_X1    g411(.A(new_n558), .ZN(new_n613));
  INV_X1    g412(.A(new_n552), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n603), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT83), .B(KEYINPUT35), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n445), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n606), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n603), .A2(new_n614), .A3(new_n613), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT35), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n611), .A2(new_n612), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n612), .B1(new_n611), .B2(new_n622), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n297), .B(new_n360), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(new_n619), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g426(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n625), .A2(new_n613), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(new_n215), .B2(new_n217), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT42), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(G8gat), .B1(new_n625), .B2(new_n613), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n631), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(G1325gat));
  INV_X1    g434(.A(new_n603), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n625), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(G15gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n605), .A2(new_n608), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n638), .B1(G15gat), .B2(new_n641), .ZN(G1326gat));
  NOR2_X1   g441(.A1(new_n625), .A2(new_n614), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT43), .B(G22gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  INV_X1    g446(.A(new_n296), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n611), .B2(new_n622), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n532), .A2(KEYINPUT82), .A3(new_n569), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT82), .B1(new_n532), .B2(new_n569), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n615), .A2(new_n617), .B1(new_n620), .B2(KEYINPUT35), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT84), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n611), .A2(new_n612), .A3(new_n622), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n648), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n651), .B1(new_n659), .B2(new_n650), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n240), .A2(new_n360), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(KEYINPUT103), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G29gat), .B1(new_n666), .B2(new_n619), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n659), .A2(new_n661), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n668), .A2(G29gat), .A3(new_n619), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT45), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(G1328gat));
  OAI21_X1  g470(.A(G36gat), .B1(new_n666), .B2(new_n613), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n668), .A2(G36gat), .A3(new_n613), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT46), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(G1329gat));
  OAI21_X1  g474(.A(G43gat), .B1(new_n662), .B2(new_n640), .ZN(new_n676));
  INV_X1    g475(.A(G43gat), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n659), .A2(new_n677), .A3(new_n603), .A4(new_n661), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(KEYINPUT47), .A3(new_n678), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n679), .A2(KEYINPUT104), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(KEYINPUT104), .ZN(new_n681));
  INV_X1    g480(.A(new_n678), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n639), .B1(new_n663), .B2(new_n665), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(new_n683), .B2(G43gat), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n680), .B(new_n681), .C1(new_n684), .C2(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g484(.A(KEYINPUT48), .B(G50gat), .C1(new_n662), .C2(new_n614), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n668), .A2(G50gat), .A3(new_n614), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n686), .B(new_n687), .C1(KEYINPUT105), .C2(KEYINPUT48), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(KEYINPUT105), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n552), .B1(new_n663), .B2(new_n665), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(G50gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n688), .B1(new_n691), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g491(.A(new_n335), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n240), .A2(new_n296), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n359), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT106), .Z(new_n696));
  NAND2_X1  g495(.A1(new_n611), .A2(new_n622), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n606), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g500(.A(new_n613), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT107), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n704), .B(new_n705), .Z(G1333gat));
  XNOR2_X1  g505(.A(new_n603), .B(KEYINPUT108), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n699), .A2(new_n205), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G71gat), .B1(new_n698), .B2(new_n640), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g510(.A1(new_n698), .A2(new_n614), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(new_n206), .ZN(G1335gat));
  XNOR2_X1  g512(.A(new_n235), .B(new_n238), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n693), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n649), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT51), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n649), .A2(new_n715), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n717), .A2(KEYINPUT109), .A3(new_n720), .ZN(new_n721));
  OR3_X1    g520(.A1(new_n718), .A2(KEYINPUT109), .A3(new_n719), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n359), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n249), .B1(new_n723), .B2(new_n619), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n660), .A2(new_n359), .A3(new_n715), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(G85gat), .A3(new_n606), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n724), .A2(new_n726), .ZN(G1336gat));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n558), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT52), .B1(new_n728), .B2(G92gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n613), .A2(G92gat), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n723), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733));
  INV_X1    g532(.A(new_n359), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n717), .B2(new_n720), .ZN(new_n735));
  AOI22_X1  g534(.A1(new_n728), .A2(G92gat), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n732), .B1(new_n733), .B2(new_n736), .ZN(G1337gat));
  XOR2_X1   g536(.A(KEYINPUT110), .B(G99gat), .Z(new_n738));
  INV_X1    g537(.A(new_n725), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(new_n640), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n636), .A2(new_n738), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n723), .B2(new_n741), .ZN(G1338gat));
  NAND4_X1  g541(.A1(new_n660), .A2(new_n552), .A3(new_n359), .A4(new_n715), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(G106gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n614), .A2(G106gat), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n735), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT53), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n715), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n296), .B1(new_n623), .B2(new_n624), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT44), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n748), .B1(new_n750), .B2(new_n651), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n751), .A2(new_n752), .A3(new_n552), .A4(new_n359), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n743), .A2(KEYINPUT111), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n754), .A3(G106gat), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n721), .A2(new_n359), .A3(new_n722), .A4(new_n745), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n755), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n756), .B1(new_n755), .B2(new_n759), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n747), .B1(new_n760), .B2(new_n761), .ZN(G1339gat));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n348), .A2(new_n763), .A3(new_n337), .A4(new_n349), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(KEYINPUT54), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n348), .A2(new_n337), .A3(new_n349), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n350), .B2(KEYINPUT113), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g569(.A(new_n337), .B(new_n770), .C1(new_n348), .C2(new_n349), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n768), .A2(new_n357), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n768), .A2(KEYINPUT55), .A3(new_n357), .A4(new_n772), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n352), .A2(new_n358), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n693), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n334), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n304), .A2(new_n306), .A3(new_n303), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n326), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n782), .A2(new_n359), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n296), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n782), .A2(new_n785), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n777), .A2(new_n296), .A3(new_n788), .A4(new_n780), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n240), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n694), .A2(new_n734), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n793), .A2(new_n606), .A3(new_n615), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n693), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n359), .ZN(new_n797));
  XOR2_X1   g596(.A(KEYINPUT116), .B(G120gat), .Z(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1341gat));
  NAND2_X1  g598(.A1(new_n794), .A2(new_n714), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G127gat), .ZN(G1342gat));
  NAND3_X1  g600(.A1(new_n794), .A2(new_n371), .A3(new_n296), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT56), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n371), .B1(new_n794), .B2(new_n296), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n803), .A2(new_n804), .ZN(G1343gat));
  AOI211_X1 g604(.A(new_n358), .B(new_n771), .C1(new_n765), .C2(new_n767), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n779), .B(new_n778), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n786), .B1(new_n335), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT118), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n811), .B(new_n786), .C1(new_n335), .C2(new_n808), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n648), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n789), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n240), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n614), .B1(new_n815), .B2(new_n792), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n793), .A2(new_n552), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818));
  MUX2_X1   g617(.A(new_n816), .B(new_n817), .S(new_n818), .Z(new_n819));
  NOR2_X1   g618(.A1(new_n639), .A2(new_n619), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n558), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n382), .B1(new_n824), .B2(new_n693), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n614), .B1(new_n791), .B2(new_n792), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n820), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n335), .A2(G141gat), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n827), .A2(new_n558), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT58), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT119), .B1(new_n826), .B2(new_n820), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n613), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n836), .B2(new_n829), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n831), .B1(new_n825), .B2(new_n837), .ZN(G1344gat));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n817), .B2(new_n818), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n826), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n815), .A2(KEYINPUT121), .A3(new_n792), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n714), .B1(new_n813), .B2(new_n789), .ZN(new_n845));
  NOR4_X1   g644(.A1(new_n240), .A2(new_n296), .A3(new_n359), .A4(new_n693), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n552), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n848), .A2(new_n849), .A3(new_n818), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n848), .B2(new_n818), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n842), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n852), .A2(KEYINPUT59), .A3(new_n359), .A4(new_n822), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n823), .A2(new_n734), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(KEYINPUT59), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n836), .A2(new_n734), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(G148gat), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n855), .A2(G148gat), .B1(new_n857), .B2(KEYINPUT59), .ZN(G1345gat));
  NOR3_X1   g657(.A1(new_n823), .A2(new_n388), .A3(new_n240), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n836), .A2(new_n240), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n388), .B2(new_n860), .ZN(G1346gat));
  NOR3_X1   g660(.A1(new_n823), .A2(new_n389), .A3(new_n648), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n836), .A2(new_n648), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n389), .B2(new_n863), .ZN(G1347gat));
  NOR2_X1   g663(.A1(new_n613), .A2(new_n606), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n791), .B2(new_n792), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n867), .A2(new_n614), .A3(new_n603), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n335), .B1(new_n476), .B2(new_n477), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(new_n614), .A3(new_n707), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n871), .A2(new_n335), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n872), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT123), .B1(new_n872), .B2(G169gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT124), .ZN(G1348gat));
  AOI21_X1  g675(.A(G176gat), .B1(new_n868), .B2(new_n359), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n871), .A2(new_n354), .A3(new_n734), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(G1349gat));
  AND2_X1   g678(.A1(new_n714), .A2(new_n455), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT125), .B1(new_n868), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G183gat), .B1(new_n871), .B2(new_n240), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n871), .B2(new_n648), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT61), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n456), .A3(new_n296), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1351gat));
  NOR2_X1   g687(.A1(new_n639), .A2(new_n866), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n817), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(G197gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n693), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n848), .A2(new_n818), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT122), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n848), .A2(new_n849), .A3(new_n818), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n895), .A2(new_n896), .B1(new_n840), .B2(new_n841), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(new_n335), .A3(new_n890), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n893), .B1(new_n898), .B2(new_n892), .ZN(G1352gat));
  NAND3_X1  g698(.A1(new_n891), .A2(new_n356), .A3(new_n359), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n900), .B(KEYINPUT62), .Z(new_n901));
  NOR3_X1   g700(.A1(new_n897), .A2(new_n734), .A3(new_n890), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n356), .ZN(G1353gat));
  INV_X1    g702(.A(new_n891), .ZN(new_n904));
  OR3_X1    g703(.A1(new_n904), .A2(new_n492), .A3(new_n240), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n852), .A2(new_n714), .A3(new_n889), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n906), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT63), .B1(new_n906), .B2(G211gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(G1354gat));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n897), .B2(new_n890), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n296), .A2(G218gat), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT127), .Z(new_n913));
  NAND3_X1  g712(.A1(new_n852), .A2(KEYINPUT126), .A3(new_n889), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(G218gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n904), .B2(new_n648), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n915), .A2(new_n917), .ZN(G1355gat));
endmodule


