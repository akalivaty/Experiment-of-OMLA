//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n209), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT64), .Z(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT65), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n209), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT0), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n201), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI22_X1  g0033(.A1(new_n226), .A2(KEYINPUT0), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  AND4_X1   g0034(.A1(new_n221), .A2(new_n223), .A3(new_n227), .A4(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  INV_X1    g0037(.A(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n212), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n239), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT69), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT68), .B(G264), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT70), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(KEYINPUT70), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n228), .A3(new_n259), .ZN(new_n260));
  XOR2_X1   g0060(.A(KEYINPUT15), .B(G87), .Z(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n229), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT8), .B(G58), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G77), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n265), .A2(new_n267), .B1(new_n229), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n260), .B1(new_n264), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G13), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n271), .A2(new_n229), .A3(G1), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n268), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n229), .A2(G1), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n260), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n270), .B(new_n273), .C1(new_n268), .C2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G107), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  OAI221_X1 g0083(.A(new_n280), .B1(new_n281), .B2(new_n214), .C1(new_n212), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(G41), .B2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n286), .A2(new_n290), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(G244), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n277), .B1(new_n296), .B2(G169), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n295), .A2(G179), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n277), .B1(new_n296), .B2(G190), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n295), .A2(G200), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  XOR2_X1   g0104(.A(new_n304), .B(KEYINPUT71), .Z(new_n305));
  INV_X1    g0105(.A(KEYINPUT7), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n278), .B2(G20), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT3), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(G33), .ZN(new_n309));
  INV_X1    g0109(.A(G33), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n311));
  OAI211_X1 g0111(.A(KEYINPUT7), .B(new_n229), .C1(new_n309), .C2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n307), .A2(KEYINPUT73), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT73), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(new_n306), .C1(new_n278), .C2(G20), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(G68), .A3(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n211), .A2(new_n213), .ZN(new_n317));
  OAI21_X1  g0117(.A(G20), .B1(new_n317), .B2(new_n201), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n266), .A2(G159), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT16), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n260), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n307), .A2(new_n312), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n320), .B1(new_n326), .B2(G68), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(new_n327), .B2(KEYINPUT16), .ZN(new_n328));
  INV_X1    g0128(.A(new_n265), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n276), .A2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n329), .A2(new_n272), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n324), .A2(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT17), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n333), .A2(KEYINPUT74), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n308), .A2(G33), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n335), .A2(new_n336), .A3(G226), .A4(G1698), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(G223), .A4(new_n282), .ZN(new_n338));
  INV_X1    g0138(.A(G87), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n337), .B(new_n338), .C1(new_n310), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n287), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n292), .B1(new_n293), .B2(G232), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n341), .A2(G190), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G200), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(new_n341), .B2(new_n342), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n333), .A2(KEYINPUT74), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n332), .A2(new_n334), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n330), .A2(new_n331), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT16), .B1(new_n316), .B2(new_n321), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n327), .A2(KEYINPUT16), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n260), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n346), .B(new_n349), .C1(new_n350), .C2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(KEYINPUT74), .A3(new_n333), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n349), .B1(new_n352), .B2(new_n350), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n341), .B2(new_n342), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n341), .A2(new_n342), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n357), .B1(G179), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n355), .A2(new_n360), .A3(KEYINPUT18), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT18), .B1(new_n355), .B2(new_n360), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n348), .B(new_n354), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n266), .A2(G50), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n364), .B1(new_n229), .B2(G68), .C1(new_n268), .C2(new_n263), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n365), .A2(new_n260), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n366), .A2(KEYINPUT11), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n272), .A2(new_n213), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT12), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n275), .A2(G68), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(KEYINPUT11), .A3(new_n260), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n367), .A2(new_n369), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  XOR2_X1   g0172(.A(new_n372), .B(KEYINPUT72), .Z(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G97), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n283), .B2(new_n238), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n281), .A2(new_n212), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n287), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT13), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n292), .B1(new_n293), .B2(G238), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n378), .B1(new_n377), .B2(new_n379), .ZN(new_n382));
  OAI21_X1  g0182(.A(G200), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n381), .A2(new_n382), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G190), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n373), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT14), .B1(new_n384), .B2(new_n356), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT14), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(G169), .C1(new_n381), .C2(new_n382), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n384), .A2(G179), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n372), .B(KEYINPUT72), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n203), .A2(G20), .ZN(new_n395));
  INV_X1    g0195(.A(G150), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n395), .B1(new_n396), .B2(new_n267), .C1(new_n265), .C2(new_n263), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n260), .B1(new_n202), .B2(new_n272), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n275), .A2(G50), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n293), .A2(G226), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n291), .B2(new_n290), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n278), .A2(G222), .A3(new_n282), .ZN(new_n404));
  INV_X1    g0204(.A(G223), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n404), .B1(new_n268), .B2(new_n278), .C1(new_n281), .C2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n403), .B1(new_n406), .B2(new_n287), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n401), .A2(KEYINPUT9), .B1(new_n344), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n407), .ZN(new_n409));
  INV_X1    g0209(.A(G190), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT9), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n409), .A2(new_n410), .B1(new_n400), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT10), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n401), .A2(KEYINPUT9), .B1(new_n407), .B2(G190), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n409), .A2(G200), .B1(new_n400), .B2(new_n411), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT10), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n409), .A2(G179), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n400), .B1(new_n407), .B2(G169), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NOR4_X1   g0222(.A1(new_n305), .A2(new_n363), .A3(new_n394), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G283), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n335), .A2(new_n336), .A3(G250), .A4(G1698), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n335), .A2(new_n336), .A3(G244), .A4(new_n282), .ZN(new_n426));
  NOR2_X1   g0226(.A1(KEYINPUT77), .A2(KEYINPUT4), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n424), .B(new_n425), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n426), .A2(new_n427), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n287), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT78), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(KEYINPUT78), .B(new_n287), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G45), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(G1), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT5), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G41), .ZN(new_n438));
  INV_X1    g0238(.A(G41), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT5), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(G257), .A3(new_n286), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n436), .A2(new_n438), .A3(new_n440), .A4(G274), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n434), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G200), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n313), .A2(G107), .A3(new_n315), .ZN(new_n448));
  AND2_X1   g0248(.A1(G97), .A2(G107), .ZN(new_n449));
  NOR2_X1   g0249(.A1(G97), .A2(G107), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n449), .A2(new_n450), .B1(KEYINPUT75), .B2(KEYINPUT6), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G97), .A2(G107), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n207), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n325), .B1(new_n448), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n272), .A2(new_n205), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT76), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n459), .B(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n274), .A2(G13), .B1(new_n289), .B2(G33), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n325), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n463), .B2(new_n205), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n426), .A2(new_n427), .ZN(new_n466));
  INV_X1    g0266(.A(new_n427), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n278), .A2(G244), .A3(new_n282), .A4(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n466), .A2(new_n468), .A3(new_n424), .A4(new_n425), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n444), .B1(new_n469), .B2(new_n287), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G190), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n447), .A2(new_n465), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G179), .ZN(new_n473));
  INV_X1    g0273(.A(new_n433), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT78), .B1(new_n469), .B2(new_n287), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n473), .B(new_n445), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT79), .ZN(new_n477));
  AOI21_X1  g0277(.A(G169), .B1(new_n430), .B2(new_n445), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n448), .A2(new_n457), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n260), .ZN(new_n480));
  INV_X1    g0280(.A(new_n464), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT79), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n434), .A2(new_n483), .A3(new_n473), .A4(new_n445), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n477), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT80), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n477), .A2(new_n482), .A3(new_n484), .A4(KEYINPUT80), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n472), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(G303), .B1(new_n309), .B2(new_n311), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n335), .A2(new_n336), .A3(G257), .A4(new_n282), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n335), .A2(new_n336), .A3(G264), .A4(G1698), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n287), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n289), .B(G45), .C1(new_n437), .C2(G41), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n439), .A2(KEYINPUT5), .ZN(new_n496));
  OAI211_X1 g0296(.A(G270), .B(new_n286), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n497), .A2(new_n443), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n356), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n256), .A2(new_n257), .B1(G1), .B2(G13), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n462), .A2(G116), .A3(new_n259), .A4(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G116), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n272), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(G20), .B1(G33), .B2(G283), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n310), .A2(G97), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n504), .A2(new_n505), .B1(G20), .B2(new_n502), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n260), .A2(KEYINPUT20), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT20), .B1(new_n260), .B2(new_n506), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n501), .B(new_n503), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n499), .A2(new_n509), .A3(KEYINPUT21), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n497), .A2(new_n443), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n287), .B2(new_n493), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n509), .A2(G179), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT21), .B1(new_n499), .B2(new_n509), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n229), .B1(new_n374), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(G87), .B2(new_n207), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n335), .A2(new_n336), .A3(new_n229), .A4(G68), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n517), .B1(new_n263), .B2(new_n205), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n260), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n325), .A2(new_n261), .A3(new_n462), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n262), .A2(new_n272), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n335), .A2(new_n336), .A3(G244), .A4(G1698), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT83), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n278), .A2(KEYINPUT83), .A3(G244), .A4(G1698), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n278), .A2(G238), .A3(new_n282), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n529), .A2(new_n530), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n287), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n436), .A2(G274), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT81), .B1(new_n435), .B2(G1), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT81), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n289), .A3(G45), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g0339(.A1(G33), .A2(G41), .ZN(new_n540));
  OAI21_X1  g0340(.A(G250), .B1(new_n540), .B2(new_n228), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n535), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n544), .B(new_n535), .C1(new_n539), .C2(new_n541), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n534), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n526), .B1(new_n356), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n534), .A2(new_n546), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n473), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n325), .A2(G87), .A3(new_n462), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n523), .A2(new_n525), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n547), .B2(G200), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n534), .A2(new_n546), .A3(G190), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n494), .A2(new_n498), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G200), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n501), .A2(new_n503), .ZN(new_n559));
  INV_X1    g0359(.A(new_n507), .ZN(new_n560));
  INV_X1    g0360(.A(new_n508), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT84), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n558), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n512), .A2(G190), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n344), .B1(new_n494), .B2(new_n498), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT84), .B1(new_n566), .B2(new_n509), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n516), .A2(new_n551), .A3(new_n556), .A4(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT86), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT25), .ZN(new_n571));
  INV_X1    g0371(.A(new_n272), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(G107), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n272), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n463), .B2(new_n206), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n278), .A2(new_n229), .A3(G87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT22), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT22), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n278), .A2(new_n579), .A3(new_n229), .A4(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT23), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n229), .B2(G107), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(G20), .B2(new_n531), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT24), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n325), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n589), .B(new_n586), .C1(new_n578), .C2(new_n580), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n576), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n278), .A2(G250), .A3(new_n282), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n278), .A2(G257), .A3(G1698), .ZN(new_n595));
  XNOR2_X1  g0395(.A(KEYINPUT85), .B(G294), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G33), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n287), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n441), .A2(G264), .A3(new_n286), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n443), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n356), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n599), .A2(new_n473), .A3(new_n600), .A4(new_n443), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n593), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(G200), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n599), .A2(G190), .A3(new_n600), .A4(new_n443), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n576), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n586), .B1(new_n578), .B2(new_n580), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n260), .B1(new_n610), .B2(KEYINPUT24), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n609), .B1(new_n611), .B2(new_n591), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n570), .B1(new_n605), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n602), .A3(new_n603), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(KEYINPUT86), .C1(new_n612), .C2(new_n608), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n569), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n423), .A2(new_n489), .A3(new_n617), .ZN(G372));
  NAND2_X1  g0418(.A1(new_n487), .A2(new_n488), .ZN(new_n619));
  INV_X1    g0419(.A(new_n472), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n516), .A2(new_n615), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n551), .A2(new_n556), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(new_n613), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n619), .A2(new_n620), .A3(new_n621), .A4(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT87), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n489), .A2(KEYINPUT87), .A3(new_n621), .A4(new_n623), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n458), .A2(new_n464), .B1(G169), .B2(new_n470), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(KEYINPUT79), .B2(new_n476), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n548), .A2(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .A4(new_n484), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n551), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n487), .A2(new_n488), .A3(new_n630), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(KEYINPUT26), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n626), .A2(new_n627), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n423), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n361), .A2(new_n362), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n386), .A2(new_n348), .A3(new_n354), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n299), .B1(new_n391), .B2(new_n392), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n418), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n421), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n637), .A2(new_n644), .ZN(G369));
  NOR2_X1   g0445(.A1(new_n271), .A2(G20), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n289), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n562), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n516), .A2(new_n568), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT88), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n654), .B1(new_n514), .B2(new_n515), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G330), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n614), .A2(new_n616), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n593), .B2(new_n653), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n615), .A2(new_n653), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n516), .A2(new_n652), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n614), .B2(new_n616), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n605), .B2(new_n653), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(G399));
  INV_X1    g0473(.A(new_n224), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G1), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n232), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT29), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n636), .A2(new_n681), .A3(new_n653), .ZN(new_n682));
  INV_X1    g0482(.A(new_n624), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT26), .B1(new_n622), .B2(new_n485), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n551), .B(new_n684), .C1(new_n634), .C2(KEYINPUT26), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n653), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT29), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n489), .A2(new_n617), .A3(new_n653), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n557), .A2(new_n473), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n549), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n470), .A2(new_n599), .A3(new_n600), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n601), .A2(new_n473), .A3(new_n557), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n446), .A2(new_n694), .A3(new_n547), .ZN(new_n695));
  INV_X1    g0495(.A(new_n692), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(KEYINPUT30), .A3(new_n690), .A4(new_n549), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT31), .B1(new_n698), .B2(new_n652), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n688), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n682), .A2(new_n687), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n680), .B1(new_n705), .B2(G1), .ZN(G364));
  NOR2_X1   g0506(.A1(new_n660), .A2(G330), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT89), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT90), .B1(new_n646), .B2(G45), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n289), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n646), .A2(KEYINPUT90), .A3(G45), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n675), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n707), .A2(KEYINPUT89), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n708), .A2(new_n661), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n278), .A2(new_n224), .ZN(new_n717));
  INV_X1    g0517(.A(G355), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(G116), .B2(new_n224), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n251), .A2(new_n435), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n279), .A2(new_n224), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n435), .B2(new_n233), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n719), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G13), .A2(G33), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n228), .B1(G20), .B2(new_n356), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n713), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n229), .A2(new_n410), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n344), .A2(G179), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n339), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n229), .A2(new_n473), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G190), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n229), .A2(G190), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n732), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n737), .A2(new_n268), .B1(new_n739), .B2(new_n206), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n735), .A2(G190), .A3(new_n344), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n734), .B(new_n740), .C1(G58), .C2(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n410), .A2(G179), .A3(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n229), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n205), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n473), .A2(new_n344), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n738), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n279), .B(new_n746), .C1(G68), .C2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n738), .A2(new_n473), .A3(new_n344), .ZN(new_n751));
  INV_X1    g0551(.A(G159), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT32), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT91), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n747), .A2(new_n731), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n755), .B1(new_n747), .B2(new_n731), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G50), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n743), .A2(new_n750), .A3(new_n754), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(G326), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT33), .B(G317), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n742), .A2(G322), .B1(new_n749), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n751), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n765), .A2(KEYINPUT93), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(KEYINPUT93), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G329), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n762), .B1(KEYINPUT94), .B2(new_n764), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n764), .A2(KEYINPUT94), .ZN(new_n771));
  INV_X1    g0571(.A(G311), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n737), .A2(new_n772), .B1(new_n739), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n745), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(new_n596), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G303), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n279), .B1(new_n733), .B2(new_n777), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT92), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT92), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n771), .A2(new_n776), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n761), .B1(new_n770), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n730), .B1(new_n782), .B2(new_n727), .ZN(new_n783));
  INV_X1    g0583(.A(new_n726), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n660), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n716), .A2(new_n785), .ZN(G396));
  NAND2_X1  g0586(.A1(new_n636), .A2(new_n653), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n277), .A2(new_n652), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n303), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n300), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n299), .A2(new_n653), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n792), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n636), .A2(new_n653), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n713), .B1(new_n796), .B2(new_n703), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n703), .B2(new_n796), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n727), .A2(new_n724), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n714), .B1(new_n268), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n727), .ZN(new_n801));
  INV_X1    g0601(.A(new_n737), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n742), .A2(G143), .B1(new_n802), .B2(G159), .ZN(new_n803));
  INV_X1    g0603(.A(G137), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n396), .B2(new_n748), .C1(new_n804), .C2(new_n758), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT34), .ZN(new_n806));
  INV_X1    g0606(.A(new_n733), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n279), .B1(new_n807), .B2(G50), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n808), .B1(new_n211), .B2(new_n745), .C1(new_n213), .C2(new_n739), .ZN(new_n809));
  INV_X1    g0609(.A(new_n768), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(G132), .B2(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G116), .A2(new_n802), .B1(new_n807), .B2(G107), .ZN(new_n812));
  INV_X1    g0612(.A(G294), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n773), .B2(new_n748), .C1(new_n813), .C2(new_n741), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n739), .A2(new_n339), .ZN(new_n815));
  NOR4_X1   g0615(.A1(new_n814), .A2(new_n278), .A3(new_n746), .A4(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n810), .A2(G311), .B1(G303), .B2(new_n759), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n806), .A2(new_n811), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n800), .B1(new_n801), .B2(new_n818), .C1(new_n794), .C2(new_n725), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n798), .A2(new_n819), .ZN(G384));
  OR2_X1    g0620(.A1(new_n456), .A2(KEYINPUT35), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n456), .A2(KEYINPUT35), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n821), .A2(G116), .A3(new_n230), .A4(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT36), .Z(new_n824));
  OR3_X1    g0624(.A1(new_n232), .A2(new_n268), .A3(new_n317), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n202), .A2(G68), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n289), .B(G13), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n702), .A2(KEYINPUT97), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT97), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n688), .A2(new_n701), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT40), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n392), .A2(new_n652), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n386), .A2(new_n393), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n391), .A2(new_n392), .A3(new_n652), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n794), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n829), .B2(new_n831), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n324), .A2(new_n328), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n359), .B1(new_n840), .B2(new_n349), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT95), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT37), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n650), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n355), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n355), .A2(new_n360), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT95), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n843), .A2(new_n353), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n846), .A2(new_n845), .A3(new_n353), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n363), .A2(new_n355), .A3(new_n844), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT96), .ZN(new_n855));
  INV_X1    g0655(.A(new_n353), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n328), .B1(KEYINPUT16), .B2(new_n327), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(new_n349), .B1(new_n359), .B2(new_n650), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT37), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n650), .B1(new_n857), .B2(new_n349), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n848), .A2(new_n859), .B1(new_n363), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n855), .B1(new_n861), .B2(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n363), .A2(new_n860), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n353), .B(new_n845), .C1(new_n841), .C2(new_n842), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n846), .B2(KEYINPUT95), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n859), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n863), .A2(new_n855), .A3(new_n867), .A4(KEYINPUT38), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n854), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n833), .B1(new_n839), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n792), .B1(new_n835), .B2(new_n836), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n688), .A2(new_n830), .A3(new_n701), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n830), .B1(new_n688), .B2(new_n701), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n863), .A2(new_n867), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n863), .A2(KEYINPUT38), .A3(new_n867), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n833), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n423), .B(new_n832), .C1(new_n871), .C2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(G330), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n879), .A2(KEYINPUT96), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n853), .B1(new_n885), .B2(new_n868), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT40), .B1(new_n875), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n832), .A2(new_n833), .A3(new_n880), .A4(new_n872), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n884), .B1(new_n829), .B2(new_n831), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n423), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n883), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n682), .A2(new_n687), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n423), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n644), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n893), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n795), .A2(new_n791), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(new_n880), .A3(new_n837), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n638), .A2(new_n844), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n393), .A2(new_n652), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n878), .B2(new_n879), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n886), .B2(new_n903), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n899), .B(new_n900), .C1(new_n902), .C2(new_n905), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n897), .A2(new_n906), .B1(new_n289), .B2(new_n646), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n897), .A2(new_n906), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n828), .B1(new_n907), .B2(new_n908), .ZN(G367));
  INV_X1    g0709(.A(new_n712), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT102), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n664), .A2(new_n666), .A3(new_n670), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT100), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n662), .A2(KEYINPUT101), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT101), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n671), .B1(new_n661), .B2(new_n916), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n915), .B1(new_n914), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n911), .B1(new_n920), .B2(new_n704), .ZN(new_n921));
  OAI211_X1 g0721(.A(KEYINPUT102), .B(new_n705), .C1(new_n918), .C2(new_n919), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n489), .B1(new_n465), .B2(new_n653), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n629), .A2(new_n484), .A3(new_n652), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n926), .A2(new_n672), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT44), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n672), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT45), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n929), .B(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n928), .A2(new_n668), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n668), .B1(new_n928), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT103), .B1(new_n923), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT103), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n934), .A2(new_n921), .A3(new_n937), .A4(new_n922), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n704), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n675), .B(KEYINPUT41), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n910), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n671), .A2(new_n489), .A3(new_n621), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT42), .ZN(new_n944));
  INV_X1    g0744(.A(new_n926), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n619), .B1(new_n945), .B2(new_n615), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n944), .B1(new_n946), .B2(new_n653), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n553), .A2(new_n652), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n551), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n630), .B2(new_n948), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT43), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT98), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n952), .A2(KEYINPUT98), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n947), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT99), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n950), .A2(new_n952), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n947), .A2(new_n955), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n668), .A2(new_n945), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n942), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n247), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n728), .B1(new_n224), .B2(new_n262), .C1(new_n966), .C2(new_n721), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n713), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n739), .A2(new_n268), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n278), .B1(new_n751), .B2(new_n804), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(G159), .C2(new_n749), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n775), .A2(G68), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n759), .A2(G143), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n202), .A2(new_n737), .B1(new_n733), .B2(new_n211), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G150), .B2(new_n742), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT104), .B(G317), .Z(new_n977));
  AOI21_X1  g0777(.A(new_n278), .B1(new_n765), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n205), .B2(new_n739), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT105), .Z(new_n980));
  OAI22_X1  g0780(.A1(new_n741), .A2(new_n777), .B1(new_n737), .B2(new_n773), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n596), .B2(new_n749), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n807), .A2(KEYINPUT46), .A3(G116), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT46), .B1(new_n807), .B2(G116), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G107), .B2(new_n775), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n759), .A2(G311), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n982), .A2(new_n983), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n976), .B1(new_n980), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT47), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n801), .B1(new_n988), .B2(new_n989), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n968), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n950), .A2(new_n726), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n965), .A2(new_n994), .ZN(G387));
  XOR2_X1   g0795(.A(new_n675), .B(KEYINPUT109), .Z(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n920), .B2(new_n704), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n923), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n242), .A2(new_n435), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n999), .A2(new_n721), .B1(new_n677), .B2(new_n717), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n265), .B2(G50), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n329), .A2(new_n1001), .A3(new_n202), .ZN(new_n1004));
  AOI21_X1  g0804(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1003), .A2(new_n677), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1000), .A2(new_n1006), .B1(new_n206), .B2(new_n674), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n713), .B1(new_n1007), .B2(new_n729), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n807), .A2(G77), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n213), .B2(new_n737), .C1(new_n396), .C2(new_n751), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G159), .B2(new_n759), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n741), .A2(new_n202), .B1(new_n748), .B2(new_n265), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n739), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n279), .B(new_n1012), .C1(G97), .C2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1011), .B(new_n1014), .C1(new_n262), .C2(new_n745), .ZN(new_n1015));
  INV_X1    g0815(.A(G322), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n758), .A2(new_n1016), .B1(new_n772), .B2(new_n748), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT107), .Z(new_n1018));
  AOI22_X1  g0818(.A1(new_n742), .A2(new_n977), .B1(new_n802), .B2(G303), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT48), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n775), .A2(G283), .B1(new_n807), .B2(new_n596), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n278), .B1(new_n765), .B2(G326), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n502), .C2(new_n739), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1023), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1015), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1008), .B1(new_n1028), .B2(new_n727), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n667), .B2(new_n784), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n998), .B(new_n1030), .C1(new_n910), .C2(new_n920), .ZN(G393));
  NAND2_X1  g0831(.A1(new_n936), .A2(new_n938), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n996), .B1(new_n923), .B2(new_n935), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n945), .A2(new_n726), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n254), .A2(new_n721), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n728), .B1(new_n205), .B2(new_n224), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n713), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n759), .A2(G150), .B1(G159), .B2(new_n742), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G143), .A2(new_n765), .B1(new_n749), .B2(G50), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n329), .A2(new_n802), .B1(new_n807), .B2(G68), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n745), .A2(new_n268), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1044), .A2(new_n279), .A3(new_n815), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n759), .A2(G317), .B1(G311), .B2(new_n742), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(KEYINPUT52), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n279), .B1(new_n739), .B2(new_n206), .C1(new_n745), .C2(new_n502), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1016), .A2(new_n751), .B1(new_n737), .B2(new_n813), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n773), .A2(new_n733), .B1(new_n748), .B2(new_n777), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1048), .A2(KEYINPUT52), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1046), .A2(new_n1047), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1038), .B1(new_n1056), .B2(new_n727), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n934), .A2(new_n712), .B1(new_n1035), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1034), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT111), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1034), .A2(KEYINPUT111), .A3(new_n1058), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(G390));
  INV_X1    g0863(.A(new_n837), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n795), .B2(new_n791), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n905), .B1(new_n1065), .B2(new_n901), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n653), .B(new_n790), .C1(new_n683), .C2(new_n685), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1067), .A2(new_n791), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT112), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n837), .B(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n902), .B(new_n870), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n890), .A2(new_n872), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n872), .A2(new_n702), .A3(G330), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1066), .A2(new_n1071), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1064), .B1(new_n703), .B2(new_n792), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1073), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n898), .ZN(new_n1081));
  OAI211_X1 g0881(.A(G330), .B(new_n794), .C1(new_n873), .C2(new_n874), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1070), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT113), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1076), .A2(new_n1067), .A3(new_n791), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1084), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1081), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n896), .A2(new_n892), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1078), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n996), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1075), .A2(new_n1088), .A3(new_n1077), .A4(new_n1089), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n714), .B1(new_n265), .B2(new_n799), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n742), .A2(G116), .B1(new_n1013), .B2(G68), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n205), .B2(new_n737), .C1(new_n206), .C2(new_n748), .ZN(new_n1097));
  NOR4_X1   g0897(.A1(new_n1097), .A2(new_n278), .A3(new_n734), .A4(new_n1044), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n810), .A2(G294), .B1(G283), .B2(new_n759), .ZN(new_n1099));
  INV_X1    g0899(.A(G128), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n758), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n742), .A2(G132), .B1(new_n1013), .B2(G50), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n804), .B2(new_n748), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(G125), .C2(new_n810), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n278), .B1(new_n737), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n733), .A2(new_n396), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1106), .B(new_n1109), .C1(G159), .C2(new_n775), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1098), .A2(new_n1099), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1095), .B1(new_n1111), .B2(new_n801), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n905), .B2(new_n724), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1078), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n712), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1094), .A2(new_n1115), .ZN(G378));
  INV_X1    g0916(.A(KEYINPUT119), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n401), .A2(new_n650), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n418), .A2(new_n421), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n418), .B2(new_n421), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1119), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1124), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n1122), .A3(new_n1118), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n889), .A2(new_n1131), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1125), .A2(new_n1128), .A3(KEYINPUT117), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT117), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n884), .B(new_n1135), .C1(new_n887), .C2(new_n888), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1132), .A2(new_n1136), .A3(new_n906), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n900), .B1(new_n905), .B2(new_n902), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n878), .A2(new_n879), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1064), .B(new_n1139), .C1(new_n795), .C2(new_n791), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(G330), .B1(new_n871), .B2(new_n882), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1130), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1135), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n889), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1141), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1117), .B1(new_n1137), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1093), .A2(new_n1089), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n906), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1143), .A2(new_n1145), .A3(new_n1141), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n1150), .A3(KEYINPUT119), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT120), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1137), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1149), .A2(new_n1150), .A3(KEYINPUT120), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1148), .A2(new_n1156), .A3(KEYINPUT57), .A4(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1154), .A2(new_n1092), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1147), .A2(new_n712), .A3(new_n1151), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n714), .B1(new_n202), .B2(new_n799), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n972), .A2(new_n439), .A3(new_n279), .A4(new_n1009), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n262), .A2(new_n737), .B1(new_n206), .B2(new_n741), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n748), .A2(new_n205), .B1(new_n739), .B2(new_n211), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n502), .B2(new_n758), .C1(new_n773), .C2(new_n768), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT58), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(G33), .A2(G41), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(G50), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n278), .B2(G41), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n804), .A2(new_n737), .B1(new_n733), .B2(new_n1105), .ZN(new_n1171));
  INV_X1    g0971(.A(G132), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n741), .A2(new_n1100), .B1(new_n748), .B2(new_n1172), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(G150), .C2(new_n775), .ZN(new_n1174));
  INV_X1    g0974(.A(G125), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n758), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT59), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT115), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1178), .A2(G124), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(G124), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n765), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n1168), .C1(new_n752), .C2(new_n739), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1167), .B(new_n1170), .C1(new_n1177), .C2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1183), .A2(KEYINPUT116), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(KEYINPUT116), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n727), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1161), .B1(new_n1184), .B2(new_n1186), .C1(new_n1144), .C2(new_n725), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT118), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1160), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1159), .A2(new_n1190), .ZN(G375));
  INV_X1    g0991(.A(new_n1088), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1089), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(new_n940), .A3(new_n1090), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1070), .A2(new_n724), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n727), .A2(G68), .A3(new_n724), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n768), .A2(new_n777), .B1(new_n813), .B2(new_n758), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G107), .A2(new_n802), .B1(new_n807), .B2(G97), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n502), .B2(new_n748), .C1(new_n773), .C2(new_n741), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n279), .B1(new_n739), .B2(new_n268), .C1(new_n745), .C2(new_n262), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT121), .Z(new_n1203));
  OAI221_X1 g1003(.A(new_n278), .B1(new_n739), .B2(new_n211), .C1(new_n745), .C2(new_n202), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n741), .A2(new_n804), .B1(new_n737), .B2(new_n396), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n752), .A2(new_n733), .B1(new_n748), .B2(new_n1105), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n1172), .B2(new_n758), .C1(new_n1100), .C2(new_n768), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1203), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(KEYINPUT122), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n801), .B1(new_n1209), .B2(KEYINPUT122), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n714), .B(new_n1197), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1088), .A2(new_n712), .B1(new_n1196), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1195), .A2(new_n1214), .ZN(G381));
  INV_X1    g1015(.A(G378), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1159), .A2(new_n1216), .A3(new_n1190), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1034), .A2(KEYINPUT111), .A3(new_n1058), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT111), .B1(new_n1034), .B2(new_n1058), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n942), .A2(new_n964), .B1(new_n993), .B2(new_n992), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1217), .B1(new_n1223), .B2(KEYINPUT123), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(KEYINPUT123), .B2(new_n1223), .ZN(G407));
  OAI211_X1 g1025(.A(G407), .B(G213), .C1(G343), .C2(new_n1217), .ZN(G409));
  INV_X1    g1026(.A(KEYINPUT60), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1194), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n996), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT124), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1194), .B2(new_n1227), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1192), .A2(KEYINPUT124), .A3(KEYINPUT60), .A4(new_n1193), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1230), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1214), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n798), .B(new_n819), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G384), .B(new_n1214), .C1(new_n1237), .C2(new_n1230), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n651), .A2(G213), .A3(G2897), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G375), .A2(G378), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1156), .A2(new_n712), .A3(new_n1157), .ZN(new_n1244));
  AND4_X1   g1044(.A1(new_n1094), .A2(new_n1244), .A3(new_n1115), .A4(new_n1187), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1152), .A2(new_n941), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1245), .A2(new_n1246), .B1(G213), .B2(new_n651), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT61), .B1(new_n1242), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1250));
  OR3_X1    g1050(.A1(new_n1248), .A2(KEYINPUT62), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1250), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(new_n1243), .A3(new_n1247), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT62), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1249), .A2(new_n1251), .A3(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT125), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1220), .B2(G387), .ZN(new_n1257));
  XOR2_X1   g1057(.A(G393), .B(G396), .Z(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1220), .A2(G387), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G390), .A2(new_n1221), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1257), .A2(new_n1259), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1220), .A2(G387), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G390), .A2(new_n1221), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1256), .A4(new_n1258), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1255), .A2(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT63), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1253), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1253), .A2(new_n1269), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1268), .A2(new_n1270), .A3(new_n1271), .A4(new_n1249), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1267), .A2(new_n1272), .ZN(G405));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1243), .A2(new_n1274), .A3(new_n1217), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n996), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1276));
  AOI211_X1 g1076(.A(G378), .B(new_n1189), .C1(new_n1276), .C2(new_n1158), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1216), .B1(new_n1159), .B2(new_n1190), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT126), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1275), .A2(new_n1279), .A3(new_n1252), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1250), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT127), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1275), .A2(new_n1279), .A3(new_n1282), .A4(new_n1252), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1284), .A2(new_n1266), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1266), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(G402));
endmodule


