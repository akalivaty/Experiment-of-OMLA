//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1224, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0005(.A(KEYINPUT65), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n206), .B1(new_n207), .B2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n209), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AND2_X1   g0013(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n207), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n202), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR4_X1   g0030(.A1(new_n214), .A2(new_n215), .A3(new_n226), .A4(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n217), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n243), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n229), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n251), .A2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G50), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G50), .B2(new_n252), .ZN(new_n259));
  INV_X1    g0059(.A(new_n255), .ZN(new_n260));
  XOR2_X1   g0060(.A(KEYINPUT8), .B(G58), .Z(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n228), .A2(new_n262), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n261), .A2(new_n263), .B1(G150), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n260), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n259), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g0069(.A(new_n269), .B(KEYINPUT9), .Z(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  AND2_X1   g0071(.A1(G1), .A2(G13), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G226), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n278), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G222), .ZN(new_n288));
  INV_X1    g0088(.A(G77), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n262), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G223), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(G1698), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n288), .B1(new_n289), .B2(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n283), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G190), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n298), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n270), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n299), .B(KEYINPUT69), .C1(new_n300), .C2(new_n298), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n303), .C1(new_n270), .C2(new_n301), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(new_n269), .C1(G169), .C2(new_n298), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n263), .A2(G77), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n313), .B1(new_n228), .B2(G68), .C1(new_n244), .C2(new_n264), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n255), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT71), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT11), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n317), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT12), .B1(new_n252), .B2(G68), .ZN(new_n320));
  OR3_X1    g0120(.A1(new_n252), .A2(KEYINPUT12), .A3(G68), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n217), .B1(new_n251), .B2(G20), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n320), .A2(new_n321), .B1(new_n256), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n318), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n293), .A2(G232), .A3(G1698), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT70), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT70), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n293), .A2(new_n327), .A3(G232), .A4(G1698), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n287), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n297), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n278), .B1(new_n218), .B2(new_n282), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n280), .B1(new_n329), .B2(new_n330), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT13), .B1(new_n337), .B2(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT14), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(G169), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(G179), .A3(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n340), .B1(new_n339), .B2(G169), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n324), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n318), .A2(new_n319), .A3(new_n323), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n339), .A2(G200), .ZN(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n346), .B(new_n347), .C1(new_n348), .C2(new_n339), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n256), .A2(G77), .A3(new_n257), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(G77), .B2(new_n252), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n261), .A2(new_n265), .B1(G20), .B2(G77), .ZN(new_n353));
  XOR2_X1   g0153(.A(KEYINPUT15), .B(G87), .Z(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n263), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n260), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G244), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n278), .B1(new_n359), .B2(new_n282), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n287), .A2(G232), .ZN(new_n361));
  INV_X1    g0161(.A(G107), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n361), .B1(new_n362), .B2(new_n293), .C1(new_n218), .C2(new_n295), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n360), .B1(new_n363), .B2(new_n297), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n358), .B1(new_n364), .B2(G190), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n300), .B2(new_n364), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n309), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(new_n358), .C1(G169), .C2(new_n364), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT68), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT7), .B1(new_n286), .B2(new_n228), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n291), .A2(KEYINPUT7), .A3(new_n228), .A4(new_n292), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(G68), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G58), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(new_n217), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(new_n201), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(KEYINPUT16), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT72), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT72), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n374), .A2(new_n381), .A3(new_n378), .A4(KEYINPUT16), .ZN(new_n382));
  XOR2_X1   g0182(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n383));
  NAND3_X1  g0183(.A1(new_n291), .A2(new_n228), .A3(new_n292), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n217), .B1(new_n386), .B2(new_n372), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n376), .A2(new_n201), .ZN(new_n388));
  INV_X1    g0188(.A(G159), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n388), .A2(new_n228), .B1(new_n389), .B2(new_n264), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n383), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n380), .A2(new_n255), .A3(new_n382), .A4(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n261), .A2(new_n257), .ZN(new_n393));
  INV_X1    g0193(.A(new_n261), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n393), .A2(new_n256), .B1(new_n253), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n282), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(G232), .B1(new_n274), .B2(new_n277), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n279), .A2(G1698), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n399), .B1(G223), .B2(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G87), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n398), .B(G179), .C1(new_n402), .C2(new_n280), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n280), .B1(new_n400), .B2(new_n401), .ZN(new_n404));
  INV_X1    g0204(.A(G232), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n278), .B1(new_n405), .B2(new_n282), .ZN(new_n406));
  OAI21_X1  g0206(.A(G169), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n403), .A2(KEYINPUT74), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT74), .B1(new_n403), .B2(new_n407), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n396), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT18), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n404), .A2(new_n406), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n348), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(G200), .B2(new_n413), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n392), .A2(new_n395), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT75), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n392), .A2(new_n395), .A3(new_n415), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n396), .A2(new_n410), .A3(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n412), .A2(new_n419), .A3(new_n421), .A4(new_n423), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n312), .A2(new_n350), .A3(new_n370), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT6), .ZN(new_n427));
  AND2_X1   g0227(.A1(G97), .A2(G107), .ZN(new_n428));
  NOR2_X1   g0228(.A1(G97), .A2(G107), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n362), .A2(KEYINPUT6), .A3(G97), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(G20), .B1(G77), .B2(new_n265), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n362), .B1(new_n386), .B2(new_n372), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(KEYINPUT76), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT76), .ZN(new_n436));
  AOI211_X1 g0236(.A(new_n436), .B(new_n362), .C1(new_n386), .C2(new_n372), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n255), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G97), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n253), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n251), .A2(G33), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n252), .A2(new_n441), .A3(new_n229), .A4(new_n254), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n442), .B2(new_n439), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n438), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT80), .ZN(new_n446));
  INV_X1    g0246(.A(G1698), .ZN(new_n447));
  OAI211_X1 g0247(.A(G244), .B(new_n447), .C1(new_n284), .C2(new_n285), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT4), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n293), .A2(KEYINPUT4), .A3(G244), .A4(new_n447), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n293), .A2(G250), .A3(G1698), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G283), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n297), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n251), .B(G45), .C1(new_n275), .C2(KEYINPUT5), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G41), .ZN(new_n458));
  OAI211_X1 g0258(.A(G257), .B(new_n280), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n274), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT77), .B1(new_n457), .B2(G41), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT77), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(new_n275), .A3(KEYINPUT5), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n457), .A2(G41), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n276), .A2(G1), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n461), .A2(new_n463), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n459), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT78), .ZN(new_n468));
  INV_X1    g0268(.A(new_n456), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(new_n274), .A3(new_n461), .A4(new_n463), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT78), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n459), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n455), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G169), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n455), .A2(new_n468), .A3(G179), .A4(new_n472), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n445), .A2(new_n446), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n438), .A2(KEYINPUT80), .A3(new_n444), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(KEYINPUT79), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT79), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n455), .A2(new_n468), .A3(new_n479), .A4(new_n472), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(G200), .A3(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n455), .A2(new_n468), .A3(G190), .A4(new_n472), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n438), .A2(new_n482), .A3(new_n444), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n476), .A2(new_n477), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(G244), .B(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n485));
  OAI211_X1 g0285(.A(G238), .B(new_n447), .C1(new_n284), .C2(new_n285), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G116), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n297), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n220), .B1(new_n276), .B2(G1), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n251), .A2(new_n271), .A3(G45), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n280), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(G169), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n488), .B2(new_n297), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n494), .B1(new_n309), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n354), .A2(new_n252), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n263), .A2(new_n498), .A3(G97), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G97), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n429), .A2(new_n219), .B1(new_n500), .B2(new_n228), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n501), .B2(new_n498), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n293), .A2(KEYINPUT81), .A3(new_n228), .A4(G68), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n228), .B(G68), .C1(new_n284), .C2(new_n285), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT81), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n497), .B1(new_n507), .B2(new_n255), .ZN(new_n508));
  INV_X1    g0308(.A(new_n354), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(new_n442), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n300), .B1(new_n489), .B2(new_n493), .ZN(new_n511));
  AOI211_X1 g0311(.A(new_n348), .B(new_n492), .C1(new_n488), .C2(new_n297), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n442), .A2(new_n219), .ZN(new_n514));
  AOI211_X1 g0314(.A(new_n497), .B(new_n514), .C1(new_n507), .C2(new_n255), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n496), .A2(new_n510), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n484), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(G270), .B(new_n280), .C1(new_n456), .C2(new_n458), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n460), .B2(new_n466), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G264), .B(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n521));
  OAI211_X1 g0321(.A(G257), .B(new_n447), .C1(new_n284), .C2(new_n285), .ZN(new_n522));
  INV_X1    g0322(.A(G303), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n293), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n297), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT85), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT82), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n256), .A2(new_n529), .A3(G116), .A4(new_n441), .ZN(new_n530));
  INV_X1    g0330(.A(G116), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT82), .B1(new_n442), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n262), .A2(G97), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT83), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n534), .A2(new_n535), .A3(new_n228), .A4(new_n453), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n254), .A2(new_n229), .B1(G20), .B2(new_n531), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n453), .B(new_n228), .C1(G33), .C2(new_n439), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT83), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(KEYINPUT20), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n536), .A3(new_n537), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT20), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n541), .A2(new_n544), .B1(new_n531), .B2(new_n253), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n527), .A2(new_n528), .A3(new_n533), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n253), .A2(new_n531), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT20), .B1(new_n538), .B2(new_n540), .ZN(new_n548));
  AND4_X1   g0348(.A1(KEYINPUT20), .A2(new_n540), .A3(new_n536), .A4(new_n537), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n533), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n300), .B1(new_n520), .B2(new_n525), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT85), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n520), .A2(new_n525), .A3(G190), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n546), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G169), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n520), .B2(new_n525), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n556), .A2(KEYINPUT21), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n520), .A2(new_n525), .A3(G179), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n550), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT84), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n550), .A2(new_n556), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT21), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI211_X1 g0364(.A(KEYINPUT84), .B(KEYINPUT21), .C1(new_n550), .C2(new_n556), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n554), .B(new_n560), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(G264), .B(new_n280), .C1(new_n456), .C2(new_n458), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n470), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G257), .B(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n570));
  OAI211_X1 g0370(.A(G250), .B(new_n447), .C1(new_n284), .C2(new_n285), .ZN(new_n571));
  INV_X1    g0371(.A(G294), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n571), .C1(new_n262), .C2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(KEYINPUT87), .A3(new_n297), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n297), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n555), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n576), .A2(G179), .A3(new_n470), .A4(new_n567), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT88), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n569), .A2(KEYINPUT88), .A3(G179), .A4(new_n576), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n228), .B(G87), .C1(new_n284), .C2(new_n285), .ZN(new_n585));
  XNOR2_X1  g0385(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT22), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(KEYINPUT86), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n293), .A2(new_n228), .A3(G87), .A4(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n487), .A2(G20), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT23), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n228), .B2(G107), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n362), .A2(KEYINPUT23), .A3(G20), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n587), .A2(new_n590), .A3(new_n595), .ZN(new_n596));
  OR2_X1    g0396(.A1(new_n596), .A2(KEYINPUT24), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(KEYINPUT24), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n260), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT25), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n252), .B2(G107), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n252), .A2(new_n600), .A3(G107), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n602), .A2(new_n603), .B1(new_n362), .B2(new_n442), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n579), .A2(new_n584), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n599), .A2(new_n604), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n578), .A2(new_n348), .A3(new_n569), .A4(new_n574), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n569), .A2(new_n576), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n300), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n566), .A2(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n426), .A2(new_n517), .A3(new_n613), .ZN(G372));
  INV_X1    g0414(.A(new_n311), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n403), .A2(new_n407), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n396), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT18), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n392), .A2(new_n395), .B1(new_n407), .B2(new_n403), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n422), .ZN(new_n620));
  INV_X1    g0420(.A(new_n345), .ZN(new_n621));
  INV_X1    g0421(.A(new_n368), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n349), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n419), .A2(new_n421), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n618), .B(new_n620), .C1(new_n623), .C2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n615), .B1(new_n626), .B2(new_n308), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT89), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(new_n629));
  INV_X1    g0429(.A(new_n579), .ZN(new_n630));
  INV_X1    g0430(.A(new_n584), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n606), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n265), .A2(G77), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n362), .A2(KEYINPUT6), .A3(G97), .ZN(new_n635));
  XNOR2_X1  g0435(.A(G97), .B(G107), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(new_n427), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n637), .B2(new_n228), .ZN(new_n638));
  OAI21_X1  g0438(.A(G107), .B1(new_n371), .B2(new_n373), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n436), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n437), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n260), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n446), .B1(new_n642), .B2(new_n443), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n474), .A2(new_n475), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n477), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n481), .A2(new_n483), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(new_n516), .A4(new_n611), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n628), .B1(new_n633), .B2(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n605), .B(new_n560), .C1(new_n564), .C2(new_n565), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n611), .A2(new_n516), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n484), .A3(new_n650), .A4(KEYINPUT89), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n496), .A2(new_n510), .ZN(new_n653));
  INV_X1    g0453(.A(new_n472), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n471), .B1(new_n470), .B2(new_n459), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n555), .B1(new_n656), .B2(new_n455), .ZN(new_n657));
  INV_X1    g0457(.A(new_n475), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT90), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT90), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n474), .A2(new_n660), .A3(new_n475), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n659), .A2(new_n445), .A3(new_n516), .A4(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT91), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT91), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(new_n666), .A3(new_n663), .ZN(new_n667));
  INV_X1    g0467(.A(new_n516), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n645), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n665), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n652), .A2(new_n653), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n627), .B1(new_n673), .B2(new_n426), .ZN(G369));
  NAND3_X1  g0474(.A1(new_n251), .A2(new_n228), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n545), .B2(new_n533), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n629), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT92), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n683), .B(KEYINPUT92), .C1(new_n566), .C2(new_n682), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n612), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n606), .B2(new_n681), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n605), .B2(new_n681), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(G330), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n629), .A2(new_n681), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n680), .B(KEYINPUT93), .Z(new_n692));
  AOI22_X1  g0492(.A1(new_n691), .A2(new_n687), .B1(new_n632), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n211), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n429), .A2(new_n219), .A3(new_n531), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n696), .A2(new_n251), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n227), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n696), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT28), .Z(new_n701));
  NAND2_X1  g0501(.A1(new_n662), .A2(KEYINPUT26), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n476), .A2(new_n663), .A3(new_n477), .A4(new_n516), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(new_n653), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n633), .A2(new_n647), .ZN(new_n705));
  OAI211_X1 g0505(.A(KEYINPUT29), .B(new_n681), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n692), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n664), .A2(KEYINPUT91), .B1(new_n669), .B2(KEYINPUT26), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n708), .A2(new_n667), .B1(new_n510), .B2(new_n496), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n707), .B1(new_n709), .B2(new_n652), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n706), .B1(new_n710), .B2(KEYINPUT29), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n495), .A2(new_n576), .A3(new_n567), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n473), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n712), .B1(new_n714), .B2(new_n559), .ZN(new_n715));
  NOR4_X1   g0515(.A1(new_n473), .A2(new_n558), .A3(new_n713), .A4(KEYINPUT30), .ZN(new_n716));
  INV_X1    g0516(.A(new_n473), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n495), .A2(G179), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(new_n608), .A3(new_n526), .ZN(new_n719));
  OAI22_X1  g0519(.A1(new_n715), .A2(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT95), .ZN(new_n721));
  XNOR2_X1  g0521(.A(KEYINPUT94), .B(KEYINPUT31), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n720), .A2(new_n721), .A3(new_n707), .A4(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n717), .A2(new_n719), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n495), .A2(new_n576), .A3(new_n567), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n559), .A2(new_n727), .A3(new_n656), .A4(new_n455), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT30), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n717), .A2(new_n712), .A3(new_n559), .A4(new_n727), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n725), .B1(new_n731), .B2(new_n681), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n707), .A2(new_n723), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT95), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n724), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n645), .A2(new_n646), .A3(new_n516), .A4(new_n692), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n736), .A2(new_n612), .A3(new_n566), .ZN(new_n737));
  OAI21_X1  g0537(.A(G330), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n711), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n701), .B1(new_n740), .B2(G1), .ZN(G364));
  NAND2_X1  g0541(.A1(new_n686), .A2(G330), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n209), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n251), .B1(new_n743), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n696), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n686), .A2(G330), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n686), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n695), .A2(new_n286), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n755), .A2(G355), .B1(new_n531), .B2(new_n695), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n695), .A2(new_n293), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G45), .B2(new_n227), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n249), .A2(new_n276), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n229), .B1(G20), .B2(new_n555), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n752), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n747), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  OR3_X1    g0563(.A1(new_n228), .A2(KEYINPUT96), .A3(G190), .ZN(new_n764));
  OAI21_X1  g0564(.A(KEYINPUT96), .B1(new_n228), .B2(G190), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G179), .A2(G200), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT97), .B(G159), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT32), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n228), .A2(new_n309), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n773), .A2(new_n348), .A3(G200), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G58), .A2(new_n774), .B1(new_n775), .B2(G77), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n348), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n777), .A2(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n776), .B1(new_n244), .B2(new_n779), .C1(new_n217), .C2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n228), .B1(new_n766), .B2(G190), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n771), .B(new_n782), .C1(G97), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n300), .A2(G179), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(G20), .A3(G190), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n764), .A2(new_n789), .A3(new_n765), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n293), .B1(new_n790), .B2(new_n219), .C1(new_n791), .C2(new_n362), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT98), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n775), .A2(G311), .B1(new_n778), .B2(G326), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n572), .B2(new_n786), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT100), .Z(new_n796));
  INV_X1    g0596(.A(new_n790), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n293), .B1(new_n797), .B2(G303), .ZN(new_n798));
  INV_X1    g0598(.A(G329), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n798), .A2(KEYINPUT101), .B1(new_n799), .B2(new_n767), .ZN(new_n800));
  INV_X1    g0600(.A(G317), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(KEYINPUT33), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(KEYINPUT33), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n780), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  INV_X1    g0605(.A(new_n774), .ZN(new_n806));
  INV_X1    g0606(.A(G322), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n804), .B1(new_n805), .B2(new_n791), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n800), .B(new_n808), .C1(KEYINPUT101), .C2(new_n798), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n788), .A2(new_n793), .B1(new_n796), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n761), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n763), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n748), .A2(new_n749), .B1(new_n754), .B2(new_n812), .ZN(G396));
  NOR2_X1   g0613(.A1(new_n368), .A2(new_n680), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n366), .B1(new_n357), .B2(new_n681), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(new_n815), .B2(new_n368), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n707), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n672), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n710), .B2(new_n816), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n746), .B1(new_n820), .B2(new_n738), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n738), .B2(new_n820), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n769), .A2(new_n775), .B1(new_n774), .B2(G143), .ZN(new_n823));
  INV_X1    g0623(.A(G150), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n781), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G137), .B2(new_n778), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT34), .Z(new_n827));
  OAI21_X1  g0627(.A(new_n293), .B1(new_n790), .B2(new_n244), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n791), .A2(new_n217), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(G132), .C2(new_n768), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n827), .B(new_n830), .C1(new_n375), .C2(new_n786), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n786), .A2(new_n439), .B1(new_n806), .B2(new_n572), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT102), .Z(new_n833));
  INV_X1    g0633(.A(new_n775), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n286), .B1(new_n362), .B2(new_n790), .C1(new_n834), .C2(new_n531), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n781), .A2(new_n805), .B1(new_n779), .B2(new_n523), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n791), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(G87), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n837), .B(new_n839), .C1(new_n840), .C2(new_n767), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n831), .B1(new_n833), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n761), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n761), .A2(new_n750), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n747), .B1(new_n289), .B2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n843), .B(new_n845), .C1(new_n816), .C2(new_n751), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n822), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  NAND3_X1  g0648(.A1(new_n345), .A2(new_n349), .A3(KEYINPUT104), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n324), .A2(new_n680), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT104), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n345), .A2(new_n349), .A3(new_n852), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n850), .A2(new_n343), .A3(new_n344), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n722), .B1(new_n731), .B2(new_n681), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(new_n613), .C2(new_n736), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n856), .A2(new_n816), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT40), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT37), .B1(new_n396), .B2(new_n410), .ZN(new_n863));
  INV_X1    g0663(.A(new_n678), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n396), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n416), .A3(new_n865), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n392), .A2(new_n395), .A3(new_n415), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n678), .B1(new_n392), .B2(new_n395), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n867), .A2(new_n619), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT106), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n618), .A2(new_n419), .A3(new_n421), .A4(new_n620), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n871), .A2(new_n872), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n617), .A2(new_n865), .A3(new_n416), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT37), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(KEYINPUT106), .A3(new_n866), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n424), .A2(new_n868), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n871), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n878), .A2(KEYINPUT108), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT108), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n873), .A2(new_n868), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n867), .A2(new_n868), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n875), .A2(KEYINPUT37), .B1(new_n886), .B2(new_n863), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(KEYINPUT106), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n877), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n883), .B1(new_n890), .B2(new_n880), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n862), .B1(new_n882), .B2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n396), .A2(new_n410), .A3(new_n422), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n422), .B1(new_n396), .B2(new_n410), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n865), .B1(new_n895), .B2(new_n624), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n884), .B1(new_n896), .B2(new_n887), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n880), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n861), .B1(new_n860), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n892), .A2(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n425), .A2(new_n859), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(G330), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT107), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n880), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n906), .B1(new_n878), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n880), .A2(new_n907), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n890), .A2(new_n910), .A3(KEYINPUT107), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT105), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n898), .B2(KEYINPUT39), .ZN(new_n913));
  AOI211_X1 g0713(.A(KEYINPUT105), .B(new_n907), .C1(new_n897), .C2(new_n880), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n909), .B(new_n911), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n621), .A2(new_n681), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n864), .B1(new_n618), .B2(new_n620), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n851), .A2(new_n855), .ZN(new_n920));
  INV_X1    g0720(.A(new_n814), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n819), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n919), .B1(new_n922), .B2(new_n898), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n425), .B(new_n706), .C1(new_n710), .C2(KEYINPUT29), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n627), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n924), .B(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n905), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n928), .A2(KEYINPUT109), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(KEYINPUT109), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n905), .A2(new_n927), .B1(new_n251), .B2(new_n743), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n432), .A2(KEYINPUT35), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n432), .A2(KEYINPUT35), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n229), .A2(new_n228), .A3(new_n531), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT36), .Z(new_n937));
  OR3_X1    g0737(.A1(new_n227), .A2(new_n289), .A3(new_n376), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n245), .B(KEYINPUT103), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n251), .B(G13), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  OR3_X1    g0740(.A1(new_n932), .A2(new_n937), .A3(new_n940), .ZN(G367));
  NAND2_X1  g0741(.A1(new_n757), .A2(new_n239), .ZN(new_n942));
  INV_X1    g0742(.A(new_n762), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n695), .B2(new_n354), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n747), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n515), .A2(new_n681), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n516), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n653), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n791), .A2(new_n439), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n286), .B1(new_n806), .B2(new_n523), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n949), .B(new_n950), .C1(G283), .C2(new_n775), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT46), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n790), .A2(new_n952), .A3(new_n531), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n790), .B2(new_n531), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n781), .B2(new_n572), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n953), .B(new_n955), .C1(G311), .C2(new_n778), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n768), .A2(G317), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n787), .A2(G107), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n951), .A2(new_n956), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n787), .A2(G68), .ZN(new_n960));
  INV_X1    g0760(.A(G143), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n960), .B1(new_n961), .B2(new_n779), .C1(new_n824), .C2(new_n806), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT110), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT111), .B(G137), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n289), .A2(new_n791), .B1(new_n767), .B2(new_n964), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n293), .B1(new_n375), .B2(new_n790), .C1(new_n834), .C2(new_n244), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n965), .B(new_n966), .C1(new_n769), .C2(new_n780), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n962), .A2(KEYINPUT110), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n959), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT47), .Z(new_n971));
  OAI221_X1 g0771(.A(new_n945), .B1(new_n753), .B2(new_n948), .C1(new_n971), .C2(new_n811), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT112), .Z(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n707), .A2(new_n445), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n484), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n659), .A2(new_n445), .A3(new_n661), .A4(new_n707), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n693), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT45), .Z(new_n980));
  NOR2_X1   g0780(.A1(new_n693), .A2(new_n978), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(new_n690), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n691), .A2(new_n687), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n689), .B2(new_n691), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n742), .B(new_n986), .Z(new_n987));
  NAND2_X1  g0787(.A1(new_n740), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n740), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n696), .B(KEYINPUT41), .Z(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n745), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n978), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n985), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT42), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n645), .B1(new_n993), .B2(new_n605), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n692), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n995), .A2(new_n997), .B1(KEYINPUT43), .B2(new_n948), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n690), .A2(new_n993), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n974), .B1(new_n992), .B2(new_n1002), .ZN(G387));
  NAND2_X1  g0803(.A1(new_n987), .A2(new_n745), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT113), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n689), .A2(new_n753), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n261), .A2(new_n244), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT50), .Z(new_n1008));
  AOI211_X1 g0808(.A(G45), .B(new_n697), .C1(G68), .C2(G77), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n757), .B(new_n1010), .C1(new_n236), .C2(new_n276), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n755), .A2(new_n697), .B1(new_n362), .B2(new_n695), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1011), .A2(KEYINPUT114), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n762), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT114), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n746), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n293), .B1(new_n806), .B2(new_n244), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n834), .A2(new_n217), .B1(new_n289), .B2(new_n790), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n261), .C2(new_n780), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n949), .B1(G150), .B2(new_n768), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n778), .A2(G159), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT115), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n787), .A2(new_n354), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n781), .A2(new_n840), .B1(new_n779), .B2(new_n807), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(KEYINPUT116), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(KEYINPUT116), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G303), .A2(new_n775), .B1(new_n774), .B2(G317), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n786), .A2(new_n805), .B1(new_n572), .B2(new_n790), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n293), .B1(new_n768), .B2(G326), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n531), .C2(new_n791), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT49), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1024), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1016), .B1(new_n1038), .B2(new_n761), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1005), .B1(new_n1006), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n740), .A2(new_n987), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n988), .A2(new_n696), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(G393));
  AOI22_X1  g0843(.A1(new_n774), .A2(G159), .B1(new_n778), .B2(G150), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT117), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n839), .B1(new_n961), .B2(new_n767), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n293), .B1(new_n217), .B2(new_n790), .C1(new_n834), .C2(new_n394), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G50), .C2(new_n780), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n787), .A2(G77), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n774), .A2(G311), .B1(new_n778), .B2(G317), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT52), .Z(new_n1054));
  OAI221_X1 g0854(.A(new_n286), .B1(new_n805), .B2(new_n790), .C1(new_n834), .C2(new_n572), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G303), .B2(new_n780), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n787), .A2(G116), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G107), .A2(new_n838), .B1(new_n768), .B2(G322), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1054), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n811), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n243), .A2(new_n757), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n943), .B1(new_n695), .B2(G97), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n747), .B(new_n1060), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT118), .Z(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n753), .B2(new_n978), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n984), .A2(new_n988), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n696), .B1(new_n984), .B2(new_n988), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1065), .B1(new_n744), .B2(new_n984), .C1(new_n1067), .C2(new_n1068), .ZN(G390));
  INV_X1    g0869(.A(new_n696), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n815), .A2(new_n368), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n681), .B(new_n1071), .C1(new_n704), .C2(new_n705), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n921), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n917), .B1(new_n856), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n882), .B2(new_n891), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n819), .A2(new_n921), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n917), .B1(new_n1076), .B2(new_n856), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n915), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n851), .A2(new_n855), .A3(new_n816), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n857), .A2(new_n858), .ZN(new_n1080));
  OAI21_X1  g0880(.A(G330), .B1(new_n737), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT119), .ZN(new_n1084));
  OAI211_X1 g0884(.A(G330), .B(new_n816), .C1(new_n735), .C2(new_n737), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1075), .B1(new_n920), .B2(new_n1085), .C1(new_n915), .C2(new_n1077), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT119), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1078), .A2(new_n1087), .A3(new_n1082), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1085), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n856), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1076), .B1(new_n1091), .B2(new_n1082), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT120), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1093), .B(G330), .C1(new_n737), .C2(new_n1080), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n816), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1093), .B1(new_n859), .B2(G330), .ZN(new_n1096));
  OAI211_X1 g0896(.A(KEYINPUT121), .B(new_n920), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1073), .B1(new_n856), .B2(new_n1090), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1081), .A2(KEYINPUT120), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(new_n816), .A3(new_n1094), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT121), .B1(new_n1101), .B2(new_n920), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1092), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n425), .A2(G330), .A3(new_n859), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n925), .A2(new_n627), .A3(new_n1104), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1103), .A2(KEYINPUT122), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT122), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1070), .B1(new_n1089), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1088), .A2(new_n1086), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1087), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT122), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1103), .A2(new_n1105), .A3(KEYINPUT122), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT123), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT123), .ZN(new_n1119));
  NOR4_X1   g0919(.A1(new_n1108), .A2(new_n1110), .A3(new_n1119), .A4(new_n1111), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1109), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n844), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n293), .B1(new_n797), .B2(G87), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n779), .B2(new_n805), .C1(new_n531), .C2(new_n806), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n829), .B(new_n1124), .C1(G294), .C2(new_n768), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G97), .A2(new_n775), .B1(new_n780), .B2(G107), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1051), .B1(new_n1127), .B2(KEYINPUT124), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(KEYINPUT124), .B2(new_n1127), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n791), .A2(new_n244), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n797), .A2(G150), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1130), .B(new_n1132), .C1(G125), .C2(new_n768), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1134), .A2(new_n779), .B1(new_n781), .B2(new_n964), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n774), .A2(G132), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(new_n293), .C1(new_n834), .C2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1135), .B(new_n1138), .C1(G159), .C2(new_n787), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1125), .A2(new_n1129), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n746), .B1(new_n261), .B2(new_n1122), .C1(new_n1140), .C2(new_n811), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n915), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n750), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1112), .B2(new_n745), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1121), .A2(new_n1144), .ZN(G378));
  NAND3_X1  g0945(.A1(new_n892), .A2(G330), .A3(new_n900), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n312), .A2(new_n269), .A3(new_n864), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n269), .A2(new_n864), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n308), .A2(new_n311), .A3(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1147), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1146), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1146), .A2(new_n1153), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n924), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1146), .A2(new_n1153), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n924), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n1154), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n744), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1153), .A2(new_n750), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n746), .B1(G50), .B2(new_n1122), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(G33), .A2(G41), .ZN(new_n1164));
  AOI211_X1 g0964(.A(G50), .B(new_n1164), .C1(new_n286), .C2(new_n275), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n362), .A2(new_n806), .B1(new_n834), .B2(new_n509), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n781), .A2(new_n439), .B1(new_n779), .B2(new_n531), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n275), .B(new_n286), .C1(new_n790), .C2(new_n289), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G58), .A2(new_n838), .B1(new_n768), .B2(G283), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n960), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT58), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1165), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n787), .A2(G150), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n775), .A2(G137), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1137), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n774), .A2(G128), .B1(new_n797), .B2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G125), .A2(new_n778), .B1(new_n780), .B2(G132), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1174), .A2(new_n1175), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n768), .A2(G124), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n838), .A2(new_n769), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1164), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1173), .B1(new_n1172), .B2(new_n1171), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1163), .B1(new_n1185), .B2(new_n761), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1162), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT125), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1161), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1105), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT57), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1105), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1119), .B1(new_n1089), .B2(new_n1108), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1110), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1195), .A2(new_n1117), .A3(KEYINPUT123), .A4(new_n1084), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1193), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1191), .A2(KEYINPUT57), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n696), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1189), .B1(new_n1192), .B2(new_n1199), .ZN(G375));
  OR2_X1    g1000(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1115), .A2(new_n1116), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n991), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n806), .A2(new_n805), .B1(new_n439), .B2(new_n790), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n293), .B(new_n1204), .C1(G107), .C2(new_n775), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G116), .A2(new_n780), .B1(new_n778), .B2(G294), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G77), .A2(new_n838), .B1(new_n768), .B2(G303), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1205), .A2(new_n1023), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n806), .A2(new_n964), .B1(new_n389), .B2(new_n790), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n286), .B(new_n1209), .C1(G150), .C2(new_n775), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n787), .A2(G50), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G132), .A2(new_n778), .B1(new_n780), .B2(new_n1176), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G58), .A2(new_n838), .B1(new_n768), .B2(G128), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1208), .A2(new_n1214), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n746), .B1(G68), .B2(new_n1122), .C1(new_n1215), .C2(new_n811), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n920), .B2(new_n750), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1103), .B2(new_n745), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1203), .A2(new_n1218), .ZN(G381));
  NOR4_X1   g1019(.A1(G390), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1220));
  INV_X1    g1020(.A(G387), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OR4_X1    g1022(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1222), .ZN(G407));
  NAND2_X1  g1023(.A1(new_n679), .A2(G213), .ZN(new_n1224));
  OR3_X1    g1024(.A1(G375), .A2(G378), .A3(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(G407), .A2(G213), .A3(new_n1225), .ZN(G409));
  OR2_X1    g1026(.A1(new_n1221), .A2(G390), .ZN(new_n1227));
  XOR2_X1   g1027(.A(G393), .B(G396), .Z(new_n1228));
  NAND2_X1  g1028(.A1(new_n1221), .A2(G390), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1228), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G378), .B(new_n1189), .C1(new_n1192), .C2(new_n1199), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1121), .A2(new_n1144), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1155), .A2(new_n1156), .A3(new_n924), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1159), .B1(new_n1158), .B2(new_n1154), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(KEYINPUT126), .B(new_n1187), .C1(new_n1238), .C2(new_n744), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT126), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1187), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1240), .B1(new_n1161), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1197), .A2(new_n990), .A3(new_n1238), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1235), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1234), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1224), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1070), .B1(new_n1201), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n1202), .B2(new_n1248), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1218), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(G384), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n679), .A2(G213), .A3(G2897), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1252), .B(new_n1253), .Z(new_n1254));
  NAND2_X1  g1054(.A1(new_n1247), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT127), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1246), .A2(new_n1224), .A3(new_n1252), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT62), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1234), .A2(new_n1245), .B1(G213), .B2(new_n679), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT62), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1261), .A3(new_n1252), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1233), .B1(new_n1257), .B2(new_n1263), .ZN(new_n1264));
  AND4_X1   g1064(.A1(KEYINPUT63), .A2(new_n1246), .A3(new_n1224), .A4(new_n1252), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT63), .B1(new_n1260), .B2(new_n1252), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1232), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT127), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1252), .B(new_n1253), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1269), .B(new_n1256), .C1(new_n1260), .C2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1264), .A2(new_n1273), .ZN(G405));
  NAND2_X1  g1074(.A1(G375), .A2(new_n1235), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1234), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1276), .A2(new_n1252), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1252), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1233), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1277), .A2(new_n1232), .A3(new_n1278), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(G402));
endmodule


