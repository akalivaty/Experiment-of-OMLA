//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT67), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(new_n202), .A3(G113gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G113gat), .B(G120gat), .ZN(new_n212));
  INV_X1    g011(.A(G127gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G134gat), .ZN(new_n214));
  INV_X1    g013(.A(G134gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G127gat), .ZN(new_n216));
  OAI22_X1  g015(.A1(new_n212), .A2(KEYINPUT1), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G155gat), .B(G162gat), .ZN(new_n219));
  INV_X1    g018(.A(G141gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G148gat), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G141gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n221), .A2(new_n223), .B1(KEYINPUT2), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n219), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(KEYINPUT2), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n222), .A2(G141gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n220), .A2(G148gat), .ZN(new_n230));
  OAI211_X1 g029(.A(KEYINPUT79), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT78), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT79), .ZN(new_n235));
  OAI211_X1 g034(.A(KEYINPUT78), .B(new_n219), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n218), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n226), .B1(new_n225), .B2(KEYINPUT79), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n226), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n239));
  XOR2_X1   g038(.A(G155gat), .B(G162gat), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n236), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n211), .A2(KEYINPUT80), .A3(new_n217), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT80), .B1(new_n211), .B2(new_n217), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n237), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT5), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(new_n242), .B2(new_n243), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n233), .A2(KEYINPUT3), .A3(new_n236), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n247), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n236), .ZN(new_n255));
  INV_X1    g054(.A(new_n218), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n237), .A2(KEYINPUT4), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n254), .A2(new_n259), .A3(new_n249), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n250), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n237), .B(new_n258), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n263), .A2(KEYINPUT5), .A3(new_n249), .A4(new_n254), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G1gat), .B(G29gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT0), .ZN(new_n267));
  XNOR2_X1  g066(.A(G57gat), .B(G85gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(KEYINPUT82), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n269), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n262), .A2(new_n273), .A3(new_n264), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT82), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n262), .B2(new_n264), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(KEYINPUT6), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT6), .A4(new_n273), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G8gat), .B(G36gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT77), .ZN(new_n282));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G226gat), .A2(G233gat), .ZN(new_n285));
  INV_X1    g084(.A(G183gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT64), .B1(new_n286), .B2(KEYINPUT27), .ZN(new_n287));
  OR2_X1    g086(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT65), .B1(new_n286), .B2(KEYINPUT27), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(G183gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n286), .A2(KEYINPUT64), .A3(KEYINPUT27), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n289), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(G183gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n286), .A2(KEYINPUT27), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n297), .B1(new_n301), .B2(KEYINPUT28), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n304));
  AND2_X1   g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n307), .A2(KEYINPUT66), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(KEYINPUT66), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(KEYINPUT24), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  INV_X1    g114(.A(G169gat), .ZN(new_n316));
  INV_X1    g115(.A(G176gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n286), .A2(new_n300), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(KEYINPUT24), .A3(new_n312), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n314), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n314), .A2(new_n320), .A3(new_n322), .A4(KEYINPUT25), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n303), .A2(new_n310), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n285), .B1(new_n327), .B2(KEYINPUT29), .ZN(new_n328));
  NAND2_X1  g127(.A1(G211gat), .A2(G218gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT22), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT73), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n329), .A2(new_n333), .A3(new_n330), .ZN(new_n334));
  XNOR2_X1  g133(.A(G197gat), .B(G204gat), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(G211gat), .A2(G218gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n329), .ZN(new_n340));
  INV_X1    g139(.A(new_n329), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT75), .B1(new_n341), .B2(new_n337), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n342), .A3(KEYINPUT74), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n345), .A2(KEYINPUT74), .A3(new_n342), .A4(new_n340), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n310), .A2(new_n296), .A3(new_n302), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n313), .B1(new_n319), .B2(new_n318), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT25), .B1(new_n350), .B2(new_n322), .ZN(new_n351));
  INV_X1    g150(.A(new_n326), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n285), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n348), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n325), .A2(new_n326), .ZN(new_n356));
  AOI211_X1 g155(.A(KEYINPUT76), .B(new_n285), .C1(new_n356), .C2(new_n349), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n328), .B(new_n347), .C1(new_n355), .C2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n347), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n327), .A2(new_n285), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n354), .B1(new_n353), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n284), .B1(new_n358), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n358), .A2(new_n363), .A3(new_n284), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n358), .A2(new_n363), .ZN(new_n370));
  INV_X1    g169(.A(new_n284), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n370), .A2(KEYINPUT30), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT83), .B1(new_n280), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n218), .A2(KEYINPUT68), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n218), .A2(KEYINPUT68), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n353), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AND2_X1   g179(.A1(G227gat), .A2(G233gat), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n356), .A2(KEYINPUT68), .A3(new_n218), .A4(new_n349), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT69), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n380), .A2(KEYINPUT69), .A3(new_n381), .A4(new_n382), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n377), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT33), .B1(new_n385), .B2(new_n386), .ZN(new_n388));
  XOR2_X1   g187(.A(G15gat), .B(G43gat), .Z(new_n389));
  XNOR2_X1  g188(.A(G71gat), .B(G99gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n387), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  AOI221_X4 g192(.A(new_n377), .B1(KEYINPUT33), .B2(new_n391), .C1(new_n385), .C2(new_n386), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT70), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n381), .B1(new_n380), .B2(new_n382), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT34), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n396), .A2(new_n397), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n392), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n387), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT70), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n387), .B1(new_n388), .B2(new_n392), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n395), .A2(new_n401), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n400), .A3(new_n408), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT29), .B1(new_n344), .B2(new_n346), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n244), .B1(new_n412), .B2(KEYINPUT3), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G228gat), .ZN(new_n416));
  INV_X1    g215(.A(G233gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n251), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n419), .B1(new_n233), .B2(new_n236), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n359), .B1(new_n420), .B2(KEYINPUT29), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n244), .B(KEYINPUT84), .C1(new_n412), .C2(KEYINPUT3), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n415), .A2(new_n418), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n347), .B1(new_n252), .B2(new_n361), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n336), .A2(new_n342), .A3(new_n340), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n340), .A2(new_n342), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n345), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n361), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n255), .B1(new_n428), .B2(new_n251), .ZN(new_n429));
  OAI22_X1  g228(.A1(new_n424), .A2(new_n429), .B1(new_n416), .B2(new_n417), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n423), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(G22gat), .ZN(new_n432));
  INV_X1    g231(.A(G22gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n423), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G78gat), .B(G106gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT31), .B(G50gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n423), .B2(new_n430), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n432), .A2(new_n440), .A3(new_n434), .A4(new_n438), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n411), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT89), .B1(new_n410), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n280), .A2(KEYINPUT83), .A3(new_n374), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n411), .A2(new_n442), .A3(new_n443), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT89), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n395), .A2(new_n401), .A3(new_n409), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n376), .A2(new_n445), .A3(new_n446), .A4(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n442), .A2(new_n443), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT35), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n279), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n270), .A2(new_n271), .A3(new_n274), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n279), .A2(new_n454), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n452), .A2(new_n453), .A3(new_n458), .A4(new_n374), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n411), .A2(KEYINPUT72), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n401), .B1(new_n393), .B2(new_n394), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT72), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n406), .A2(new_n462), .A3(new_n400), .A4(new_n408), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT88), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n367), .A2(new_n364), .A3(new_n365), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(new_n372), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(KEYINPUT35), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n452), .A2(new_n468), .A3(new_n458), .ZN(new_n469));
  INV_X1    g268(.A(new_n464), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n451), .A2(KEYINPUT35), .B1(new_n465), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT71), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n411), .A2(KEYINPUT36), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n474), .B1(new_n410), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT36), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n464), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n449), .A2(KEYINPUT71), .A3(KEYINPUT36), .A4(new_n411), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n442), .A2(new_n443), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT83), .ZN(new_n482));
  AOI211_X1 g281(.A(new_n482), .B(new_n467), .C1(new_n278), .C2(new_n279), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n375), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n274), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n263), .A2(new_n254), .ZN(new_n486));
  INV_X1    g285(.A(new_n249), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n269), .B1(new_n488), .B2(KEYINPUT39), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n248), .B2(new_n249), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n489), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT40), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT86), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n485), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(new_n467), .C1(new_n494), .C2(new_n492), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n370), .A2(KEYINPUT37), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n371), .B1(new_n370), .B2(KEYINPUT37), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT38), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n328), .B(new_n359), .C1(new_n355), .C2(new_n357), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n347), .B1(new_n360), .B2(new_n362), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(KEYINPUT37), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT38), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n499), .B(new_n368), .C1(new_n498), .C2(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n496), .B(new_n452), .C1(new_n458), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n480), .A2(new_n484), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n473), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G120gat), .B(G148gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(G176gat), .B(G204gat), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n510), .B(new_n511), .Z(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G71gat), .B(G78gat), .ZN(new_n514));
  XOR2_X1   g313(.A(G57gat), .B(G64gat), .Z(new_n515));
  INV_X1    g314(.A(KEYINPUT9), .ZN(new_n516));
  INV_X1    g315(.A(G71gat), .ZN(new_n517));
  INV_X1    g316(.A(G78gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n514), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n515), .A2(new_n514), .A3(new_n519), .ZN(new_n522));
  NAND2_X1  g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  OR2_X1    g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(KEYINPUT8), .B2(new_n526), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT98), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  AND4_X1   g331(.A1(new_n521), .A2(new_n522), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n524), .A2(new_n529), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n526), .A3(new_n525), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT97), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n530), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT94), .B1(new_n521), .B2(new_n522), .ZN(new_n539));
  INV_X1    g338(.A(new_n522), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n540), .A2(new_n541), .A3(new_n520), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n541), .B1(new_n540), .B2(new_n520), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n521), .A2(KEYINPUT94), .A3(new_n522), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n537), .B1(new_n547), .B2(new_n538), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n536), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT99), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT99), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n549), .A2(new_n554), .A3(new_n551), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT10), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n557), .B(new_n536), .C1(new_n544), .C2(new_n548), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n539), .A2(new_n542), .ZN(new_n559));
  INV_X1    g358(.A(new_n538), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(KEYINPUT10), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n551), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n513), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n558), .A2(new_n561), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n550), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n565), .A2(new_n553), .A3(new_n512), .A4(new_n555), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n559), .A2(KEYINPUT21), .ZN(new_n569));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G15gat), .B(G22gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT16), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(G1gat), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(G1gat), .B2(new_n572), .ZN(new_n575));
  INV_X1    g374(.A(G8gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n578), .B1(new_n559), .B2(KEYINPUT21), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n571), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT95), .ZN(new_n583));
  XOR2_X1   g382(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n581), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT96), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT14), .ZN(new_n591));
  INV_X1    g390(.A(G29gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n594));
  AOI21_X1  g393(.A(G36gat), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n592), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n596));
  OR3_X1    g395(.A1(new_n595), .A2(KEYINPUT15), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT15), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  XNOR2_X1  g397(.A(G43gat), .B(G50gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT91), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT17), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT91), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT17), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n607), .A2(new_n608), .A3(new_n538), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n603), .A2(new_n606), .A3(new_n560), .ZN(new_n610));
  INV_X1    g409(.A(G232gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(new_n417), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n590), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n607), .A2(new_n608), .A3(new_n538), .ZN(new_n616));
  INV_X1    g415(.A(new_n590), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n616), .A2(new_n617), .A3(new_n610), .A4(new_n613), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n620));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n615), .A2(new_n622), .A3(new_n618), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n568), .A2(new_n588), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n607), .A2(new_n577), .A3(new_n608), .ZN(new_n628));
  NAND2_X1  g427(.A1(G229gat), .A2(G233gat), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n603), .A2(new_n578), .A3(new_n606), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT92), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n628), .A2(KEYINPUT92), .A3(new_n629), .A4(new_n630), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n628), .A2(KEYINPUT18), .A3(new_n629), .A4(new_n630), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n603), .A2(new_n606), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n577), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n630), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n629), .B(KEYINPUT13), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G113gat), .B(G141gat), .Z(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G169gat), .B(G197gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT12), .Z(new_n649));
  AND3_X1   g448(.A1(new_n636), .A2(new_n643), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n636), .B2(new_n643), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n627), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n509), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n280), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g456(.A(new_n576), .B1(new_n654), .B2(new_n467), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT16), .B(G8gat), .ZN(new_n659));
  NOR4_X1   g458(.A1(new_n509), .A2(new_n374), .A3(new_n653), .A4(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT42), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(KEYINPUT42), .B2(new_n660), .ZN(G1325gat));
  AOI21_X1  g461(.A(G15gat), .B1(new_n654), .B2(new_n470), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT100), .Z(new_n664));
  INV_X1    g463(.A(new_n480), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n665), .A2(G15gat), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n654), .B2(new_n666), .ZN(G1326gat));
  NAND2_X1  g466(.A1(new_n654), .A2(new_n481), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT43), .B(G22gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  AND3_X1   g469(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n448), .B1(new_n447), .B2(new_n449), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n375), .A2(new_n483), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n453), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n472), .A2(new_n465), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n507), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n626), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n652), .A2(new_n588), .A3(new_n567), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(G29gat), .A3(new_n280), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n615), .A2(new_n622), .A3(new_n618), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n622), .B1(new_n615), .B2(new_n618), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n624), .A2(KEYINPUT103), .A3(new_n625), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n507), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n480), .A2(new_n484), .A3(KEYINPUT102), .A4(new_n506), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n473), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n691), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n677), .B2(new_n678), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n679), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n700), .A2(new_n280), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n683), .B1(new_n702), .B2(new_n592), .ZN(G1328gat));
  NOR3_X1   g502(.A1(new_n680), .A2(G36gat), .A3(new_n374), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT46), .ZN(new_n705));
  OAI21_X1  g504(.A(G36gat), .B1(new_n700), .B2(new_n374), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1329gat));
  OAI211_X1 g506(.A(new_n665), .B(new_n679), .C1(new_n697), .C2(new_n699), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G43gat), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n464), .A2(G43gat), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n677), .A2(new_n678), .A3(new_n679), .A4(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT47), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717));
  AOI211_X1 g516(.A(KEYINPUT104), .B(new_n717), .C1(new_n709), .C2(new_n713), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n716), .A2(new_n718), .ZN(G1330gat));
  OR2_X1    g518(.A1(new_n452), .A2(G50gat), .ZN(new_n720));
  OAI22_X1  g519(.A1(new_n680), .A2(new_n720), .B1(KEYINPUT106), .B2(KEYINPUT48), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n481), .B(new_n679), .C1(new_n697), .C2(new_n699), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(G50gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n723), .B(new_n724), .Z(G1331gat));
  AOI21_X1  g524(.A(new_n473), .B1(new_n693), .B2(new_n694), .ZN(new_n726));
  INV_X1    g525(.A(new_n652), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n588), .A2(new_n626), .A3(new_n567), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n655), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n467), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT49), .B(G64gat), .Z(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(G1333gat));
  NAND3_X1  g534(.A1(new_n729), .A2(new_n517), .A3(new_n470), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n729), .A2(new_n665), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(new_n517), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1334gat));
  NAND2_X1  g539(.A1(new_n729), .A2(new_n481), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g541(.A1(new_n727), .A2(new_n588), .A3(new_n568), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n697), .B2(new_n699), .ZN(new_n744));
  OAI21_X1  g543(.A(G85gat), .B1(new_n744), .B2(new_n280), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n695), .A2(new_n696), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n727), .A2(new_n588), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n678), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(KEYINPUT51), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n726), .B2(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(G85gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n655), .A2(new_n755), .A3(new_n567), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n745), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT107), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n745), .B(new_n759), .C1(new_n754), .C2(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1336gat));
  OAI211_X1 g560(.A(new_n467), .B(new_n743), .C1(new_n697), .C2(new_n699), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G92gat), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n568), .A2(G92gat), .A3(new_n374), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT108), .Z(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n750), .B2(new_n752), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n763), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n767), .A2(new_n764), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT52), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n765), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n763), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(G1337gat));
  INV_X1    g573(.A(G99gat), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n753), .A2(new_n775), .A3(new_n470), .A4(new_n567), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n744), .A2(new_n480), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n778), .B2(new_n775), .ZN(G1338gat));
  OAI21_X1  g578(.A(G106gat), .B1(new_n744), .B2(new_n452), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n568), .A2(new_n452), .A3(G106gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n753), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(G1339gat));
  NOR2_X1   g584(.A1(new_n280), .A2(new_n467), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n470), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n627), .A2(new_n727), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n636), .A2(new_n643), .A3(new_n649), .ZN(new_n789));
  INV_X1    g588(.A(new_n648), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n640), .A2(new_n641), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n629), .B1(new_n628), .B2(new_n630), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n567), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n558), .A2(new_n551), .A3(new_n561), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n565), .A2(KEYINPUT54), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n513), .B1(new_n565), .B2(KEYINPUT54), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n565), .A2(KEYINPUT54), .A3(new_n796), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n512), .B1(new_n562), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(new_n566), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n794), .B1(new_n804), .B2(new_n652), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n689), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n793), .ZN(new_n807));
  OR3_X1    g606(.A1(new_n804), .A2(new_n689), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n588), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n788), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT112), .B1(new_n811), .B2(new_n481), .ZN(new_n812));
  INV_X1    g611(.A(new_n788), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n804), .A2(new_n689), .A3(new_n807), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n689), .B2(new_n805), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n815), .B2(new_n588), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n817), .A3(new_n452), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n787), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n204), .B1(new_n819), .B2(new_n727), .ZN(new_n820));
  INV_X1    g619(.A(new_n673), .ZN(new_n821));
  INV_X1    g620(.A(new_n786), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n811), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n652), .A2(G113gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n820), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT114), .ZN(G1340gat));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n202), .A3(new_n567), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n202), .B1(new_n819), .B2(new_n567), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(G1341gat));
  NAND3_X1  g633(.A1(new_n823), .A2(new_n213), .A3(new_n588), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n819), .A2(new_n588), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n213), .ZN(G1342gat));
  NAND3_X1  g636(.A1(new_n823), .A2(new_n215), .A3(new_n678), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT116), .Z(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n838), .B(KEYINPUT116), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n819), .A2(new_n678), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n840), .B(new_n843), .C1(new_n215), .C2(new_n844), .ZN(G1343gat));
  NOR2_X1   g644(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n665), .A2(new_n822), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n452), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n797), .B2(new_n798), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n566), .A3(new_n803), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n794), .B1(new_n854), .B2(new_n652), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n626), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n814), .B1(new_n856), .B2(KEYINPUT118), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n855), .A2(new_n858), .A3(new_n626), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n588), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n849), .B(new_n851), .C1(new_n860), .C2(new_n788), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n850), .B1(new_n811), .B2(new_n452), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n855), .A2(new_n858), .A3(new_n626), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n858), .B1(new_n855), .B2(new_n626), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n864), .A2(new_n865), .A3(new_n814), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n813), .B1(new_n866), .B2(new_n588), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n849), .B1(new_n867), .B2(new_n851), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n727), .B(new_n848), .C1(new_n863), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G141gat), .ZN(new_n870));
  NAND2_X1  g669(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n811), .A2(new_n452), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n848), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n652), .A2(G141gat), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n871), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n847), .B1(new_n870), .B2(new_n877), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n846), .B(new_n876), .C1(new_n869), .C2(G141gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(G1344gat));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n848), .B1(new_n863), .B2(new_n868), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n881), .B(G148gat), .C1(new_n882), .C2(new_n568), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n816), .A2(new_n851), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n804), .A2(new_n626), .A3(new_n807), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n626), .B2(new_n855), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n813), .B1(new_n886), .B2(new_n588), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n481), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n568), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n222), .B1(new_n890), .B2(new_n848), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n883), .B1(new_n881), .B2(new_n891), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n872), .A2(new_n222), .A3(new_n567), .A4(new_n848), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1345gat));
  INV_X1    g693(.A(new_n882), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n588), .A2(G155gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n873), .A2(new_n810), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(KEYINPUT121), .ZN(new_n898));
  AOI21_X1  g697(.A(G155gat), .B1(new_n897), .B2(KEYINPUT121), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n895), .A2(new_n896), .B1(new_n898), .B2(new_n899), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n882), .B2(new_n689), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n626), .A2(G162gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n873), .B2(new_n902), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n655), .A2(new_n374), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n673), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n811), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n727), .ZN(new_n907));
  INV_X1    g706(.A(new_n904), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(new_n464), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n812), .B2(new_n818), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n652), .A2(new_n316), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(G1348gat));
  NAND3_X1  g712(.A1(new_n906), .A2(new_n317), .A3(new_n567), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n911), .A2(new_n567), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n317), .ZN(G1349gat));
  AND3_X1   g715(.A1(new_n588), .A2(new_n298), .A3(new_n299), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n906), .A2(new_n917), .ZN(new_n918));
  AOI211_X1 g717(.A(new_n810), .B(new_n910), .C1(new_n812), .C2(new_n818), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n286), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT123), .B1(new_n920), .B2(KEYINPUT60), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n811), .A2(KEYINPUT112), .A3(new_n481), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n817), .B1(new_n816), .B2(new_n452), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n588), .B(new_n909), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n924), .A2(G183gat), .B1(new_n906), .B2(new_n917), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n920), .A2(new_n930), .A3(KEYINPUT60), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT122), .B1(new_n925), .B2(new_n927), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n929), .A2(new_n933), .ZN(G1350gat));
  NAND2_X1  g733(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G190gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n911), .B2(new_n678), .ZN(new_n937));
  NOR2_X1   g736(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n937), .B(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n689), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n906), .A2(new_n300), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1351gat));
  NOR2_X1   g741(.A1(new_n665), .A2(new_n908), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n872), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n944), .A2(G197gat), .A3(new_n652), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n727), .B(new_n943), .C1(new_n884), .C2(new_n888), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(G197gat), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT125), .ZN(G1352gat));
  INV_X1    g747(.A(new_n944), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950));
  AOI21_X1  g749(.A(G204gat), .B1(new_n950), .B2(KEYINPUT62), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n949), .A2(new_n567), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n890), .A2(new_n943), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G204gat), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1353gat));
  OR3_X1    g756(.A1(new_n944), .A2(G211gat), .A3(new_n810), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n588), .B(new_n943), .C1(new_n884), .C2(new_n888), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT127), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n964), .B(new_n958), .C1(new_n960), .C2(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1354gat));
  INV_X1    g765(.A(G218gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n967), .A3(new_n940), .ZN(new_n968));
  NOR4_X1   g767(.A1(new_n889), .A2(new_n665), .A3(new_n626), .A4(new_n908), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(new_n967), .ZN(G1355gat));
endmodule


