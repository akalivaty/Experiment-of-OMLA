//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(KEYINPUT71), .A3(KEYINPUT23), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT71), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G128), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n190), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n189), .B1(new_n195), .B2(new_n188), .ZN(new_n196));
  INV_X1    g010(.A(new_n188), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(KEYINPUT70), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n192), .A2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  XOR2_X1   g015(.A(KEYINPUT24), .B(G110), .Z(new_n202));
  OAI22_X1  g016(.A1(new_n196), .A2(G110), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT72), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n206), .A3(G125), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n204), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G140), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(KEYINPUT16), .ZN(new_n214));
  OAI21_X1  g028(.A(G146), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(G140), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n208), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n203), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT72), .B1(new_n212), .B2(G140), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n210), .B1(new_n220), .B2(new_n213), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n214), .B1(new_n221), .B2(KEYINPUT16), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n217), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n196), .A2(G110), .B1(new_n201), .B2(new_n202), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(KEYINPUT73), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT73), .B1(new_n224), .B2(new_n225), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n219), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT22), .B(G137), .ZN(new_n230));
  INV_X1    g044(.A(G953), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n231), .A2(G221), .A3(G234), .ZN(new_n232));
  XOR2_X1   g046(.A(new_n230), .B(new_n232), .Z(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n219), .B(new_n233), .C1(new_n227), .C2(new_n228), .ZN(new_n236));
  INV_X1    g050(.A(G217), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(G234), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G902), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n235), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n241), .B(KEYINPUT74), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n235), .A2(new_n238), .A3(new_n236), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT25), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n235), .A2(new_n245), .A3(new_n238), .A4(new_n236), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n246), .A3(new_n239), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n242), .A2(KEYINPUT75), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT75), .B1(new_n242), .B2(new_n247), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n191), .A2(G116), .ZN(new_n252));
  INV_X1    g066(.A(G116), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G119), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT2), .B(G113), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n255), .B(new_n256), .Z(new_n257));
  NAND2_X1  g071(.A1(new_n217), .A2(G143), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G128), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G137), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n264), .A2(G137), .ZN(new_n267));
  OAI21_X1  g081(.A(G131), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT11), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n264), .B2(G137), .ZN(new_n270));
  INV_X1    g084(.A(G137), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT11), .A3(G134), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n270), .A2(new_n272), .A3(new_n273), .A4(new_n265), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n258), .B(new_n260), .C1(KEYINPUT1), .C2(new_n187), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n263), .A2(new_n268), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n270), .A2(new_n272), .A3(new_n265), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G131), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n278), .A2(new_n274), .ZN(new_n279));
  XNOR2_X1  g093(.A(G143), .B(G146), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT0), .B(G128), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT64), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT0), .A2(G128), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT64), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n261), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n280), .A2(new_n283), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n282), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n257), .B(new_n276), .C1(new_n279), .C2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n290), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n261), .A2(new_n285), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n295), .A2(KEYINPUT64), .B1(new_n280), .B2(new_n283), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n278), .A2(new_n274), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n287), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n257), .B1(new_n298), .B2(new_n276), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT28), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n293), .B1(new_n300), .B2(KEYINPUT66), .ZN(new_n301));
  NOR2_X1   g115(.A1(G237), .A2(G953), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G210), .ZN(new_n303));
  INV_X1    g117(.A(G101), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n292), .A2(new_n308), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n301), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT30), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT65), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n276), .B(new_n312), .C1(new_n279), .C2(new_n289), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n311), .A2(KEYINPUT65), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n314), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n298), .A2(new_n276), .A3(new_n312), .A4(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n257), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n307), .B1(new_n318), .B2(new_n294), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n251), .B1(new_n310), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n276), .B1(new_n279), .B2(new_n289), .ZN(new_n323));
  INV_X1    g137(.A(new_n257), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n291), .B1(new_n325), .B2(new_n290), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n292), .B1(new_n326), .B2(new_n308), .ZN(new_n327));
  INV_X1    g141(.A(new_n307), .ZN(new_n328));
  INV_X1    g142(.A(new_n309), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n327), .A2(KEYINPUT29), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n330), .A2(new_n238), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n332), .A2(KEYINPUT68), .A3(new_n320), .A4(new_n319), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n322), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G472), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT69), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT69), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n337), .A3(G472), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n318), .A2(new_n307), .A3(new_n294), .ZN(new_n340));
  AOI21_X1  g154(.A(G902), .B1(new_n340), .B2(KEYINPUT31), .ZN(new_n341));
  INV_X1    g155(.A(G472), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n328), .B1(new_n327), .B2(new_n329), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n315), .A2(new_n317), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n324), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n328), .A3(new_n290), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT31), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT32), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n307), .B1(new_n301), .B2(new_n309), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(new_n347), .A3(new_n346), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(KEYINPUT32), .A3(new_n342), .A4(new_n341), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(KEYINPUT67), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT67), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n349), .A2(new_n356), .A3(new_n350), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n250), .B1(new_n339), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n231), .A2(G227), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT76), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G140), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(KEYINPUT77), .A2(G104), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT78), .A2(G107), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(KEYINPUT78), .A2(G107), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n367), .B(new_n368), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G107), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G104), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(G104), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n374), .B1(KEYINPUT3), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n376), .A3(new_n304), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n372), .A2(new_n376), .A3(KEYINPUT80), .A4(new_n304), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n263), .A2(new_n275), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  OR2_X1    g197(.A1(KEYINPUT78), .A2(G107), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(new_n369), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n384), .A2(KEYINPUT81), .A3(new_n385), .A4(new_n369), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n375), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G101), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n381), .A2(KEYINPUT10), .A3(new_n383), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT82), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n379), .A2(new_n380), .B1(G101), .B2(new_n390), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT10), .A4(new_n383), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n380), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n385), .A2(G107), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n385), .A2(G107), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(new_n366), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n384), .A2(new_n369), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n367), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n399), .B1(new_n404), .B2(new_n304), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n372), .A2(new_n376), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n406), .A2(KEYINPUT79), .A3(KEYINPUT4), .A4(G101), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n398), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n289), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n381), .A2(new_n383), .A3(new_n391), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT10), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n408), .A2(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n397), .A2(new_n279), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT12), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n279), .B1(KEYINPUT83), .B2(new_n414), .ZN(new_n415));
  AOI221_X4 g229(.A(new_n382), .B1(new_n390), .B2(G101), .C1(new_n379), .C2(new_n380), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n383), .B1(new_n381), .B2(new_n391), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n414), .A2(KEYINPUT83), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI221_X1 g234(.A(new_n415), .B1(KEYINPUT83), .B2(new_n414), .C1(new_n416), .C2(new_n417), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n364), .B1(new_n413), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n397), .A2(new_n412), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n297), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n397), .A2(new_n412), .A3(new_n279), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n363), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G469), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n423), .A2(new_n427), .A3(new_n428), .A4(new_n238), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n238), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n363), .B1(new_n413), .B2(new_n422), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n425), .A2(new_n364), .A3(new_n426), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(G469), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G221), .ZN(new_n436));
  XOR2_X1   g250(.A(KEYINPUT9), .B(G234), .Z(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(new_n238), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G214), .B1(G237), .B2(G902), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G210), .B1(G237), .B2(G902), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n445));
  XOR2_X1   g259(.A(G110), .B(G122), .Z(new_n446));
  AOI22_X1  g260(.A1(new_n406), .A2(G101), .B1(KEYINPUT79), .B2(KEYINPUT4), .ZN(new_n447));
  AOI211_X1 g261(.A(new_n304), .B(new_n399), .C1(new_n372), .C2(new_n376), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n257), .B1(new_n449), .B2(new_n398), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n255), .A2(new_n256), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n452), .A2(G113), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n252), .A2(new_n254), .A3(KEYINPUT5), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n381), .A2(new_n391), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n446), .B1(new_n450), .B2(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n380), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n405), .A2(new_n407), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n324), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n394), .A2(new_n455), .ZN(new_n461));
  INV_X1    g275(.A(new_n446), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n457), .A2(new_n463), .A3(KEYINPUT6), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n465), .B(new_n446), .C1(new_n450), .C2(new_n456), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n445), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n408), .A2(new_n324), .B1(new_n394), .B2(new_n455), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n465), .B1(new_n468), .B2(new_n462), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT84), .B1(new_n469), .B2(new_n457), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n289), .A2(G125), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n382), .A2(new_n212), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G224), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(G953), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n473), .A2(new_n475), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n467), .A2(new_n470), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n394), .ZN(new_n481));
  OR3_X1    g295(.A1(new_n481), .A2(KEYINPUT85), .A3(new_n455), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n455), .B1(new_n481), .B2(KEYINPUT85), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n446), .B(KEYINPUT8), .Z(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n486));
  OR3_X1    g300(.A1(new_n473), .A2(new_n486), .A3(new_n475), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n473), .B1(new_n486), .B2(new_n475), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n485), .A2(new_n463), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n238), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n444), .B1(new_n480), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n464), .A2(new_n445), .ZN(new_n492));
  INV_X1    g306(.A(new_n466), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n457), .B2(new_n469), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n492), .B(new_n478), .C1(new_n494), .C2(new_n445), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n489), .A2(new_n238), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n443), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n442), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n440), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(G475), .A2(G902), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n502));
  INV_X1    g316(.A(G237), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n231), .A3(G214), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n259), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n302), .A2(G143), .A3(G214), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n273), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT87), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n509));
  INV_X1    g323(.A(new_n506), .ZN(new_n510));
  AOI21_X1  g324(.A(G143), .B1(new_n302), .B2(G214), .ZN(new_n511));
  OAI21_X1  g325(.A(G131), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n505), .A2(new_n513), .A3(new_n273), .A4(new_n506), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n508), .A2(new_n509), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n505), .A2(new_n506), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT17), .A3(G131), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n515), .A2(new_n223), .A3(new_n215), .A4(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G113), .B(G122), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(new_n385), .ZN(new_n520));
  OAI211_X1 g334(.A(KEYINPUT18), .B(G131), .C1(new_n510), .C2(new_n511), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT86), .ZN(new_n522));
  INV_X1    g336(.A(new_n221), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n218), .B1(new_n523), .B2(new_n217), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT86), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n516), .A2(new_n525), .A3(KEYINPUT18), .A4(G131), .ZN(new_n526));
  NAND2_X1  g340(.A1(KEYINPUT18), .A2(G131), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n505), .A2(new_n506), .A3(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n522), .A2(new_n524), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n518), .A2(new_n520), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n508), .A2(new_n512), .A3(new_n514), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT19), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n208), .A2(new_n216), .A3(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n217), .B(new_n533), .C1(new_n523), .C2(new_n532), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n215), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n520), .B1(new_n535), .B2(new_n529), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n502), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n529), .ZN(new_n538));
  INV_X1    g352(.A(new_n520), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n518), .A2(new_n520), .A3(new_n529), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(KEYINPUT88), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n501), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT20), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT89), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n540), .A2(KEYINPUT88), .A3(new_n541), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT88), .B1(new_n540), .B2(new_n541), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n500), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT20), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n544), .B(new_n500), .C1(new_n530), .C2(new_n536), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n545), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n520), .B1(new_n518), .B2(new_n529), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n238), .B1(new_n530), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT90), .B(G475), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n552), .A2(KEYINPUT91), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT91), .B1(new_n552), .B2(new_n556), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n253), .A2(G122), .ZN(new_n560));
  INV_X1    g374(.A(G122), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G116), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n560), .A2(new_n562), .A3(KEYINPUT92), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n384), .A2(new_n369), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n560), .A2(KEYINPUT14), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n562), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n560), .A2(KEYINPUT14), .ZN(new_n572));
  OAI21_X1  g386(.A(G107), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G128), .B(G143), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(new_n264), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n569), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT94), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n569), .A2(new_n578), .A3(new_n573), .A4(new_n575), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n567), .B(new_n568), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n574), .A2(new_n264), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n187), .A2(G143), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n187), .A2(G143), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(KEYINPUT13), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n585), .A2(KEYINPUT93), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(KEYINPUT93), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n584), .A2(KEYINPUT13), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n581), .B(new_n582), .C1(new_n264), .C2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n437), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n591), .A2(new_n237), .A3(G953), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n580), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n592), .B1(new_n580), .B2(new_n590), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n238), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G478), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(KEYINPUT15), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n595), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n231), .A2(G952), .ZN(new_n601));
  NAND2_X1  g415(.A1(G234), .A2(G237), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(G902), .A3(G953), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT95), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT21), .B(G898), .Z(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n604), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n600), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT96), .B1(new_n559), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n552), .A2(new_n556), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT91), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n552), .A2(KEYINPUT91), .A3(new_n556), .ZN(new_n616));
  AND4_X1   g430(.A1(KEYINPUT96), .A2(new_n615), .A3(new_n616), .A4(new_n611), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n359), .B(new_n499), .C1(new_n612), .C2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  OAI21_X1  g433(.A(new_n341), .B1(new_n343), .B2(new_n348), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G472), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n349), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n248), .B2(new_n249), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n435), .A2(new_n439), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT97), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n242), .A2(new_n247), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT75), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n242), .A2(KEYINPUT75), .A3(new_n247), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT97), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(new_n440), .A3(new_n632), .A4(new_n623), .ZN(new_n633));
  INV_X1    g447(.A(new_n610), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n498), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n626), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(new_n593), .B2(new_n594), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n637), .B(KEYINPUT33), .C1(new_n593), .C2(new_n594), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(G478), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n596), .A2(new_n238), .ZN(new_n643));
  INV_X1    g457(.A(new_n595), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n643), .B1(new_n644), .B2(new_n596), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT99), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n642), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n650), .B1(new_n557), .B2(new_n558), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n636), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT34), .B(G104), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT100), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n652), .B(new_n654), .ZN(G6));
  OAI211_X1 g469(.A(new_n545), .B(new_n550), .C1(KEYINPUT20), .C2(new_n548), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n556), .A3(new_n600), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n636), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT35), .B(G107), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  OR2_X1    g474(.A1(new_n234), .A2(KEYINPUT36), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n229), .B(new_n661), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n240), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n622), .B1(new_n247), .B2(new_n663), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n499), .B(new_n664), .C1(new_n612), .C2(new_n617), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND2_X1  g481(.A1(new_n247), .A2(new_n663), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n440), .A2(new_n498), .A3(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n334), .A2(new_n337), .A3(G472), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n337), .B1(new_n334), .B2(G472), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n358), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n603), .B(KEYINPUT101), .Z(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(new_n607), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n657), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n669), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XNOR2_X1  g492(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n675), .B(new_n679), .Z(new_n680));
  AND2_X1   g494(.A1(new_n440), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n328), .B1(new_n325), .B2(new_n290), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT102), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n238), .B1(new_n685), .B2(new_n340), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(G472), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT103), .B1(new_n358), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n689));
  INV_X1    g503(.A(new_n687), .ZN(new_n690));
  AOI211_X1 g504(.A(new_n689), .B(new_n690), .C1(new_n355), .C2(new_n357), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n668), .A2(new_n442), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n600), .B(new_n693), .C1(new_n557), .C2(new_n558), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n491), .A2(new_n497), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT38), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR4_X1   g511(.A1(new_n683), .A2(new_n692), .A3(new_n694), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n259), .ZN(G45));
  INV_X1    g513(.A(new_n675), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n650), .B(new_n700), .C1(new_n557), .C2(new_n558), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n669), .A3(new_n672), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT106), .B(G146), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G48));
  INV_X1    g519(.A(new_n651), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n423), .A2(new_n238), .A3(new_n427), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G469), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n439), .A3(new_n429), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT107), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n708), .A2(new_n711), .A3(new_n439), .A4(new_n429), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n359), .A2(new_n706), .A3(new_n635), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND3_X1  g530(.A1(new_n710), .A2(new_n498), .A3(new_n712), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n336), .A2(new_n338), .B1(new_n357), .B2(new_n355), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n250), .A2(new_n610), .A3(new_n657), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  OAI211_X1 g536(.A(new_n719), .B(new_n668), .C1(new_n612), .C2(new_n617), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NAND2_X1  g538(.A1(new_n615), .A2(new_n616), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n725), .A2(new_n600), .A3(new_n498), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n622), .A2(new_n627), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n634), .A3(new_n713), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NAND4_X1  g543(.A1(new_n702), .A2(new_n713), .A3(new_n498), .A4(new_n664), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  INV_X1    g545(.A(new_n349), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n733), .A3(KEYINPUT32), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n354), .A2(KEYINPUT109), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n734), .A2(new_n351), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n627), .B1(new_n339), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n432), .B2(new_n433), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n279), .B1(new_n397), .B2(new_n412), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n413), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT108), .B1(new_n741), .B2(new_n364), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n739), .A2(new_n742), .A3(new_n428), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n429), .A2(new_n431), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n439), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n491), .A2(new_n441), .A3(new_n497), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n737), .A2(KEYINPUT42), .A3(new_n702), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n746), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n739), .A2(new_n742), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(G469), .ZN(new_n753));
  INV_X1    g567(.A(new_n744), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n751), .A2(new_n755), .A3(new_n439), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n737), .A3(KEYINPUT110), .A4(new_n702), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n359), .A2(new_n702), .A3(new_n747), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n757), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n750), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  NAND4_X1  g577(.A1(new_n747), .A2(new_n672), .A3(new_n631), .A4(new_n676), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n359), .A2(KEYINPUT111), .A3(new_n676), .A4(new_n747), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  NAND2_X1  g583(.A1(new_n752), .A2(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n432), .A2(new_n433), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n428), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n430), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n429), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n439), .B(new_n680), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT112), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n650), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n725), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n780), .B(new_n781), .C1(new_n725), .C2(new_n783), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n622), .A2(new_n668), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n779), .B1(new_n789), .B2(KEYINPUT44), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(KEYINPUT44), .A3(new_n788), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT113), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n787), .A2(new_n793), .A3(KEYINPUT44), .A4(new_n788), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n751), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n792), .A2(KEYINPUT114), .A3(new_n751), .A4(new_n794), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n790), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g613(.A(KEYINPUT115), .B(G137), .Z(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(G39));
  OAI21_X1  g615(.A(new_n439), .B1(new_n776), .B2(new_n777), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT47), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT47), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n804), .B(new_n439), .C1(new_n776), .C2(new_n777), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n672), .A2(new_n701), .A3(new_n631), .A4(new_n746), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  NAND2_X1  g622(.A1(new_n708), .A2(new_n429), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(KEYINPUT49), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(KEYINPUT49), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n242), .A2(new_n247), .A3(new_n441), .A4(new_n439), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n692), .A2(new_n697), .A3(new_n784), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n672), .B(new_n669), .C1(new_n702), .C2(new_n676), .ZN(new_n816));
  INV_X1    g630(.A(new_n694), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n695), .A2(new_n700), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n745), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n817), .B(new_n819), .C1(new_n688), .C2(new_n691), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n820), .A3(new_n730), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT52), .ZN(new_n822));
  INV_X1    g636(.A(new_n600), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n651), .B1(new_n725), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n626), .A3(new_n633), .A4(new_n635), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n618), .A2(new_n665), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n746), .A2(new_n625), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n600), .A2(new_n675), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n556), .A2(new_n828), .A3(new_n668), .A4(new_n656), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n670), .A2(new_n671), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n355), .A2(new_n357), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n827), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n725), .A2(new_n650), .A3(new_n664), .A4(new_n700), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(new_n756), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n766), .B2(new_n767), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n816), .A2(new_n820), .A3(new_n730), .A4(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n822), .A2(new_n826), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n728), .A2(new_n721), .A3(new_n714), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n762), .A2(new_n723), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(KEYINPUT53), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(KEYINPUT53), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n815), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n837), .A2(new_n822), .A3(new_n826), .A4(new_n835), .ZN(new_n845));
  INV_X1    g659(.A(new_n840), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n826), .A2(new_n835), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(KEYINPUT116), .A3(new_n837), .A4(new_n822), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n847), .A2(KEYINPUT53), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT53), .B1(new_n838), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n841), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT54), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n844), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n787), .A2(new_n673), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n713), .A2(new_n751), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT119), .Z(new_n858));
  AND2_X1   g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(KEYINPUT48), .A3(new_n737), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n250), .A2(new_n603), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n858), .A2(new_n692), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n706), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n856), .A2(new_n727), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n863), .B(new_n601), .C1(new_n717), .C2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT48), .B1(new_n859), .B2(new_n737), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(KEYINPUT50), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n713), .A2(new_n442), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n696), .B1(new_n870), .B2(KEYINPUT117), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(KEYINPUT117), .B2(new_n870), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n864), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n869), .B1(new_n864), .B2(new_n872), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n864), .A2(new_n746), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n803), .A2(new_n805), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n809), .A2(new_n439), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n862), .A2(new_n559), .A3(new_n783), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n859), .A2(new_n664), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n875), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n860), .B(new_n867), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n855), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(G952), .A2(G953), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n814), .B1(new_n886), .B2(new_n887), .ZN(G75));
  XOR2_X1   g702(.A(new_n478), .B(KEYINPUT55), .Z(new_n889));
  NAND4_X1  g703(.A1(new_n850), .A2(G210), .A3(G902), .A4(new_n853), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n492), .B1(new_n494), .B2(new_n445), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT120), .Z(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n890), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n894), .B1(new_n890), .B2(new_n891), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n889), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n890), .A2(new_n891), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n893), .ZN(new_n900));
  INV_X1    g714(.A(new_n889), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n895), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n231), .A2(G952), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n898), .A2(new_n902), .A3(new_n904), .ZN(G51));
  AOI211_X1 g719(.A(new_n840), .B(new_n838), .C1(new_n851), .C2(KEYINPUT53), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n852), .A2(new_n841), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n815), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n850), .A2(KEYINPUT54), .A3(new_n853), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(KEYINPUT121), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n850), .A2(new_n853), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n912), .A3(new_n815), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n430), .B(KEYINPUT57), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n423), .A2(new_n427), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT122), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n911), .A2(new_n238), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n770), .A3(new_n773), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n903), .B1(new_n918), .B2(new_n920), .ZN(G54));
  NAND3_X1  g735(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n537), .A2(new_n542), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n922), .A2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n903), .ZN(G60));
  AND2_X1   g741(.A1(new_n640), .A2(new_n641), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n643), .B(KEYINPUT59), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n910), .A2(new_n913), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n910), .A2(new_n933), .A3(new_n913), .A4(new_n930), .ZN(new_n934));
  INV_X1    g748(.A(new_n929), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n844), .B2(new_n854), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n903), .B1(new_n936), .B2(new_n928), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n932), .A2(new_n934), .A3(new_n937), .ZN(G63));
  NOR2_X1   g752(.A1(new_n906), .A2(new_n907), .ZN(new_n939));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT60), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n235), .A2(new_n236), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n939), .A2(new_n662), .A3(new_n941), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n904), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n944), .A2(KEYINPUT61), .A3(new_n904), .A4(new_n945), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(G66));
  NAND3_X1  g764(.A1(new_n826), .A2(new_n839), .A3(new_n723), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n231), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT124), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n609), .B2(new_n474), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n893), .B1(G898), .B2(new_n231), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  OAI21_X1  g771(.A(new_n533), .B1(new_n523), .B2(new_n532), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n344), .B(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(G227), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n231), .B1(new_n961), .B2(G900), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n726), .A2(new_n737), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT126), .B1(new_n778), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n807), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n816), .A2(new_n730), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n762), .A2(new_n768), .A3(new_n966), .ZN(new_n967));
  OR3_X1    g781(.A1(new_n778), .A2(KEYINPUT126), .A3(new_n963), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n231), .B1(new_n799), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n959), .B1(new_n960), .B2(G953), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n962), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n797), .A2(new_n798), .ZN(new_n974));
  INV_X1    g788(.A(new_n790), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n824), .A2(new_n359), .A3(new_n681), .A4(new_n751), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n977), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n799), .A2(KEYINPUT125), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n966), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n698), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n807), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n959), .A2(new_n231), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n972), .B1(new_n986), .B2(new_n987), .ZN(G72));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n799), .A2(new_n951), .A3(new_n969), .ZN(new_n990));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n989), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n951), .ZN(new_n995));
  INV_X1    g809(.A(new_n969), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n976), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(KEYINPUT127), .A3(new_n992), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n318), .A2(new_n294), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(new_n328), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n994), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n842), .A2(new_n843), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n993), .B1(new_n346), .B2(new_n319), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n903), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1000), .A2(new_n328), .ZN(new_n1007));
  INV_X1    g821(.A(new_n985), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n995), .B(new_n1008), .C1(new_n978), .C2(new_n980), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1007), .B1(new_n1009), .B2(new_n992), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1006), .A2(new_n1010), .ZN(G57));
endmodule


