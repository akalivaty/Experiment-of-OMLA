

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n759), .A2(n758), .ZN(n760) );
  AND2_X2 U550 ( .A1(n517), .A2(G2105), .ZN(n593) );
  INV_X1 U551 ( .A(KEYINPUT103), .ZN(n708) );
  XNOR2_X1 U552 ( .A(n709), .B(n708), .ZN(n716) );
  INV_X1 U553 ( .A(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U554 ( .A(n723), .B(n722), .ZN(n727) );
  INV_X1 U555 ( .A(KEYINPUT105), .ZN(n741) );
  XNOR2_X1 U556 ( .A(n694), .B(KEYINPUT64), .ZN(n695) );
  NOR2_X1 U557 ( .A1(G164), .A2(G1384), .ZN(n692) );
  NOR2_X1 U558 ( .A1(G651), .A2(n620), .ZN(n641) );
  XNOR2_X1 U559 ( .A(G2104), .B(KEYINPUT65), .ZN(n517) );
  NAND2_X1 U560 ( .A1(G126), .A2(n593), .ZN(n515) );
  AND2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n882) );
  NAND2_X1 U562 ( .A1(G114), .A2(n882), .ZN(n514) );
  NAND2_X1 U563 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U564 ( .A(n516), .B(KEYINPUT90), .ZN(n522) );
  NOR2_X2 U565 ( .A1(n517), .A2(G2105), .ZN(n879) );
  NAND2_X1 U566 ( .A1(n879), .A2(G102), .ZN(n520) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n518), .Z(n878) );
  NAND2_X1 U569 ( .A1(n878), .A2(G138), .ZN(n519) );
  NAND2_X1 U570 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U571 ( .A1(n522), .A2(n521), .ZN(G164) );
  NAND2_X1 U572 ( .A1(G137), .A2(n878), .ZN(n523) );
  XNOR2_X1 U573 ( .A(n523), .B(KEYINPUT66), .ZN(n676) );
  NAND2_X1 U574 ( .A1(G101), .A2(n879), .ZN(n524) );
  XOR2_X1 U575 ( .A(KEYINPUT23), .B(n524), .Z(n675) );
  AND2_X1 U576 ( .A1(n676), .A2(n675), .ZN(n527) );
  NAND2_X1 U577 ( .A1(G125), .A2(n593), .ZN(n526) );
  NAND2_X1 U578 ( .A1(G113), .A2(n882), .ZN(n525) );
  AND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n673) );
  AND2_X1 U580 ( .A1(n527), .A2(n673), .ZN(G160) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n620) );
  NAND2_X1 U582 ( .A1(n641), .A2(G52), .ZN(n530) );
  XNOR2_X1 U583 ( .A(KEYINPUT67), .B(G651), .ZN(n531) );
  NOR2_X1 U584 ( .A1(G543), .A2(n531), .ZN(n528) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n528), .Z(n637) );
  NAND2_X1 U586 ( .A1(G64), .A2(n637), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n530), .A2(n529), .ZN(n537) );
  NOR2_X1 U588 ( .A1(n620), .A2(n531), .ZN(n633) );
  NAND2_X1 U589 ( .A1(G77), .A2(n633), .ZN(n532) );
  XNOR2_X1 U590 ( .A(n532), .B(KEYINPUT70), .ZN(n534) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n632) );
  NAND2_X1 U592 ( .A1(G90), .A2(n632), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U594 ( .A(KEYINPUT9), .B(n535), .Z(n536) );
  NOR2_X1 U595 ( .A1(n537), .A2(n536), .ZN(G171) );
  AND2_X1 U596 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U597 ( .A(G108), .ZN(G238) );
  INV_X1 U598 ( .A(G132), .ZN(G219) );
  INV_X1 U599 ( .A(G82), .ZN(G220) );
  NAND2_X1 U600 ( .A1(n641), .A2(G50), .ZN(n539) );
  NAND2_X1 U601 ( .A1(G62), .A2(n637), .ZN(n538) );
  NAND2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U603 ( .A(KEYINPUT83), .B(n540), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n633), .A2(G75), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n632), .A2(G88), .ZN(n541) );
  AND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(G303) );
  NAND2_X1 U608 ( .A1(G7), .A2(G661), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n545), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U610 ( .A(G223), .ZN(n815) );
  NAND2_X1 U611 ( .A1(n815), .A2(G567), .ZN(n546) );
  XOR2_X1 U612 ( .A(KEYINPUT11), .B(n546), .Z(G234) );
  NAND2_X1 U613 ( .A1(G81), .A2(n632), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(KEYINPUT12), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(KEYINPUT72), .ZN(n550) );
  NAND2_X1 U616 ( .A1(G68), .A2(n633), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT13), .B(n551), .ZN(n557) );
  NAND2_X1 U619 ( .A1(n637), .A2(G56), .ZN(n552) );
  XOR2_X1 U620 ( .A(KEYINPUT14), .B(n552), .Z(n555) );
  NAND2_X1 U621 ( .A1(G43), .A2(n641), .ZN(n553) );
  XNOR2_X1 U622 ( .A(KEYINPUT73), .B(n553), .ZN(n554) );
  NOR2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n931) );
  INV_X1 U625 ( .A(G860), .ZN(n606) );
  OR2_X1 U626 ( .A1(n931), .A2(n606), .ZN(G153) );
  INV_X1 U627 ( .A(G171), .ZN(G301) );
  NAND2_X1 U628 ( .A1(G868), .A2(G301), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G54), .A2(n641), .ZN(n564) );
  NAND2_X1 U630 ( .A1(n632), .A2(G92), .ZN(n559) );
  NAND2_X1 U631 ( .A1(G66), .A2(n637), .ZN(n558) );
  NAND2_X1 U632 ( .A1(n559), .A2(n558), .ZN(n562) );
  NAND2_X1 U633 ( .A1(n633), .A2(G79), .ZN(n560) );
  XOR2_X1 U634 ( .A(KEYINPUT74), .B(n560), .Z(n561) );
  NOR2_X1 U635 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U636 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U637 ( .A(n565), .B(KEYINPUT15), .ZN(n930) );
  OR2_X1 U638 ( .A1(n930), .A2(G868), .ZN(n566) );
  NAND2_X1 U639 ( .A1(n567), .A2(n566), .ZN(G284) );
  NAND2_X1 U640 ( .A1(n641), .A2(G53), .ZN(n569) );
  NAND2_X1 U641 ( .A1(G65), .A2(n637), .ZN(n568) );
  NAND2_X1 U642 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U643 ( .A1(n632), .A2(G91), .ZN(n571) );
  NAND2_X1 U644 ( .A1(G78), .A2(n633), .ZN(n570) );
  NAND2_X1 U645 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U646 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U647 ( .A(n574), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U648 ( .A1(n632), .A2(G89), .ZN(n575) );
  XNOR2_X1 U649 ( .A(n575), .B(KEYINPUT4), .ZN(n577) );
  NAND2_X1 U650 ( .A1(G76), .A2(n633), .ZN(n576) );
  NAND2_X1 U651 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U652 ( .A(n578), .B(KEYINPUT5), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n641), .A2(G51), .ZN(n580) );
  NAND2_X1 U654 ( .A1(G63), .A2(n637), .ZN(n579) );
  NAND2_X1 U655 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U656 ( .A(KEYINPUT6), .B(n581), .Z(n582) );
  NAND2_X1 U657 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U658 ( .A(n584), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U659 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U660 ( .A(G299), .ZN(n936) );
  INV_X1 U661 ( .A(G868), .ZN(n653) );
  NAND2_X1 U662 ( .A1(n936), .A2(n653), .ZN(n585) );
  XNOR2_X1 U663 ( .A(n585), .B(KEYINPUT75), .ZN(n587) );
  NOR2_X1 U664 ( .A1(n653), .A2(G286), .ZN(n586) );
  NOR2_X1 U665 ( .A1(n587), .A2(n586), .ZN(G297) );
  NAND2_X1 U666 ( .A1(n606), .A2(G559), .ZN(n588) );
  NAND2_X1 U667 ( .A1(n588), .A2(n930), .ZN(n589) );
  XNOR2_X1 U668 ( .A(n589), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n931), .ZN(n592) );
  NAND2_X1 U670 ( .A1(G868), .A2(n930), .ZN(n590) );
  NOR2_X1 U671 ( .A1(G559), .A2(n590), .ZN(n591) );
  NOR2_X1 U672 ( .A1(n592), .A2(n591), .ZN(G282) );
  NAND2_X1 U673 ( .A1(n593), .A2(G123), .ZN(n594) );
  XNOR2_X1 U674 ( .A(n594), .B(KEYINPUT18), .ZN(n596) );
  NAND2_X1 U675 ( .A1(G135), .A2(n878), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U677 ( .A(KEYINPUT76), .B(n597), .Z(n599) );
  NAND2_X1 U678 ( .A1(n879), .A2(G99), .ZN(n598) );
  NAND2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U680 ( .A1(G111), .A2(n882), .ZN(n600) );
  XNOR2_X1 U681 ( .A(KEYINPUT77), .B(n600), .ZN(n601) );
  NOR2_X1 U682 ( .A1(n602), .A2(n601), .ZN(n975) );
  XNOR2_X1 U683 ( .A(G2096), .B(n975), .ZN(n604) );
  INV_X1 U684 ( .A(G2100), .ZN(n603) );
  NAND2_X1 U685 ( .A1(n604), .A2(n603), .ZN(G156) );
  NAND2_X1 U686 ( .A1(G559), .A2(n930), .ZN(n605) );
  XOR2_X1 U687 ( .A(n931), .B(n605), .Z(n650) );
  NAND2_X1 U688 ( .A1(n606), .A2(n650), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G93), .A2(n632), .ZN(n608) );
  NAND2_X1 U690 ( .A1(G55), .A2(n641), .ZN(n607) );
  NAND2_X1 U691 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n637), .A2(G67), .ZN(n609) );
  XOR2_X1 U693 ( .A(KEYINPUT78), .B(n609), .Z(n610) );
  NOR2_X1 U694 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U695 ( .A1(G80), .A2(n633), .ZN(n612) );
  AND2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n652) );
  XOR2_X1 U697 ( .A(n614), .B(n652), .Z(G145) );
  NAND2_X1 U698 ( .A1(G74), .A2(G651), .ZN(n615) );
  XNOR2_X1 U699 ( .A(n615), .B(KEYINPUT80), .ZN(n618) );
  NAND2_X1 U700 ( .A1(G49), .A2(n641), .ZN(n616) );
  XOR2_X1 U701 ( .A(KEYINPUT79), .B(n616), .Z(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n637), .A2(n619), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n620), .A2(G87), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(G288) );
  NAND2_X1 U706 ( .A1(G73), .A2(n633), .ZN(n623) );
  XNOR2_X1 U707 ( .A(n623), .B(KEYINPUT2), .ZN(n625) );
  NAND2_X1 U708 ( .A1(G61), .A2(n637), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G86), .A2(n632), .ZN(n626) );
  XNOR2_X1 U711 ( .A(KEYINPUT81), .B(n626), .ZN(n627) );
  NOR2_X1 U712 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U713 ( .A(n629), .B(KEYINPUT82), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G48), .A2(n641), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(G305) );
  NAND2_X1 U716 ( .A1(n632), .A2(G85), .ZN(n635) );
  NAND2_X1 U717 ( .A1(G72), .A2(n633), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U719 ( .A(KEYINPUT68), .B(n636), .ZN(n640) );
  NAND2_X1 U720 ( .A1(G60), .A2(n637), .ZN(n638) );
  XNOR2_X1 U721 ( .A(KEYINPUT69), .B(n638), .ZN(n639) );
  NOR2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n641), .A2(G47), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(G290) );
  XNOR2_X1 U725 ( .A(KEYINPUT84), .B(G288), .ZN(n644) );
  XOR2_X1 U726 ( .A(n644), .B(n652), .Z(n647) );
  XNOR2_X1 U727 ( .A(n936), .B(G303), .ZN(n645) );
  XNOR2_X1 U728 ( .A(n645), .B(G305), .ZN(n646) );
  XNOR2_X1 U729 ( .A(n647), .B(n646), .ZN(n649) );
  XNOR2_X1 U730 ( .A(G290), .B(KEYINPUT19), .ZN(n648) );
  XNOR2_X1 U731 ( .A(n649), .B(n648), .ZN(n894) );
  XNOR2_X1 U732 ( .A(n650), .B(n894), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n651), .A2(G868), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U736 ( .A(KEYINPUT85), .B(n656), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n658) );
  XOR2_X1 U738 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n657) );
  XNOR2_X1 U739 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U744 ( .A1(G220), .A2(G219), .ZN(n662) );
  XOR2_X1 U745 ( .A(KEYINPUT22), .B(n662), .Z(n663) );
  NOR2_X1 U746 ( .A1(G218), .A2(n663), .ZN(n664) );
  XOR2_X1 U747 ( .A(KEYINPUT87), .B(n664), .Z(n665) );
  NAND2_X1 U748 ( .A1(G96), .A2(n665), .ZN(n820) );
  NAND2_X1 U749 ( .A1(n820), .A2(G2106), .ZN(n671) );
  NAND2_X1 U750 ( .A1(G120), .A2(G69), .ZN(n666) );
  XOR2_X1 U751 ( .A(KEYINPUT88), .B(n666), .Z(n667) );
  NAND2_X1 U752 ( .A1(G57), .A2(n667), .ZN(n668) );
  NOR2_X1 U753 ( .A1(G238), .A2(n668), .ZN(n669) );
  XNOR2_X1 U754 ( .A(KEYINPUT89), .B(n669), .ZN(n821) );
  NAND2_X1 U755 ( .A1(n821), .A2(G567), .ZN(n670) );
  NAND2_X1 U756 ( .A1(n671), .A2(n670), .ZN(n822) );
  NAND2_X1 U757 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U758 ( .A1(n822), .A2(n672), .ZN(n817) );
  NAND2_X1 U759 ( .A1(n817), .A2(G36), .ZN(G176) );
  AND2_X1 U760 ( .A1(G40), .A2(n673), .ZN(n674) );
  AND2_X1 U761 ( .A1(n675), .A2(n674), .ZN(n677) );
  NAND2_X1 U762 ( .A1(n677), .A2(n676), .ZN(n691) );
  NOR2_X1 U763 ( .A1(n692), .A2(n691), .ZN(n678) );
  XOR2_X1 U764 ( .A(KEYINPUT91), .B(n678), .Z(n810) );
  XNOR2_X1 U765 ( .A(KEYINPUT34), .B(KEYINPUT92), .ZN(n682) );
  NAND2_X1 U766 ( .A1(G140), .A2(n878), .ZN(n680) );
  NAND2_X1 U767 ( .A1(G104), .A2(n879), .ZN(n679) );
  NAND2_X1 U768 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U769 ( .A(n682), .B(n681), .ZN(n688) );
  XNOR2_X1 U770 ( .A(KEYINPUT93), .B(KEYINPUT35), .ZN(n686) );
  NAND2_X1 U771 ( .A1(G128), .A2(n593), .ZN(n684) );
  NAND2_X1 U772 ( .A1(G116), .A2(n882), .ZN(n683) );
  NAND2_X1 U773 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U774 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U775 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U776 ( .A(n689), .B(KEYINPUT36), .ZN(n690) );
  XNOR2_X1 U777 ( .A(n690), .B(KEYINPUT94), .ZN(n873) );
  XNOR2_X1 U778 ( .A(G2067), .B(KEYINPUT37), .ZN(n808) );
  NOR2_X1 U779 ( .A1(n873), .A2(n808), .ZN(n974) );
  NAND2_X1 U780 ( .A1(n810), .A2(n974), .ZN(n806) );
  INV_X1 U781 ( .A(n691), .ZN(n693) );
  NAND2_X1 U782 ( .A1(n693), .A2(n692), .ZN(n694) );
  BUF_X2 U783 ( .A(n695), .Z(n746) );
  NOR2_X1 U784 ( .A1(n746), .A2(G2084), .ZN(n729) );
  NAND2_X1 U785 ( .A1(G8), .A2(n729), .ZN(n744) );
  XNOR2_X1 U786 ( .A(G1996), .B(KEYINPUT101), .ZN(n918) );
  NOR2_X1 U787 ( .A1(n695), .A2(n918), .ZN(n696) );
  XOR2_X1 U788 ( .A(n696), .B(KEYINPUT26), .Z(n698) );
  NAND2_X1 U789 ( .A1(n746), .A2(G1341), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U791 ( .A1(n931), .A2(n699), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n705), .A2(n930), .ZN(n704) );
  AND2_X1 U793 ( .A1(n746), .A2(G1348), .ZN(n700) );
  XOR2_X1 U794 ( .A(n700), .B(KEYINPUT102), .Z(n702) );
  INV_X1 U795 ( .A(n746), .ZN(n711) );
  NAND2_X1 U796 ( .A1(n711), .A2(G2067), .ZN(n701) );
  NAND2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n707) );
  OR2_X1 U799 ( .A1(n930), .A2(n705), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U801 ( .A1(G2072), .A2(n711), .ZN(n710) );
  XNOR2_X1 U802 ( .A(KEYINPUT27), .B(n710), .ZN(n714) );
  XOR2_X1 U803 ( .A(G1956), .B(KEYINPUT98), .Z(n998) );
  NOR2_X1 U804 ( .A1(n998), .A2(n711), .ZN(n712) );
  XOR2_X1 U805 ( .A(KEYINPUT99), .B(n712), .Z(n713) );
  NOR2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U807 ( .A1(n717), .A2(n936), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n721) );
  NOR2_X1 U809 ( .A1(n717), .A2(n936), .ZN(n719) );
  XOR2_X1 U810 ( .A(KEYINPUT28), .B(KEYINPUT100), .Z(n718) );
  XNOR2_X1 U811 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n723) );
  AND2_X1 U813 ( .A1(n746), .A2(G1961), .ZN(n725) );
  XNOR2_X1 U814 ( .A(G2078), .B(KEYINPUT25), .ZN(n912) );
  NOR2_X1 U815 ( .A1(n746), .A2(n912), .ZN(n724) );
  NOR2_X1 U816 ( .A1(n725), .A2(n724), .ZN(n728) );
  NAND2_X1 U817 ( .A1(G171), .A2(n728), .ZN(n726) );
  NAND2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n738) );
  NOR2_X1 U819 ( .A1(G171), .A2(n728), .ZN(n735) );
  NAND2_X1 U820 ( .A1(G8), .A2(n746), .ZN(n772) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n772), .ZN(n739) );
  NOR2_X1 U822 ( .A1(n729), .A2(n739), .ZN(n730) );
  XNOR2_X1 U823 ( .A(KEYINPUT104), .B(n730), .ZN(n731) );
  NAND2_X1 U824 ( .A1(n731), .A2(G8), .ZN(n732) );
  XNOR2_X1 U825 ( .A(KEYINPUT30), .B(n732), .ZN(n733) );
  NOR2_X1 U826 ( .A1(G168), .A2(n733), .ZN(n734) );
  NOR2_X1 U827 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U828 ( .A(KEYINPUT31), .B(n736), .Z(n737) );
  NAND2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n745) );
  INV_X1 U830 ( .A(n745), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X1 U832 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n755) );
  NAND2_X1 U834 ( .A1(n745), .A2(G286), .ZN(n751) );
  NOR2_X1 U835 ( .A1(n746), .A2(G2090), .ZN(n748) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n772), .ZN(n747) );
  NOR2_X1 U837 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U838 ( .A1(n749), .A2(G303), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n752), .A2(G8), .ZN(n753) );
  XNOR2_X1 U841 ( .A(KEYINPUT32), .B(n753), .ZN(n754) );
  NAND2_X1 U842 ( .A1(n755), .A2(n754), .ZN(n771) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n761) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U845 ( .A1(n761), .A2(n756), .ZN(n942) );
  AND2_X1 U846 ( .A1(n771), .A2(n942), .ZN(n759) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n935) );
  INV_X1 U848 ( .A(n772), .ZN(n757) );
  NAND2_X1 U849 ( .A1(n935), .A2(n757), .ZN(n758) );
  NOR2_X1 U850 ( .A1(n760), .A2(KEYINPUT33), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n761), .A2(KEYINPUT33), .ZN(n762) );
  NOR2_X1 U852 ( .A1(n762), .A2(n772), .ZN(n763) );
  NOR2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n766) );
  XOR2_X1 U854 ( .A(G1981), .B(KEYINPUT106), .Z(n765) );
  XNOR2_X1 U855 ( .A(G305), .B(n765), .ZN(n948) );
  NAND2_X1 U856 ( .A1(n766), .A2(n948), .ZN(n777) );
  NOR2_X1 U857 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XOR2_X1 U858 ( .A(n767), .B(KEYINPUT24), .Z(n768) );
  OR2_X1 U859 ( .A1(n772), .A2(n768), .ZN(n775) );
  NOR2_X1 U860 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U861 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  AND2_X1 U866 ( .A1(n806), .A2(n778), .ZN(n799) );
  NAND2_X1 U867 ( .A1(G129), .A2(n593), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G117), .A2(n882), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U870 ( .A(n781), .B(KEYINPUT97), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G141), .A2(n878), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n879), .A2(G105), .ZN(n784) );
  XOR2_X1 U874 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n867) );
  INV_X1 U876 ( .A(G1996), .ZN(n800) );
  NOR2_X1 U877 ( .A1(n867), .A2(n800), .ZN(n796) );
  NAND2_X1 U878 ( .A1(G107), .A2(n882), .ZN(n788) );
  NAND2_X1 U879 ( .A1(G131), .A2(n878), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G95), .A2(n879), .ZN(n789) );
  XNOR2_X1 U882 ( .A(KEYINPUT95), .B(n789), .ZN(n790) );
  NOR2_X1 U883 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n593), .A2(G119), .ZN(n792) );
  NAND2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n869) );
  NAND2_X1 U886 ( .A1(G1991), .A2(n869), .ZN(n794) );
  XOR2_X1 U887 ( .A(KEYINPUT96), .B(n794), .Z(n795) );
  NOR2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n801) );
  XOR2_X1 U889 ( .A(G1986), .B(G290), .Z(n937) );
  NAND2_X1 U890 ( .A1(n801), .A2(n937), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n797), .A2(n810), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n813) );
  AND2_X1 U893 ( .A1(n800), .A2(n867), .ZN(n966) );
  INV_X1 U894 ( .A(n801), .ZN(n973) );
  NOR2_X1 U895 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U896 ( .A1(G1991), .A2(n869), .ZN(n976) );
  NOR2_X1 U897 ( .A1(n802), .A2(n976), .ZN(n803) );
  NOR2_X1 U898 ( .A1(n973), .A2(n803), .ZN(n804) );
  NOR2_X1 U899 ( .A1(n966), .A2(n804), .ZN(n805) );
  XNOR2_X1 U900 ( .A(KEYINPUT39), .B(n805), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n873), .A2(n808), .ZN(n963) );
  NAND2_X1 U903 ( .A1(n809), .A2(n963), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U906 ( .A(n814), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n815), .ZN(G217) );
  AND2_X1 U908 ( .A1(G15), .A2(G2), .ZN(n816) );
  NAND2_X1 U909 ( .A1(G661), .A2(n816), .ZN(G259) );
  NAND2_X1 U910 ( .A1(G1), .A2(G3), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U912 ( .A(n819), .B(KEYINPUT108), .ZN(G188) );
  XNOR2_X1 U913 ( .A(G69), .B(KEYINPUT109), .ZN(G235) );
  INV_X1 U915 ( .A(G120), .ZN(G236) );
  INV_X1 U916 ( .A(G96), .ZN(G221) );
  INV_X1 U917 ( .A(G57), .ZN(G237) );
  NOR2_X1 U918 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U919 ( .A(G325), .ZN(G261) );
  INV_X1 U920 ( .A(n822), .ZN(G319) );
  XNOR2_X1 U921 ( .A(G1348), .B(G2435), .ZN(n823) );
  XNOR2_X1 U922 ( .A(n823), .B(G2438), .ZN(n824) );
  XNOR2_X1 U923 ( .A(n824), .B(G1341), .ZN(n830) );
  XOR2_X1 U924 ( .A(G2451), .B(G2446), .Z(n826) );
  XNOR2_X1 U925 ( .A(G2427), .B(G2443), .ZN(n825) );
  XNOR2_X1 U926 ( .A(n826), .B(n825), .ZN(n828) );
  XOR2_X1 U927 ( .A(G2430), .B(G2454), .Z(n827) );
  XNOR2_X1 U928 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U929 ( .A(n830), .B(n829), .ZN(n831) );
  NAND2_X1 U930 ( .A1(n831), .A2(G14), .ZN(n832) );
  XNOR2_X1 U931 ( .A(KEYINPUT107), .B(n832), .ZN(G401) );
  XOR2_X1 U932 ( .A(KEYINPUT41), .B(G1956), .Z(n834) );
  XNOR2_X1 U933 ( .A(G1996), .B(G1991), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U935 ( .A(n835), .B(KEYINPUT111), .Z(n837) );
  XNOR2_X1 U936 ( .A(G1966), .B(G1981), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U938 ( .A(G1976), .B(G1971), .Z(n839) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1961), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U942 ( .A(KEYINPUT112), .B(G2474), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(G229) );
  XOR2_X1 U944 ( .A(G2096), .B(KEYINPUT43), .Z(n845) );
  XNOR2_X1 U945 ( .A(G2090), .B(G2678), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U947 ( .A(n846), .B(KEYINPUT110), .Z(n848) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U950 ( .A(KEYINPUT42), .B(G2100), .Z(n850) );
  XNOR2_X1 U951 ( .A(G2084), .B(G2078), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(G227) );
  NAND2_X1 U954 ( .A1(G112), .A2(n882), .ZN(n854) );
  NAND2_X1 U955 ( .A1(G136), .A2(n878), .ZN(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n593), .A2(G124), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U959 ( .A1(G100), .A2(n879), .ZN(n856) );
  NAND2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U961 ( .A1(n859), .A2(n858), .ZN(G162) );
  NAND2_X1 U962 ( .A1(G130), .A2(n593), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G118), .A2(n882), .ZN(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G142), .A2(n878), .ZN(n863) );
  NAND2_X1 U966 ( .A1(G106), .A2(n879), .ZN(n862) );
  NAND2_X1 U967 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U968 ( .A(n864), .B(KEYINPUT45), .Z(n865) );
  NOR2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n868) );
  XOR2_X1 U970 ( .A(n868), .B(n867), .Z(n877) );
  XNOR2_X1 U971 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n869), .B(KEYINPUT48), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(n872), .B(KEYINPUT114), .Z(n875) );
  XNOR2_X1 U975 ( .A(n873), .B(KEYINPUT115), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n891) );
  NAND2_X1 U978 ( .A1(G139), .A2(n878), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G103), .A2(n879), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n887) );
  NAND2_X1 U981 ( .A1(G127), .A2(n593), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G115), .A2(n882), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n959) );
  XOR2_X1 U986 ( .A(G162), .B(n959), .Z(n889) );
  XNOR2_X1 U987 ( .A(G164), .B(G160), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n892), .B(n975), .ZN(n893) );
  NOR2_X1 U991 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U992 ( .A(n931), .B(n894), .ZN(n896) );
  XNOR2_X1 U993 ( .A(G171), .B(n930), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U995 ( .A(G286), .B(n897), .Z(n898) );
  NOR2_X1 U996 ( .A1(G37), .A2(n898), .ZN(G397) );
  NOR2_X1 U997 ( .A1(G229), .A2(G227), .ZN(n900) );
  XNOR2_X1 U998 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(G401), .A2(n901), .ZN(n902) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n902), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(KEYINPUT117), .B(n903), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1006 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n983) );
  XNOR2_X1 U1007 ( .A(KEYINPUT54), .B(G34), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(n906), .B(KEYINPUT123), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(G2084), .B(n907), .ZN(n925) );
  XNOR2_X1 U1010 ( .A(G2090), .B(G35), .ZN(n923) );
  XNOR2_X1 U1011 ( .A(KEYINPUT121), .B(G2067), .ZN(n908) );
  XNOR2_X1 U1012 ( .A(n908), .B(G26), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(G1991), .B(G25), .ZN(n910) );
  XNOR2_X1 U1014 ( .A(G33), .B(G2072), .ZN(n909) );
  NOR2_X1 U1015 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1016 ( .A1(G28), .A2(n911), .ZN(n915) );
  XOR2_X1 U1017 ( .A(G27), .B(n912), .Z(n913) );
  XNOR2_X1 U1018 ( .A(KEYINPUT122), .B(n913), .ZN(n914) );
  NOR2_X1 U1019 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1020 ( .A1(n917), .A2(n916), .ZN(n920) );
  XOR2_X1 U1021 ( .A(G32), .B(n918), .Z(n919) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1023 ( .A(KEYINPUT53), .B(n921), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n983), .B(n926), .ZN(n928) );
  INV_X1 U1027 ( .A(G29), .ZN(n927) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(G11), .A2(n929), .ZN(n958) );
  XNOR2_X1 U1030 ( .A(G171), .B(G1961), .ZN(n947) );
  XNOR2_X1 U1031 ( .A(n930), .B(G1348), .ZN(n933) );
  XOR2_X1 U1032 ( .A(G1341), .B(n931), .Z(n932) );
  NAND2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n945) );
  NAND2_X1 U1034 ( .A1(G1971), .A2(G303), .ZN(n934) );
  NAND2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(n936), .B(G1956), .ZN(n938) );
  NAND2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1040 ( .A(KEYINPUT125), .B(n943), .Z(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G168), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(n950), .B(KEYINPUT57), .ZN(n951) );
  XOR2_X1 U1046 ( .A(KEYINPUT124), .B(n951), .Z(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n955) );
  XOR2_X1 U1048 ( .A(KEYINPUT56), .B(G16), .Z(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n956), .B(KEYINPUT126), .ZN(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n987) );
  XOR2_X1 U1052 ( .A(G2072), .B(n959), .Z(n961) );
  XOR2_X1 U1053 ( .A(G164), .B(G2078), .Z(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(KEYINPUT50), .B(n962), .ZN(n972) );
  XNOR2_X1 U1056 ( .A(G2084), .B(G160), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n970) );
  XOR2_X1 U1058 ( .A(G2090), .B(G162), .Z(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1060 ( .A(KEYINPUT51), .B(n967), .Z(n968) );
  XNOR2_X1 U1061 ( .A(n968), .B(KEYINPUT119), .ZN(n969) );
  NOR2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n981) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n979) );
  NOR2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(n977), .B(KEYINPUT118), .ZN(n978) );
  NAND2_X1 U1067 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1068 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1069 ( .A(KEYINPUT52), .B(n982), .ZN(n984) );
  NAND2_X1 U1070 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1071 ( .A1(n985), .A2(G29), .ZN(n986) );
  NAND2_X1 U1072 ( .A1(n987), .A2(n986), .ZN(n1012) );
  XOR2_X1 U1073 ( .A(G1986), .B(G24), .Z(n991) );
  XNOR2_X1 U1074 ( .A(G1971), .B(G22), .ZN(n989) );
  XNOR2_X1 U1075 ( .A(G23), .B(G1976), .ZN(n988) );
  NOR2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n993) );
  XNOR2_X1 U1078 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(n993), .B(n992), .ZN(n997) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G21), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G5), .B(G1961), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n1008) );
  XNOR2_X1 U1084 ( .A(n998), .B(G20), .ZN(n1002) );
  XNOR2_X1 U1085 ( .A(G1341), .B(G19), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(G1981), .B(G6), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1089 ( .A(KEYINPUT59), .B(G1348), .Z(n1003) );
  XNOR2_X1 U1090 ( .A(G4), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1092 ( .A(KEYINPUT60), .B(n1006), .Z(n1007) );
  NOR2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(KEYINPUT61), .B(n1009), .Z(n1010) );
  NOR2_X1 U1095 ( .A1(G16), .A2(n1010), .ZN(n1011) );
  NOR2_X1 U1096 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(n1013), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1098 ( .A(G311), .ZN(G150) );
  INV_X1 U1099 ( .A(G303), .ZN(G166) );
endmodule

