//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  XNOR2_X1  g000(.A(G119), .B(G128), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT24), .B(G110), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n192));
  INV_X1    g006(.A(G110), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT23), .B1(new_n194), .B2(G119), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT76), .B1(new_n196), .B2(G128), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n195), .B(new_n197), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n191), .A2(new_n192), .B1(new_n193), .B2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n192), .B2(new_n191), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n205));
  OR3_X1    g019(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G146), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n207), .B(KEYINPUT79), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n204), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT80), .B1(new_n209), .B2(G146), .ZN(new_n210));
  XNOR2_X1  g024(.A(G125), .B(G140), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT80), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n200), .A2(new_n208), .A3(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n198), .A2(new_n193), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n217), .B(KEYINPUT77), .ZN(new_n218));
  INV_X1    g032(.A(new_n207), .ZN(new_n219));
  AOI21_X1  g033(.A(G146), .B1(new_n205), .B2(new_n206), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n218), .B(new_n222), .C1(new_n189), .C2(new_n190), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT22), .B(G137), .ZN(new_n225));
  INV_X1    g039(.A(G221), .ZN(new_n226));
  INV_X1    g040(.A(G234), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n226), .A2(new_n227), .A3(G953), .ZN(new_n228));
  XOR2_X1   g042(.A(new_n225), .B(new_n228), .Z(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n216), .A2(new_n223), .A3(new_n229), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n233));
  AOI21_X1  g047(.A(G902), .B1(new_n233), .B2(KEYINPUT81), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n233), .A2(KEYINPUT81), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n236), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n231), .A2(new_n238), .A3(new_n232), .A4(new_n234), .ZN(new_n239));
  OAI21_X1  g053(.A(G217), .B1(new_n227), .B2(G902), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT74), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n237), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n231), .A2(new_n232), .ZN(new_n244));
  AOI21_X1  g058(.A(G902), .B1(new_n227), .B2(G217), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT72), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n196), .A2(G116), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(KEYINPUT66), .A2(G116), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT66), .A2(G116), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(G119), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT2), .B(G113), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n251), .A2(KEYINPUT67), .A3(G119), .A4(new_n252), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n257), .B1(new_n255), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n262));
  INV_X1    g076(.A(G137), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(G134), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G137), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n267), .B2(KEYINPUT11), .ZN(new_n268));
  INV_X1    g082(.A(G131), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT11), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n265), .B(new_n270), .C1(new_n266), .C2(G137), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n266), .A2(G137), .ZN(new_n273));
  OAI21_X1  g087(.A(G131), .B1(new_n273), .B2(new_n264), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n276));
  INV_X1    g090(.A(G143), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G146), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n213), .A2(G143), .ZN(new_n279));
  OAI22_X1  g093(.A1(new_n276), .A2(new_n278), .B1(new_n279), .B2(G128), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(G143), .B(G146), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT65), .A3(new_n276), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n280), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n262), .B1(new_n275), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n280), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT65), .B1(new_n284), .B2(new_n276), .ZN(new_n289));
  AND4_X1   g103(.A1(KEYINPUT65), .A2(new_n276), .A3(new_n278), .A4(new_n279), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n291), .A2(KEYINPUT69), .A3(new_n274), .A4(new_n272), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n278), .A2(new_n279), .A3(new_n294), .ZN(new_n295));
  OR2_X1    g109(.A1(KEYINPUT0), .A2(G128), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n294), .B1(new_n278), .B2(new_n279), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n293), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n298), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n300), .A2(KEYINPUT68), .A3(new_n296), .A4(new_n295), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n269), .B1(new_n268), .B2(new_n271), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n299), .B(new_n301), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n261), .A2(new_n287), .A3(new_n292), .A4(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n287), .A2(new_n292), .A3(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT30), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n291), .A2(new_n274), .A3(new_n272), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT30), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n302), .A2(new_n303), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n297), .A2(new_n298), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n310), .B(new_n311), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n261), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT26), .B(G101), .ZN(new_n316));
  NOR2_X1   g130(.A1(G237), .A2(G953), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G210), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n316), .B(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n307), .A2(new_n315), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT31), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n248), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n261), .A2(new_n310), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT28), .B1(new_n325), .B2(new_n304), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n292), .A2(new_n304), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n328), .A2(new_n306), .A3(new_n261), .A4(new_n287), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n255), .A2(new_n258), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n256), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n329), .A2(new_n330), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n327), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n321), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n309), .A2(new_n314), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n340), .A2(new_n334), .B1(new_n329), .B2(new_n330), .ZN(new_n341));
  INV_X1    g155(.A(new_n321), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n323), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n334), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n329), .A2(new_n330), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n324), .A2(new_n339), .A3(new_n343), .A4(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT32), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT32), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n348), .A2(new_n352), .A3(new_n349), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n335), .A2(new_n334), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n345), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n326), .B1(new_n356), .B2(KEYINPUT28), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT73), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n342), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT73), .B1(new_n338), .B2(new_n321), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n341), .A2(new_n342), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(KEYINPUT29), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n308), .A2(new_n334), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n345), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n326), .B1(new_n365), .B2(KEYINPUT28), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n342), .A2(KEYINPUT29), .ZN(new_n367));
  AOI21_X1  g181(.A(G902), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G472), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n247), .B1(new_n354), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n291), .A2(G125), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n297), .A2(new_n203), .A3(new_n298), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n373), .A2(KEYINPUT91), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(KEYINPUT91), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G224), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G953), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n376), .B(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT6), .ZN(new_n381));
  XOR2_X1   g195(.A(KEYINPUT89), .B(KEYINPUT5), .Z(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G113), .B1(new_n383), .B2(new_n249), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n253), .A2(new_n254), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n385), .A2(new_n258), .A3(new_n249), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n386), .B2(new_n383), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(G107), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT3), .A3(G104), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n391), .B2(G104), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(KEYINPUT82), .A3(G107), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n393), .A2(new_n394), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n389), .A2(G107), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n391), .A2(G104), .ZN(new_n400));
  OAI21_X1  g214(.A(G101), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n333), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n387), .A2(new_n403), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n391), .A2(KEYINPUT3), .A3(G104), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT3), .B1(new_n391), .B2(G104), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n396), .A2(new_n397), .ZN(new_n408));
  OAI21_X1  g222(.A(G101), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(KEYINPUT4), .A3(new_n398), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n411), .B(G101), .C1(new_n407), .C2(new_n408), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n410), .B(new_n412), .C1(new_n259), .C2(new_n260), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT88), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n334), .A2(KEYINPUT88), .A3(new_n412), .A4(new_n410), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n404), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G122), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n381), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n404), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n410), .A2(new_n412), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT88), .B1(new_n421), .B2(new_n334), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n413), .A2(new_n414), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n418), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n417), .A2(KEYINPUT90), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n419), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n418), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n417), .B2(KEYINPUT90), .ZN(new_n430));
  AOI211_X1 g244(.A(new_n425), .B(new_n404), .C1(new_n415), .C2(new_n416), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n430), .A2(new_n381), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n380), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G210), .B1(G237), .B2(G902), .ZN(new_n434));
  INV_X1    g248(.A(G902), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n418), .B(KEYINPUT8), .ZN(new_n436));
  INV_X1    g250(.A(new_n387), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n402), .B1(new_n437), .B2(new_n333), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n384), .B1(new_n386), .B2(KEYINPUT5), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(new_n403), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n436), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT7), .ZN(new_n442));
  OAI22_X1  g256(.A1(new_n372), .A2(new_n373), .B1(new_n442), .B2(new_n378), .ZN(new_n443));
  INV_X1    g257(.A(new_n378), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n376), .A2(KEYINPUT7), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n420), .B(new_n418), .C1(new_n422), .C2(new_n423), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n435), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n433), .A2(new_n434), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n434), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n447), .A2(KEYINPUT6), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n430), .B2(new_n431), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n424), .A2(new_n425), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n455), .A2(KEYINPUT6), .A3(new_n427), .A4(new_n429), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n379), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n452), .B1(new_n457), .B2(new_n449), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G214), .B1(G237), .B2(G902), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT92), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT92), .ZN(new_n462));
  INV_X1    g276(.A(new_n460), .ZN(new_n463));
  AOI211_X1 g277(.A(new_n462), .B(new_n463), .C1(new_n451), .C2(new_n458), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT9), .B(G234), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n226), .B1(new_n467), .B2(new_n435), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT94), .A2(KEYINPUT18), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n277), .A2(KEYINPUT93), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(G214), .A3(new_n317), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT93), .B(G143), .ZN(new_n473));
  INV_X1    g287(.A(G237), .ZN(new_n474));
  INV_X1    g288(.A(G953), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n474), .A2(new_n475), .A3(G214), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n472), .B(new_n269), .C1(new_n473), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT93), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G143), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n471), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n317), .A2(G214), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n269), .B1(new_n483), .B2(new_n472), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n470), .B1(new_n478), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n209), .A2(G146), .ZN(new_n486));
  INV_X1    g300(.A(new_n472), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n480), .A2(new_n471), .B1(new_n317), .B2(G214), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n215), .A2(new_n486), .B1(new_n489), .B2(new_n469), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n484), .A2(KEYINPUT17), .ZN(new_n492));
  OAI21_X1  g306(.A(G131), .B1(new_n487), .B2(new_n488), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n477), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n221), .B(new_n492), .C1(new_n494), .C2(KEYINPUT17), .ZN(new_n495));
  XNOR2_X1  g309(.A(G113), .B(G122), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(new_n389), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n491), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(new_n491), .B2(new_n495), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n435), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G475), .ZN(new_n501));
  NOR2_X1   g315(.A1(G475), .A2(G902), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT19), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n209), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n211), .A2(KEYINPUT19), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n493), .A2(new_n477), .B1(new_n506), .B2(new_n213), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n208), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n497), .B1(new_n491), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n502), .B1(new_n498), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(KEYINPUT20), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT20), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n491), .A2(new_n495), .A3(new_n497), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n485), .A2(new_n490), .B1(new_n208), .B2(new_n507), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n513), .B1(new_n514), .B2(new_n497), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n512), .B1(new_n515), .B2(new_n502), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n501), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT95), .ZN(new_n518));
  INV_X1    g332(.A(G952), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(G953), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n227), .B2(new_n474), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI211_X1 g336(.A(new_n435), .B(new_n475), .C1(G234), .C2(G237), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT21), .B(G898), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n501), .C1(new_n511), .C2(new_n516), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT97), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n251), .A2(G122), .A3(new_n252), .ZN(new_n530));
  INV_X1    g344(.A(G122), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G116), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n391), .ZN(new_n535));
  XNOR2_X1  g349(.A(G128), .B(G143), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT96), .B(G134), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n530), .A2(KEYINPUT14), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G107), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n530), .A2(KEYINPUT14), .A3(new_n533), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n535), .B(new_n538), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT13), .B1(new_n194), .B2(G143), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(new_n266), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(new_n536), .ZN(new_n545));
  INV_X1    g359(.A(new_n530), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n391), .B1(new_n546), .B2(new_n532), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n530), .A2(G107), .A3(new_n533), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n467), .A2(G217), .A3(new_n475), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n529), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n552), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n542), .A2(new_n549), .A3(KEYINPUT97), .A4(new_n551), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n435), .ZN(new_n557));
  INV_X1    g371(.A(G478), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(KEYINPUT15), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n559), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n556), .B2(new_n435), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n518), .A2(new_n526), .A3(new_n528), .A4(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G469), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(new_n435), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT83), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n398), .A2(new_n401), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(new_n568), .B2(new_n286), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n291), .A2(KEYINPUT83), .A3(new_n398), .A4(new_n401), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT10), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT84), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT84), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n569), .A2(new_n570), .A3(new_n574), .A4(new_n571), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n410), .A2(new_n299), .A3(new_n301), .A4(new_n412), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n402), .A2(KEYINPUT10), .A3(new_n291), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n576), .A2(new_n312), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(G110), .B(G140), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n475), .A2(G227), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n312), .B1(new_n576), .B2(new_n580), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT85), .ZN(new_n589));
  INV_X1    g403(.A(new_n312), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n590), .B(new_n579), .C1(new_n573), .C2(new_n575), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n568), .A2(new_n286), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n569), .A2(new_n570), .A3(new_n592), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n593), .A2(KEYINPUT12), .A3(new_n590), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT12), .B1(new_n593), .B2(new_n590), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n589), .B1(new_n591), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n595), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n593), .A2(KEYINPUT12), .A3(new_n590), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n581), .A2(new_n600), .A3(KEYINPUT85), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n588), .B1(new_n602), .B2(new_n584), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n566), .B1(new_n603), .B2(G469), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT87), .B1(new_n591), .B2(new_n584), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT87), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n581), .A2(new_n606), .A3(new_n585), .ZN(new_n607));
  OR3_X1    g421(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT86), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n600), .A2(KEYINPUT86), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n605), .A2(new_n607), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n584), .B1(new_n587), .B2(new_n591), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n565), .A3(new_n435), .ZN(new_n613));
  AOI211_X1 g427(.A(new_n468), .B(new_n564), .C1(new_n604), .C2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n371), .A2(new_n465), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  INV_X1    g430(.A(G472), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n348), .B2(new_n435), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n349), .B2(new_n348), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n468), .B1(new_n604), .B2(new_n613), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n241), .B1(new_n235), .B2(new_n236), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n621), .A2(new_n239), .B1(new_n244), .B2(new_n245), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n459), .A2(new_n460), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n556), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n550), .A2(new_n628), .A3(new_n551), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n542), .A2(new_n549), .B1(KEYINPUT98), .B2(new_n552), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT33), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n627), .A2(G478), .A3(new_n435), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n557), .A2(new_n558), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n528), .B2(new_n518), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n625), .A2(new_n525), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n624), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NAND2_X1  g455(.A1(new_n510), .A2(KEYINPUT20), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n515), .A2(new_n512), .A3(new_n502), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(KEYINPUT99), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(KEYINPUT99), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n646), .A2(new_n647), .B1(G475), .B2(new_n500), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n560), .A2(new_n562), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n463), .B1(new_n451), .B2(new_n458), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n651), .A3(new_n526), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n623), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT100), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT35), .B(G107), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  INV_X1    g470(.A(new_n618), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n230), .A2(KEYINPUT36), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT101), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n224), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n245), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n243), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n657), .A2(new_n658), .A3(new_n350), .A4(new_n663), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n248), .B(new_n323), .C1(new_n341), .C2(new_n342), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT72), .B1(new_n346), .B2(KEYINPUT31), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n321), .A2(new_n338), .B1(new_n322), .B2(new_n323), .ZN(new_n668));
  AOI21_X1  g482(.A(G902), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n350), .B(new_n663), .C1(new_n669), .C2(new_n617), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT102), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n465), .A2(new_n614), .A3(new_n664), .A4(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  AND3_X1   g488(.A1(new_n348), .A2(new_n352), .A3(new_n349), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n352), .B1(new_n348), .B2(new_n349), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n370), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n523), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n521), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n648), .A2(new_n649), .A3(new_n680), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n243), .A2(new_n662), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n677), .A2(new_n683), .A3(new_n651), .A4(new_n620), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XNOR2_X1  g499(.A(new_n680), .B(KEYINPUT39), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n620), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT40), .ZN(new_n688));
  INV_X1    g502(.A(new_n341), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n342), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n690), .B(new_n435), .C1(new_n342), .C2(new_n365), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G472), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n675), .B2(new_n676), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT38), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n459), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n518), .A2(new_n528), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n682), .A2(new_n460), .A3(new_n697), .A4(new_n649), .ZN(new_n698));
  NOR4_X1   g512(.A1(new_n688), .A2(new_n694), .A3(new_n696), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n277), .ZN(G45));
  AND3_X1   g514(.A1(new_n636), .A2(new_n663), .A3(new_n680), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n677), .A2(new_n651), .A3(new_n620), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  NAND2_X1  g517(.A1(new_n612), .A2(new_n435), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  INV_X1    g519(.A(new_n468), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n613), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT103), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n565), .B1(new_n612), .B2(new_n435), .ZN(new_n709));
  AOI211_X1 g523(.A(G469), .B(G902), .C1(new_n610), .C2(new_n611), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n709), .A2(new_n710), .A3(new_n468), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n371), .A2(new_n638), .A3(new_n708), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n371), .A2(new_n708), .A3(new_n713), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n717), .B1(new_n718), .B2(new_n652), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n713), .A2(new_n708), .ZN(new_n720));
  INV_X1    g534(.A(new_n652), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(KEYINPUT104), .A3(new_n371), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G116), .ZN(G18));
  NOR2_X1   g538(.A1(new_n682), .A2(new_n564), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n677), .A2(new_n651), .A3(new_n711), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  NOR2_X1   g541(.A1(new_n366), .A2(new_n342), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n346), .A2(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n343), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n349), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n622), .B(new_n731), .C1(new_n669), .C2(new_n617), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n657), .A2(KEYINPUT105), .A3(new_n622), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n528), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n527), .B1(new_n644), .B2(new_n501), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n649), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n625), .A2(new_n525), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n736), .A2(new_n708), .A3(new_n713), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT106), .B(G122), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G24));
  INV_X1    g557(.A(new_n731), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n618), .A2(new_n682), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n680), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n637), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n745), .A2(new_n711), .A3(new_n747), .A4(new_n651), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  NOR2_X1   g563(.A1(new_n468), .A2(new_n463), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n451), .A2(new_n458), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n603), .A2(G469), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT107), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n585), .B1(new_n597), .B2(new_n601), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n754), .A2(KEYINPUT107), .A3(new_n588), .A4(new_n565), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n710), .A2(new_n566), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n371), .A2(new_n747), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n371), .A2(KEYINPUT42), .A3(new_n747), .A4(new_n759), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  XNOR2_X1  g579(.A(new_n681), .B(KEYINPUT108), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n371), .A3(new_n759), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  NOR3_X1   g582(.A1(new_n591), .A2(new_n596), .A3(new_n589), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT85), .B1(new_n581), .B2(new_n600), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n584), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n588), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT109), .B1(new_n773), .B2(new_n565), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n775), .B(G469), .C1(new_n603), .C2(KEYINPUT45), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n603), .A2(KEYINPUT45), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n566), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n566), .A2(new_n781), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n710), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n706), .A3(new_n686), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n451), .A2(new_n458), .A3(new_n460), .ZN(new_n788));
  INV_X1    g602(.A(new_n619), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n518), .A2(new_n634), .A3(new_n528), .ZN(new_n790));
  NOR2_X1   g604(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n791), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n789), .B(new_n663), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT44), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n788), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n787), .B(new_n798), .C1(new_n797), .C2(new_n796), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  NAND2_X1  g614(.A1(new_n778), .A2(new_n783), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n613), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT46), .B1(new_n778), .B2(new_n779), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n706), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT47), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g622(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n785), .B2(new_n706), .ZN(new_n810));
  INV_X1    g624(.A(new_n788), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n747), .A2(new_n811), .A3(new_n247), .ZN(new_n812));
  OR4_X1    g626(.A1(new_n677), .A2(new_n808), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  NAND3_X1  g628(.A1(new_n741), .A2(new_n714), .A3(new_n726), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n719), .B2(new_n722), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n625), .A2(new_n462), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n651), .A2(KEYINPUT92), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n614), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n677), .A2(new_n622), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n697), .A2(new_n649), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n634), .B1(new_n518), .B2(new_n528), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n822), .A2(new_n525), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n818), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  OAI22_X1  g639(.A1(new_n820), .A2(new_n821), .B1(new_n825), .B2(new_n623), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n465), .A2(new_n614), .A3(new_n664), .A4(new_n671), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n817), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n624), .A2(new_n465), .A3(new_n824), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n615), .A3(KEYINPUT113), .A4(new_n672), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT107), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n603), .B2(G469), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n613), .B(new_n779), .C1(new_n834), .C2(new_n755), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n663), .A2(new_n468), .A3(new_n746), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n836), .B1(new_n835), .B2(new_n837), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n463), .B(new_n739), .C1(new_n458), .C2(new_n451), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n693), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n684), .A2(new_n702), .A3(new_n748), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n832), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n835), .A2(new_n837), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT115), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n693), .A3(new_n847), .A4(new_n840), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n620), .A2(new_n651), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n849), .B(new_n677), .C1(new_n683), .C2(new_n701), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n848), .A2(KEYINPUT52), .A3(new_n850), .A4(new_n748), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n844), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n560), .A2(new_n562), .A3(new_n746), .ZN(new_n853));
  INV_X1    g667(.A(new_n647), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n853), .B(new_n501), .C1(new_n854), .C2(new_n645), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT114), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n663), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n855), .A2(KEYINPUT114), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n857), .A2(new_n788), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n677), .A3(new_n620), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n759), .A2(new_n747), .A3(new_n745), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n767), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n763), .B2(new_n762), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n816), .A2(new_n831), .A3(new_n852), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT54), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n816), .A2(new_n831), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT53), .A3(new_n852), .A4(new_n863), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n864), .A2(new_n865), .ZN(new_n871));
  XOR2_X1   g685(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n522), .B1(new_n793), .B2(new_n795), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n734), .B2(new_n735), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n651), .A3(new_n711), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n707), .A2(new_n788), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n247), .A2(new_n521), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n694), .A3(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n876), .B(new_n520), .C1(new_n637), .C2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n795), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n521), .B1(new_n881), .B2(new_n792), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n877), .A2(KEYINPUT118), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT118), .B1(new_n877), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n885), .A2(KEYINPUT48), .A3(new_n821), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT48), .B1(new_n885), .B2(new_n821), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n880), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n745), .B1(new_n883), .B2(new_n884), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n635), .A2(new_n528), .A3(new_n518), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n879), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n618), .A2(new_n744), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT105), .B1(new_n892), .B2(new_n622), .ZN(new_n893));
  NOR4_X1   g707(.A1(new_n618), .A2(new_n744), .A3(new_n247), .A4(new_n733), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n882), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n696), .A2(new_n463), .A3(new_n711), .ZN(new_n896));
  NOR2_X1   g710(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n897), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n459), .A2(new_n695), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT38), .B1(new_n451), .B2(new_n458), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n463), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n707), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n900), .B1(new_n904), .B2(new_n875), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n889), .B(new_n891), .C1(new_n898), .C2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n705), .A2(new_n613), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n706), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n808), .B2(new_n810), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n895), .A2(new_n788), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n888), .B1(new_n912), .B2(KEYINPUT51), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n895), .A2(new_n896), .B1(new_n899), .B2(new_n897), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n904), .A2(new_n875), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n897), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n916), .A2(KEYINPUT51), .A3(new_n889), .A4(new_n891), .ZN(new_n917));
  INV_X1    g731(.A(new_n911), .ZN(new_n918));
  INV_X1    g732(.A(new_n809), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n804), .A2(new_n919), .ZN(new_n920));
  OAI221_X1 g734(.A(new_n706), .B1(new_n805), .B2(new_n806), .C1(new_n802), .C2(new_n803), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n908), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n918), .B1(new_n922), .B2(KEYINPUT119), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n910), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n917), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n913), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n868), .A2(new_n873), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n519), .A2(new_n475), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT120), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n907), .B(KEYINPUT49), .Z(new_n932));
  INV_X1    g746(.A(new_n790), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n622), .A3(new_n750), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT112), .Z(new_n935));
  NAND4_X1  g749(.A1(new_n932), .A2(new_n694), .A3(new_n696), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT121), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n931), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(G75));
  AOI21_X1  g755(.A(new_n435), .B1(new_n870), .B2(new_n871), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(G210), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT56), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n428), .A2(new_n432), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n379), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n433), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT55), .Z(new_n948));
  AND3_X1   g762(.A1(new_n943), .A2(new_n944), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n943), .B2(new_n944), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n475), .A2(G952), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(G51));
  INV_X1    g766(.A(new_n778), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n942), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT123), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n566), .B(KEYINPUT122), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT57), .Z(new_n957));
  INV_X1    g771(.A(new_n873), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n872), .B1(new_n870), .B2(new_n871), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n612), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n951), .B1(new_n955), .B2(new_n961), .ZN(G54));
  INV_X1    g776(.A(new_n951), .ZN(new_n963));
  NAND2_X1  g777(.A1(KEYINPUT58), .A2(G475), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT124), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n942), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n515), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n967), .B2(new_n966), .ZN(G60));
  AND2_X1   g783(.A1(new_n627), .A2(new_n631), .ZN(new_n970));
  NAND2_X1  g784(.A1(G478), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT59), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n970), .B(new_n972), .C1(new_n958), .C2(new_n959), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n963), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n868), .A2(new_n873), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n975), .B2(new_n972), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n974), .A2(new_n976), .ZN(G63));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT60), .Z(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n866), .B2(new_n867), .ZN(new_n980));
  INV_X1    g794(.A(new_n244), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n661), .B(new_n979), .C1(new_n866), .C2(new_n867), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n982), .A2(new_n963), .A3(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT61), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(G66));
  NOR3_X1   g800(.A1(new_n524), .A2(new_n377), .A3(new_n475), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n869), .B2(new_n475), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n945), .B1(G898), .B2(new_n475), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(G69));
  NAND2_X1  g804(.A1(G900), .A2(G953), .ZN(new_n991));
  AND4_X1   g805(.A1(new_n748), .A2(new_n764), .A3(new_n767), .A4(new_n850), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n787), .A2(new_n371), .A3(new_n840), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n813), .A2(new_n992), .A3(new_n799), .A4(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n991), .B1(new_n994), .B2(G953), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n340), .B(KEYINPUT125), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(new_n506), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n699), .A2(new_n843), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT62), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n822), .A2(new_n823), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT126), .Z(new_n1001));
  OR4_X1    g815(.A1(new_n821), .A2(new_n1001), .A3(new_n687), .A4(new_n788), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n999), .A2(new_n799), .A3(new_n813), .A4(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n997), .A2(G953), .ZN(new_n1004));
  AOI22_X1  g818(.A1(new_n995), .A2(new_n997), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n475), .B1(G227), .B2(G900), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(G72));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1003), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(new_n869), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n963), .B1(new_n1012), .B2(new_n690), .ZN(new_n1013));
  INV_X1    g827(.A(new_n869), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n994), .A2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g829(.A(new_n342), .B(new_n689), .C1(new_n1015), .C2(new_n1009), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n346), .A2(KEYINPUT127), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(new_n361), .ZN(new_n1018));
  AOI211_X1 g832(.A(new_n1010), .B(new_n1018), .C1(new_n870), .C2(new_n871), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n1013), .A2(new_n1016), .A3(new_n1019), .ZN(G57));
endmodule


