//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n440, new_n442, new_n444, new_n449, new_n450, new_n451, new_n454,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(new_n440));
  INV_X1    g015(.A(new_n440), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT66), .B(G108), .Z(new_n442));
  INV_X1    g017(.A(new_n442), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT69), .ZN(new_n450));
  AND2_X1   g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(G223));
  NAND2_X1  g027(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g028(.A1(new_n451), .A2(G2106), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT70), .Z(G217));
  OR4_X1    g030(.A1(G221), .A2(G218), .A3(G219), .A4(G220), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT2), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n442), .A2(G69), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n440), .A2(G120), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(new_n460), .ZN(G261));
  INV_X1    g036(.A(G261), .ZN(G325));
  INV_X1    g037(.A(new_n457), .ZN(new_n463));
  OAI21_X1  g038(.A(G567), .B1(new_n458), .B2(new_n459), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G2106), .B1(KEYINPUT71), .B2(new_n465), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n465), .A2(KEYINPUT71), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(G319));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(G137), .B(new_n477), .C1(new_n470), .C2(new_n471), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT72), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n481), .A2(KEYINPUT72), .A3(G137), .A4(new_n477), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n477), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G101), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n476), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  OAI21_X1  g062(.A(KEYINPUT75), .B1(G100), .B2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n477), .A2(G112), .ZN(new_n490));
  NOR3_X1   g065(.A1(KEYINPUT75), .A2(G100), .A3(G2105), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n472), .B2(new_n477), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n481), .A2(KEYINPUT74), .A3(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n496), .A2(G124), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n472), .A2(G2105), .ZN(new_n498));
  XNOR2_X1  g073(.A(new_n498), .B(KEYINPUT73), .ZN(new_n499));
  AOI211_X1 g074(.A(new_n492), .B(new_n497), .C1(G136), .C2(new_n499), .ZN(G162));
  OAI211_X1 g075(.A(G138), .B(new_n477), .C1(new_n470), .C2(new_n471), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n481), .A2(new_n503), .A3(G138), .A4(new_n477), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n484), .A2(G102), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n481), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(new_n477), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n506), .A2(new_n509), .ZN(G164));
  AND2_X1   g085(.A1(G75), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT77), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT77), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(G543), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n513), .A2(new_n516), .B1(KEYINPUT5), .B2(new_n512), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n511), .B1(new_n517), .B2(G62), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(KEYINPUT6), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G651), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n517), .A2(G88), .A3(new_n524), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n521), .A2(new_n523), .A3(G50), .A4(G543), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT76), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n520), .A2(KEYINPUT78), .A3(new_n525), .A4(new_n528), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n528), .B(new_n525), .C1(new_n519), .C2(new_n518), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT78), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(new_n532), .ZN(G166));
  NAND2_X1  g108(.A1(G63), .A2(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n521), .A2(new_n523), .ZN(new_n535));
  INV_X1    g110(.A(G89), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT79), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n524), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n535), .A2(KEYINPUT79), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(G543), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G51), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n538), .B(new_n540), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(G168));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n517), .A2(new_n524), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n544), .A2(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n519), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n551), .A2(new_n553), .ZN(G171));
  INV_X1    g129(.A(G43), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n544), .A2(new_n555), .B1(new_n556), .B2(new_n550), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n519), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  NAND4_X1  g141(.A1(new_n542), .A2(G53), .A3(G543), .A4(new_n543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n513), .A2(new_n516), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g147(.A(KEYINPUT80), .B(G65), .Z(new_n573));
  OAI21_X1  g148(.A(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n550), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n574), .A2(G651), .B1(new_n575), .B2(G91), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n568), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  XNOR2_X1  g153(.A(new_n546), .B(KEYINPUT81), .ZN(G286));
  AND2_X1   g154(.A1(new_n529), .A2(new_n532), .ZN(G303));
  AND3_X1   g155(.A1(new_n542), .A2(G543), .A3(new_n543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G49), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n575), .A2(G87), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n572), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G48), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT82), .B1(new_n535), .B2(new_n589), .ZN(new_n590));
  OR3_X1    g165(.A1(new_n535), .A2(KEYINPUT82), .A3(new_n589), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n588), .A2(G651), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n575), .A2(G86), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n581), .A2(G47), .B1(new_n575), .B2(G85), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT83), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n519), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT84), .B(G66), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n517), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT85), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n603), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(G651), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n581), .A2(G54), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n517), .A2(G92), .A3(new_n524), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n609), .A2(KEYINPUT86), .A3(new_n610), .A4(new_n613), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n601), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n601), .B1(new_n618), .B2(G868), .ZN(G321));
  MUX2_X1   g195(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g196(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n618), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n618), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n498), .A2(G2104), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n499), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n496), .A2(G123), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(KEYINPUT87), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(KEYINPUT87), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n636), .B(new_n637), .C1(G111), .C2(new_n477), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n633), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n632), .A2(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(KEYINPUT89), .B(G2438), .Z(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT88), .B(KEYINPUT14), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT90), .B(G1341), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2443), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n657), .A2(G14), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT91), .Z(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT17), .Z(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n659), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n660), .ZN(new_n666));
  INV_X1    g241(.A(new_n662), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n663), .A3(new_n659), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n664), .A2(new_n659), .A3(new_n660), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2096), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(G2100), .Z(G227));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT92), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n674), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n683), .A2(new_n680), .A3(new_n678), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n678), .A2(new_n674), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n685), .A2(new_n682), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n681), .B(new_n684), .C1(new_n686), .C2(new_n680), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  NAND2_X1  g268(.A1(new_n499), .A2(G141), .ZN(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT26), .Z(new_n696));
  AOI22_X1  g271(.A1(new_n496), .A2(G129), .B1(G105), .B2(new_n484), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT98), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G29), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G29), .B2(G32), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT27), .B(G1996), .ZN(new_n706));
  OR2_X1    g281(.A1(KEYINPUT24), .A2(G34), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(KEYINPUT24), .A2(G34), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G160), .B2(new_n708), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n705), .A2(new_n706), .B1(G2084), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n484), .A2(G103), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT97), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n499), .A2(new_n717), .A3(G139), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n499), .B2(G139), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n715), .B1(new_n477), .B2(new_n716), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G33), .B(new_n720), .S(G29), .Z(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(G2072), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n712), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT99), .Z(new_n724));
  NAND2_X1  g299(.A1(G168), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G16), .B2(G21), .ZN(new_n726));
  INV_X1    g301(.A(G1966), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT100), .Z(new_n729));
  NOR2_X1   g304(.A1(new_n726), .A2(new_n727), .ZN(new_n730));
  AND2_X1   g305(.A1(KEYINPUT30), .A2(G28), .ZN(new_n731));
  NOR2_X1   g306(.A1(KEYINPUT30), .A2(G28), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n708), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n639), .B2(new_n708), .ZN(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  NOR2_X1   g310(.A1(G164), .A2(new_n708), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G27), .B2(new_n708), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT31), .B(G11), .ZN(new_n739));
  NOR2_X1   g314(.A1(G16), .A2(G19), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n560), .B2(G16), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G1341), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(G1341), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n738), .A2(new_n739), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  OAI22_X1  g319(.A1(new_n737), .A2(new_n735), .B1(G2084), .B2(new_n711), .ZN(new_n745));
  NOR4_X1   g320(.A1(new_n729), .A2(new_n730), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n708), .A2(G35), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G162), .B2(new_n708), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT29), .B(G2090), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT23), .ZN(new_n751));
  INV_X1    g326(.A(G16), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n751), .B(new_n753), .C1(G299), .C2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n751), .B2(new_n753), .ZN(new_n755));
  INV_X1    g330(.A(G1956), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n746), .A2(new_n750), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n752), .A2(G5), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G171), .B2(new_n752), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT101), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT28), .ZN(new_n762));
  INV_X1    g337(.A(G26), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(G29), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(G29), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n499), .A2(G140), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n496), .A2(G128), .ZN(new_n767));
  NOR2_X1   g342(.A1(G104), .A2(G2105), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(new_n477), .B2(G116), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n765), .B1(new_n770), .B2(G29), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(new_n762), .ZN(new_n772));
  AOI22_X1  g347(.A1(G1961), .A2(new_n761), .B1(new_n772), .B2(G2067), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n773), .B1(G1961), .B2(new_n761), .C1(new_n705), .C2(new_n706), .ZN(new_n774));
  NOR2_X1   g349(.A1(G4), .A2(G16), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n618), .B2(G16), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(G1348), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n776), .A2(G1348), .ZN(new_n778));
  OR3_X1    g353(.A1(new_n774), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n724), .A2(new_n758), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n752), .A2(G24), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n599), .B2(new_n752), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1986), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n752), .A2(G23), .ZN(new_n784));
  INV_X1    g359(.A(G288), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n752), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT33), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1976), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n752), .A2(G6), .ZN(new_n789));
  INV_X1    g364(.A(G305), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n752), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT32), .B(G1981), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G22), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G166), .B2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G1971), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n788), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n783), .B1(new_n799), .B2(KEYINPUT34), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n708), .A2(G25), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(new_n477), .B2(G107), .ZN(new_n802));
  INV_X1    g377(.A(G95), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n477), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n499), .B2(G131), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n496), .A2(G119), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n801), .B1(new_n808), .B2(new_n708), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT93), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT35), .B(G1991), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n800), .B(new_n812), .C1(KEYINPUT34), .C2(new_n799), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n772), .A2(G2067), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n813), .A2(new_n814), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n780), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  NAND2_X1  g394(.A1(new_n618), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n581), .A2(G55), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n575), .A2(G93), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n822), .B(new_n823), .C1(new_n519), .C2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n560), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT39), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n821), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(G860), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT102), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n825), .A2(G860), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT37), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(G145));
  XNOR2_X1  g408(.A(new_n702), .B(new_n770), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n720), .ZN(new_n835));
  NAND2_X1  g410(.A1(G114), .A2(G2104), .ZN(new_n836));
  INV_X1    g411(.A(G126), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n472), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n838), .A2(G2105), .B1(G102), .B2(new_n484), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT103), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT103), .B1(new_n502), .B2(new_n504), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n835), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n835), .A2(new_n842), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n499), .A2(G142), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n496), .A2(G130), .ZN(new_n847));
  NOR2_X1   g422(.A1(G106), .A2(G2105), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(new_n477), .B2(G118), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n630), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n639), .B(new_n486), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n808), .B(G162), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n845), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  INV_X1    g432(.A(new_n855), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n843), .A2(new_n844), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n825), .A2(G868), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n625), .B(new_n826), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n614), .B(G299), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT41), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n826), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n625), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n866), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(G166), .B(G288), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(G305), .ZN(new_n875));
  NOR2_X1   g450(.A1(G303), .A2(G288), .ZN(new_n876));
  NOR2_X1   g451(.A1(G166), .A2(new_n785), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n790), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n875), .A2(new_n599), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n599), .B1(new_n875), .B2(new_n878), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n880), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n875), .A2(new_n599), .A3(new_n878), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n873), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n879), .A2(new_n880), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n881), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n882), .B1(new_n879), .B2(new_n880), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n868), .A4(new_n872), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n891), .A3(KEYINPUT105), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n873), .B(new_n893), .C1(new_n883), .C2(new_n886), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G868), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n862), .B(new_n864), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n896), .B1(new_n892), .B2(new_n894), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT106), .B1(new_n898), .B2(new_n863), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(G295));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n863), .ZN(G331));
  NOR2_X1   g476(.A1(G171), .A2(new_n546), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(G286), .A2(G171), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n826), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n902), .B(KEYINPUT107), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n869), .A3(new_n905), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n909), .A3(new_n866), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n907), .A2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n911), .B2(new_n867), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n912), .A2(new_n888), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n857), .B1(new_n912), .B2(new_n888), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT108), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n916), .B(new_n857), .C1(new_n912), .C2(new_n888), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n913), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n913), .A2(new_n914), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT44), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OR3_X1    g497(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT43), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n918), .B2(new_n920), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(G397));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n505), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT103), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n509), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(G1384), .ZN(new_n932));
  XOR2_X1   g507(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(KEYINPUT110), .B(G40), .ZN(new_n935));
  AND4_X1   g510(.A1(new_n476), .A2(new_n483), .A3(new_n485), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT111), .ZN(new_n938));
  INV_X1    g513(.A(G1996), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT126), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n940), .B1(new_n941), .B2(KEYINPUT46), .ZN(new_n942));
  INV_X1    g517(.A(G2067), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n770), .B(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n938), .B1(new_n702), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT126), .B(KEYINPUT46), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n942), .B(new_n946), .C1(new_n940), .C2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n703), .A2(new_n939), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n702), .A2(G1996), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n944), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n808), .A2(new_n811), .ZN(new_n954));
  OAI22_X1  g529(.A1(new_n953), .A2(new_n954), .B1(G2067), .B2(new_n770), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n938), .ZN(new_n956));
  INV_X1    g531(.A(G1986), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n938), .A2(new_n957), .A3(new_n599), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT48), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n807), .B(new_n811), .Z(new_n960));
  OAI21_X1  g535(.A(new_n938), .B1(new_n953), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n950), .A2(new_n956), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n842), .A2(new_n936), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G8), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT52), .B1(G288), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n968), .B(new_n970), .C1(new_n969), .C2(G288), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT49), .ZN(new_n972));
  NOR2_X1   g547(.A1(G305), .A2(G1981), .ZN(new_n973));
  INV_X1    g548(.A(G1981), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT117), .B(G86), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n575), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n592), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n972), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n592), .A2(new_n976), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(G1981), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n980), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n981), .A3(new_n968), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n965), .B(G8), .C1(new_n969), .C2(G288), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n983), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT116), .B1(new_n983), .B2(KEYINPUT52), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n971), .B(new_n982), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n529), .A2(new_n532), .A3(G8), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(KEYINPUT115), .A3(new_n988), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n991), .B(new_n992), .C1(new_n988), .C2(new_n987), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n476), .A2(new_n483), .A3(new_n485), .A4(new_n935), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n964), .B1(new_n506), .B2(new_n509), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n842), .A2(new_n997), .A3(new_n964), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT113), .B(G2090), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n842), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1002));
  INV_X1    g577(.A(new_n933), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n995), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n936), .A3(new_n1004), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n1000), .A2(new_n1001), .B1(new_n1005), .B2(new_n797), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n967), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n986), .B1(new_n993), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n992), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT115), .B1(new_n987), .B2(new_n988), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n987), .A2(new_n988), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1384), .B1(new_n839), .B2(new_n505), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n997), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n936), .B(new_n1015), .C1(new_n932), .C2(new_n997), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1017), .A2(new_n999), .B1(new_n797), .B2(new_n1005), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1013), .B1(new_n1018), .B2(new_n967), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1009), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n1005), .B2(G2078), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n996), .A2(new_n998), .ZN(new_n1024));
  INV_X1    g599(.A(G1961), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n931), .B2(G1384), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n994), .B1(new_n1014), .B2(new_n933), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1029), .A2(KEYINPUT53), .A3(new_n735), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G171), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n934), .A2(new_n1022), .A3(G2078), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(G40), .A3(G160), .A4(new_n1002), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(new_n1027), .A3(G301), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1021), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1020), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1023), .A2(G301), .A3(new_n1026), .A4(new_n1031), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT54), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1035), .A2(new_n1027), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(G171), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n546), .A2(G8), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT45), .B1(new_n842), .B2(new_n964), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n964), .B(new_n933), .C1(new_n506), .C2(new_n509), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n936), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n727), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G2084), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n996), .A2(new_n998), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1043), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n996), .A2(new_n998), .A3(new_n1048), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1966), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1052), .B1(new_n1055), .B2(new_n1043), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n967), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1043), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1057), .A2(KEYINPUT51), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1051), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT122), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1055), .A2(new_n1052), .A3(new_n1043), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT51), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(KEYINPUT122), .A3(new_n1051), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1042), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n964), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n994), .B1(new_n1069), .B2(KEYINPUT50), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1956), .B1(new_n1070), .B2(new_n1015), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n568), .A2(KEYINPUT57), .A3(new_n576), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n568), .B2(new_n576), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1002), .A2(new_n936), .A3(new_n1004), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1071), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1073), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n568), .A2(KEYINPUT57), .A3(new_n576), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1016), .A2(new_n756), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(new_n1076), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1068), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n616), .A2(new_n617), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n966), .A2(new_n943), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1024), .A2(new_n649), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1074), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1082), .A2(new_n1081), .A3(new_n1076), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(KEYINPUT61), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n618), .A2(new_n1094), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1084), .A2(new_n1090), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1002), .A2(new_n936), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(KEYINPUT120), .A3(new_n939), .A4(new_n1004), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1005), .B2(G1996), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n965), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n560), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1104), .B1(new_n1103), .B2(new_n560), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT59), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1103), .A2(new_n560), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n1105), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1096), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1091), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1038), .B(new_n1067), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n986), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1008), .A2(new_n993), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1055), .A2(G286), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1117), .A2(new_n1019), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1009), .A2(KEYINPUT119), .A3(new_n1019), .A4(new_n1119), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1008), .A2(new_n993), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1009), .A2(KEYINPUT63), .A3(new_n1119), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1118), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n982), .A2(new_n969), .A3(new_n785), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n973), .B(KEYINPUT118), .Z(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1129), .A2(new_n1117), .B1(new_n968), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1116), .A2(new_n1128), .A3(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1009), .A2(G171), .A3(new_n1019), .A4(new_n1032), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT122), .B1(new_n1065), .B2(new_n1051), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1061), .B(new_n1050), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1135), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT124), .B1(new_n1141), .B2(KEYINPUT62), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1143), .B(new_n1139), .C1(new_n1062), .C2(new_n1066), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1140), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT125), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1140), .B(new_n1147), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1134), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n938), .A2(G1986), .A3(G290), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n958), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT112), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n961), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n963), .B1(new_n1149), .B2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g729(.A1(G229), .A2(new_n468), .ZN(new_n1156));
  AOI21_X1  g730(.A(G227), .B1(new_n657), .B2(G14), .ZN(new_n1157));
  NAND4_X1  g731(.A1(new_n924), .A2(new_n860), .A3(new_n1156), .A4(new_n1157), .ZN(G225));
  INV_X1    g732(.A(G225), .ZN(G308));
endmodule


