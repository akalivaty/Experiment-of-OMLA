

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(G1384), .A2(G164), .ZN(n764) );
  INV_X1 U554 ( .A(n733), .ZN(n710) );
  INV_X1 U555 ( .A(n932), .ZN(n747) );
  AND2_X1 U556 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U557 ( .A1(G543), .A2(G651), .ZN(n640) );
  INV_X1 U558 ( .A(G2104), .ZN(n520) );
  INV_X1 U559 ( .A(G2105), .ZN(n525) );
  NOR2_X1 U560 ( .A1(n520), .A2(n525), .ZN(n867) );
  NAND2_X1 U561 ( .A1(n867), .A2(G113), .ZN(n523) );
  NOR2_X4 U562 ( .A1(G2105), .A2(n520), .ZN(n874) );
  NAND2_X1 U563 ( .A1(G101), .A2(n874), .ZN(n521) );
  XOR2_X1 U564 ( .A(KEYINPUT23), .B(n521), .Z(n522) );
  NAND2_X1 U565 ( .A1(n523), .A2(n522), .ZN(n529) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XOR2_X2 U567 ( .A(KEYINPUT17), .B(n524), .Z(n865) );
  NAND2_X1 U568 ( .A1(G137), .A2(n865), .ZN(n527) );
  NOR2_X1 U569 ( .A1(n525), .A2(G2104), .ZN(n868) );
  NAND2_X1 U570 ( .A1(G125), .A2(n868), .ZN(n526) );
  NAND2_X1 U571 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U572 ( .A1(n529), .A2(n528), .ZN(G160) );
  AND2_X1 U573 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U574 ( .A(G860), .ZN(n591) );
  NAND2_X1 U575 ( .A1(n640), .A2(G81), .ZN(n530) );
  XNOR2_X1 U576 ( .A(n530), .B(KEYINPUT12), .ZN(n532) );
  XOR2_X1 U577 ( .A(G543), .B(KEYINPUT0), .Z(n630) );
  INV_X1 U578 ( .A(G651), .ZN(n536) );
  NOR2_X1 U579 ( .A1(n630), .A2(n536), .ZN(n642) );
  NAND2_X1 U580 ( .A1(G68), .A2(n642), .ZN(n531) );
  NAND2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U582 ( .A(n533), .B(KEYINPUT13), .ZN(n535) );
  NOR2_X1 U583 ( .A1(G651), .A2(n630), .ZN(n643) );
  NAND2_X1 U584 ( .A1(G43), .A2(n643), .ZN(n534) );
  NAND2_X1 U585 ( .A1(n535), .A2(n534), .ZN(n540) );
  NOR2_X1 U586 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n537), .Z(n646) );
  NAND2_X1 U588 ( .A1(n646), .A2(G56), .ZN(n538) );
  XOR2_X1 U589 ( .A(KEYINPUT14), .B(n538), .Z(n539) );
  NOR2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U591 ( .A(KEYINPUT72), .B(n541), .Z(n927) );
  OR2_X1 U592 ( .A1(n591), .A2(n927), .ZN(G153) );
  INV_X1 U593 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U594 ( .A(KEYINPUT6), .B(KEYINPUT74), .ZN(n545) );
  NAND2_X1 U595 ( .A1(G51), .A2(n643), .ZN(n543) );
  NAND2_X1 U596 ( .A1(G63), .A2(n646), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U598 ( .A(n545), .B(n544), .ZN(n552) );
  NAND2_X1 U599 ( .A1(n640), .A2(G89), .ZN(n546) );
  XNOR2_X1 U600 ( .A(n546), .B(KEYINPUT4), .ZN(n548) );
  NAND2_X1 U601 ( .A1(G76), .A2(n642), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U603 ( .A(KEYINPUT5), .B(n549), .ZN(n550) );
  XNOR2_X1 U604 ( .A(KEYINPUT73), .B(n550), .ZN(n551) );
  NOR2_X1 U605 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U606 ( .A(KEYINPUT7), .B(n553), .Z(G168) );
  XOR2_X1 U607 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U608 ( .A1(G126), .A2(n868), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G138), .A2(n865), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U611 ( .A1(G114), .A2(n867), .ZN(n557) );
  NAND2_X1 U612 ( .A1(G102), .A2(n874), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U615 ( .A(n560), .B(KEYINPUT88), .ZN(G164) );
  NAND2_X1 U616 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U617 ( .A(n561), .B(KEYINPUT10), .ZN(n562) );
  XNOR2_X1 U618 ( .A(KEYINPUT70), .B(n562), .ZN(G223) );
  INV_X1 U619 ( .A(G223), .ZN(n821) );
  NAND2_X1 U620 ( .A1(n821), .A2(G567), .ZN(n563) );
  XNOR2_X1 U621 ( .A(n563), .B(KEYINPUT71), .ZN(n564) );
  XNOR2_X1 U622 ( .A(KEYINPUT11), .B(n564), .ZN(G234) );
  NAND2_X1 U623 ( .A1(G52), .A2(n643), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G64), .A2(n646), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n571) );
  NAND2_X1 U626 ( .A1(G90), .A2(n640), .ZN(n568) );
  NAND2_X1 U627 ( .A1(G77), .A2(n642), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U629 ( .A(KEYINPUT9), .B(n569), .Z(n570) );
  NOR2_X1 U630 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U631 ( .A(KEYINPUT68), .B(n572), .ZN(G171) );
  INV_X1 U632 ( .A(G171), .ZN(G301) );
  NAND2_X1 U633 ( .A1(G301), .A2(G868), .ZN(n581) );
  NAND2_X1 U634 ( .A1(G92), .A2(n640), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G79), .A2(n642), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G54), .A2(n643), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G66), .A2(n646), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT15), .B(n579), .Z(n922) );
  OR2_X1 U642 ( .A1(n922), .A2(G868), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U644 ( .A1(G53), .A2(n643), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G65), .A2(n646), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT69), .B(n584), .ZN(n588) );
  NAND2_X1 U648 ( .A1(G91), .A2(n640), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G78), .A2(n642), .ZN(n585) );
  AND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(G299) );
  INV_X1 U652 ( .A(G868), .ZN(n660) );
  NOR2_X1 U653 ( .A1(G286), .A2(n660), .ZN(n590) );
  NOR2_X1 U654 ( .A1(G868), .A2(G299), .ZN(n589) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(G297) );
  NAND2_X1 U656 ( .A1(n591), .A2(G559), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n592), .A2(n922), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n593), .B(KEYINPUT16), .ZN(n594) );
  XOR2_X1 U659 ( .A(KEYINPUT75), .B(n594), .Z(G148) );
  NAND2_X1 U660 ( .A1(n922), .A2(G868), .ZN(n595) );
  XNOR2_X1 U661 ( .A(KEYINPUT76), .B(n595), .ZN(n596) );
  NOR2_X1 U662 ( .A1(G559), .A2(n596), .ZN(n598) );
  NOR2_X1 U663 ( .A1(n927), .A2(G868), .ZN(n597) );
  NOR2_X1 U664 ( .A1(n598), .A2(n597), .ZN(G282) );
  NAND2_X1 U665 ( .A1(G111), .A2(n867), .ZN(n600) );
  NAND2_X1 U666 ( .A1(G99), .A2(n874), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U668 ( .A(KEYINPUT78), .B(n601), .ZN(n607) );
  NAND2_X1 U669 ( .A1(G123), .A2(n868), .ZN(n602) );
  XOR2_X1 U670 ( .A(KEYINPUT77), .B(n602), .Z(n603) );
  XNOR2_X1 U671 ( .A(n603), .B(KEYINPUT18), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G135), .A2(n865), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U674 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U675 ( .A(KEYINPUT79), .B(n608), .Z(n988) );
  XNOR2_X1 U676 ( .A(n988), .B(G2096), .ZN(n610) );
  INV_X1 U677 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U679 ( .A1(G85), .A2(n640), .ZN(n612) );
  NAND2_X1 U680 ( .A1(G72), .A2(n642), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U682 ( .A(KEYINPUT66), .B(n613), .ZN(n616) );
  NAND2_X1 U683 ( .A1(G47), .A2(n643), .ZN(n614) );
  XNOR2_X1 U684 ( .A(KEYINPUT67), .B(n614), .ZN(n615) );
  NOR2_X1 U685 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n646), .A2(G60), .ZN(n617) );
  NAND2_X1 U687 ( .A1(n618), .A2(n617), .ZN(G290) );
  NAND2_X1 U688 ( .A1(G73), .A2(n642), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n619), .B(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U690 ( .A1(G48), .A2(n643), .ZN(n621) );
  NAND2_X1 U691 ( .A1(G61), .A2(n646), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U693 ( .A1(G86), .A2(n640), .ZN(n622) );
  XNOR2_X1 U694 ( .A(KEYINPUT83), .B(n622), .ZN(n623) );
  NOR2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n626), .A2(n625), .ZN(G305) );
  NAND2_X1 U697 ( .A1(G49), .A2(n643), .ZN(n628) );
  NAND2_X1 U698 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U700 ( .A1(n646), .A2(n629), .ZN(n632) );
  NAND2_X1 U701 ( .A1(n630), .A2(G87), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U703 ( .A1(G50), .A2(n643), .ZN(n634) );
  NAND2_X1 U704 ( .A1(G62), .A2(n646), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U706 ( .A(KEYINPUT84), .B(n635), .Z(n639) );
  NAND2_X1 U707 ( .A1(G88), .A2(n640), .ZN(n637) );
  NAND2_X1 U708 ( .A1(G75), .A2(n642), .ZN(n636) );
  AND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n639), .A2(n638), .ZN(G303) );
  INV_X1 U711 ( .A(G303), .ZN(G166) );
  NAND2_X1 U712 ( .A1(n922), .A2(G559), .ZN(n912) );
  NAND2_X1 U713 ( .A1(G93), .A2(n640), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n641), .B(KEYINPUT80), .ZN(n651) );
  NAND2_X1 U715 ( .A1(G80), .A2(n642), .ZN(n645) );
  NAND2_X1 U716 ( .A1(G55), .A2(n643), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U718 ( .A1(G67), .A2(n646), .ZN(n647) );
  XNOR2_X1 U719 ( .A(KEYINPUT81), .B(n647), .ZN(n648) );
  NOR2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U722 ( .A(KEYINPUT82), .B(n652), .ZN(n915) );
  XNOR2_X1 U723 ( .A(KEYINPUT19), .B(G305), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n653), .B(G288), .ZN(n654) );
  XNOR2_X1 U725 ( .A(G290), .B(n654), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n927), .B(G166), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n915), .B(n657), .ZN(n658) );
  XNOR2_X1 U729 ( .A(n658), .B(G299), .ZN(n894) );
  XNOR2_X1 U730 ( .A(n912), .B(n894), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n659), .A2(G868), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n915), .A2(n660), .ZN(n661) );
  NAND2_X1 U733 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U734 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XOR2_X1 U735 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U736 ( .A1(G2090), .A2(n664), .ZN(n666) );
  XOR2_X1 U737 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n665) );
  XNOR2_X1 U738 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U739 ( .A1(n667), .A2(G2072), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n668), .B(KEYINPUT86), .ZN(G158) );
  XNOR2_X1 U741 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U742 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n670) );
  NAND2_X1 U743 ( .A1(G132), .A2(G82), .ZN(n669) );
  XNOR2_X1 U744 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X1 U745 ( .A1(n671), .A2(G218), .ZN(n672) );
  NAND2_X1 U746 ( .A1(G96), .A2(n672), .ZN(n916) );
  NAND2_X1 U747 ( .A1(n916), .A2(G2106), .ZN(n676) );
  NAND2_X1 U748 ( .A1(G69), .A2(G120), .ZN(n673) );
  NOR2_X1 U749 ( .A1(G237), .A2(n673), .ZN(n674) );
  NAND2_X1 U750 ( .A1(G108), .A2(n674), .ZN(n917) );
  NAND2_X1 U751 ( .A1(n917), .A2(G567), .ZN(n675) );
  NAND2_X1 U752 ( .A1(n676), .A2(n675), .ZN(n827) );
  NAND2_X1 U753 ( .A1(G661), .A2(G483), .ZN(n677) );
  NOR2_X1 U754 ( .A1(n827), .A2(n677), .ZN(n826) );
  NAND2_X1 U755 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U756 ( .A1(G40), .A2(G160), .ZN(n678) );
  XOR2_X1 U757 ( .A(n678), .B(KEYINPUT89), .Z(n763) );
  INV_X1 U758 ( .A(n763), .ZN(n679) );
  NAND2_X2 U759 ( .A1(n764), .A2(n679), .ZN(n733) );
  NAND2_X1 U760 ( .A1(G8), .A2(n733), .ZN(n811) );
  NOR2_X1 U761 ( .A1(G1976), .A2(G288), .ZN(n930) );
  NAND2_X1 U762 ( .A1(n930), .A2(KEYINPUT33), .ZN(n680) );
  NOR2_X1 U763 ( .A1(n811), .A2(n680), .ZN(n752) );
  NOR2_X1 U764 ( .A1(G2084), .A2(n733), .ZN(n715) );
  NAND2_X1 U765 ( .A1(G8), .A2(n715), .ZN(n730) );
  NOR2_X1 U766 ( .A1(G1966), .A2(n811), .ZN(n681) );
  XOR2_X1 U767 ( .A(KEYINPUT93), .B(n681), .Z(n728) );
  AND2_X1 U768 ( .A1(n710), .A2(G1996), .ZN(n683) );
  XOR2_X1 U769 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n682) );
  XNOR2_X1 U770 ( .A(n683), .B(n682), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n733), .A2(G1341), .ZN(n684) );
  NAND2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U773 ( .A1(n927), .A2(n686), .ZN(n687) );
  XOR2_X1 U774 ( .A(KEYINPUT65), .B(n687), .Z(n689) );
  NOR2_X1 U775 ( .A1(n689), .A2(n922), .ZN(n688) );
  XNOR2_X1 U776 ( .A(n688), .B(KEYINPUT95), .ZN(n701) );
  NAND2_X1 U777 ( .A1(n689), .A2(n922), .ZN(n694) );
  NAND2_X1 U778 ( .A1(G1348), .A2(n733), .ZN(n691) );
  NAND2_X1 U779 ( .A1(G2067), .A2(n710), .ZN(n690) );
  NAND2_X1 U780 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U781 ( .A(KEYINPUT94), .B(n692), .ZN(n693) );
  NAND2_X1 U782 ( .A1(n694), .A2(n693), .ZN(n699) );
  NAND2_X1 U783 ( .A1(n710), .A2(G2072), .ZN(n695) );
  XOR2_X1 U784 ( .A(KEYINPUT27), .B(n695), .Z(n697) );
  NAND2_X1 U785 ( .A1(G1956), .A2(n733), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n697), .A2(n696), .ZN(n703) );
  NAND2_X1 U787 ( .A1(G299), .A2(n703), .ZN(n698) );
  XNOR2_X1 U788 ( .A(n698), .B(KEYINPUT28), .ZN(n702) );
  AND2_X1 U789 ( .A1(n699), .A2(n702), .ZN(n700) );
  NAND2_X1 U790 ( .A1(n701), .A2(n700), .ZN(n708) );
  INV_X1 U791 ( .A(n702), .ZN(n706) );
  NOR2_X1 U792 ( .A1(G299), .A2(n703), .ZN(n704) );
  XOR2_X1 U793 ( .A(KEYINPUT96), .B(n704), .Z(n705) );
  OR2_X1 U794 ( .A1(n706), .A2(n705), .ZN(n707) );
  AND2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U796 ( .A(KEYINPUT29), .B(n709), .Z(n714) );
  XNOR2_X1 U797 ( .A(G2078), .B(KEYINPUT25), .ZN(n1010) );
  NOR2_X1 U798 ( .A1(n733), .A2(n1010), .ZN(n712) );
  INV_X1 U799 ( .A(G1961), .ZN(n948) );
  NOR2_X1 U800 ( .A1(n710), .A2(n948), .ZN(n711) );
  NOR2_X1 U801 ( .A1(n712), .A2(n711), .ZN(n720) );
  NAND2_X1 U802 ( .A1(G171), .A2(n720), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n714), .A2(n713), .ZN(n725) );
  NOR2_X1 U804 ( .A1(n728), .A2(n715), .ZN(n716) );
  NAND2_X1 U805 ( .A1(G8), .A2(n716), .ZN(n717) );
  XNOR2_X1 U806 ( .A(KEYINPUT30), .B(n717), .ZN(n718) );
  XOR2_X1 U807 ( .A(KEYINPUT97), .B(n718), .Z(n719) );
  NOR2_X1 U808 ( .A1(G168), .A2(n719), .ZN(n722) );
  NOR2_X1 U809 ( .A1(n720), .A2(G171), .ZN(n721) );
  NOR2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U811 ( .A(KEYINPUT31), .B(n723), .Z(n724) );
  NAND2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n732) );
  INV_X1 U813 ( .A(KEYINPUT98), .ZN(n726) );
  XNOR2_X1 U814 ( .A(n732), .B(n726), .ZN(n727) );
  NOR2_X1 U815 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U816 ( .A1(n730), .A2(n729), .ZN(n743) );
  AND2_X1 U817 ( .A1(G286), .A2(G8), .ZN(n731) );
  NAND2_X1 U818 ( .A1(n732), .A2(n731), .ZN(n740) );
  INV_X1 U819 ( .A(G8), .ZN(n738) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n811), .ZN(n735) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U823 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U824 ( .A1(n738), .A2(n737), .ZN(n739) );
  AND2_X1 U825 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U826 ( .A(n741), .B(KEYINPUT32), .ZN(n742) );
  NAND2_X1 U827 ( .A1(n743), .A2(n742), .ZN(n807) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n937) );
  NOR2_X1 U829 ( .A1(n930), .A2(n937), .ZN(n744) );
  XOR2_X1 U830 ( .A(KEYINPUT99), .B(n744), .Z(n745) );
  NAND2_X1 U831 ( .A1(n807), .A2(n745), .ZN(n749) );
  NAND2_X1 U832 ( .A1(G288), .A2(G1976), .ZN(n746) );
  XNOR2_X1 U833 ( .A(n746), .B(KEYINPUT100), .ZN(n932) );
  NOR2_X1 U834 ( .A1(n811), .A2(n747), .ZN(n748) );
  NOR2_X1 U835 ( .A1(KEYINPUT33), .A2(n750), .ZN(n751) );
  NOR2_X1 U836 ( .A1(n752), .A2(n751), .ZN(n803) );
  XOR2_X1 U837 ( .A(G1981), .B(G305), .Z(n919) );
  XNOR2_X1 U838 ( .A(KEYINPUT37), .B(G2067), .ZN(n762) );
  NAND2_X1 U839 ( .A1(G116), .A2(n867), .ZN(n754) );
  NAND2_X1 U840 ( .A1(G128), .A2(n868), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U842 ( .A(n755), .B(KEYINPUT35), .ZN(n760) );
  NAND2_X1 U843 ( .A1(G104), .A2(n874), .ZN(n757) );
  NAND2_X1 U844 ( .A1(G140), .A2(n865), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U846 ( .A(KEYINPUT34), .B(n758), .Z(n759) );
  NAND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U848 ( .A(n761), .B(KEYINPUT36), .Z(n882) );
  AND2_X1 U849 ( .A1(n762), .A2(n882), .ZN(n981) );
  NOR2_X1 U850 ( .A1(n762), .A2(n882), .ZN(n982) );
  NOR2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n793) );
  NAND2_X1 U852 ( .A1(n982), .A2(n793), .ZN(n796) );
  NAND2_X1 U853 ( .A1(G117), .A2(n867), .ZN(n766) );
  NAND2_X1 U854 ( .A1(G129), .A2(n868), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n874), .A2(G105), .ZN(n767) );
  XOR2_X1 U857 ( .A(KEYINPUT38), .B(n767), .Z(n768) );
  NOR2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U859 ( .A(n770), .B(KEYINPUT92), .ZN(n772) );
  NAND2_X1 U860 ( .A1(G141), .A2(n865), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n887) );
  NOR2_X1 U862 ( .A1(G1996), .A2(n887), .ZN(n986) );
  NAND2_X1 U863 ( .A1(G107), .A2(n867), .ZN(n773) );
  XOR2_X1 U864 ( .A(KEYINPUT90), .B(n773), .Z(n778) );
  NAND2_X1 U865 ( .A1(G95), .A2(n874), .ZN(n775) );
  NAND2_X1 U866 ( .A1(G131), .A2(n865), .ZN(n774) );
  NAND2_X1 U867 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U868 ( .A(KEYINPUT91), .B(n776), .Z(n777) );
  NOR2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n868), .A2(G119), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n862) );
  NAND2_X1 U872 ( .A1(G1991), .A2(n862), .ZN(n782) );
  NAND2_X1 U873 ( .A1(G1996), .A2(n887), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n980) );
  NOR2_X1 U875 ( .A1(G1986), .A2(G290), .ZN(n783) );
  NOR2_X1 U876 ( .A1(G1991), .A2(n862), .ZN(n989) );
  NOR2_X1 U877 ( .A1(n783), .A2(n989), .ZN(n784) );
  XOR2_X1 U878 ( .A(KEYINPUT101), .B(n784), .Z(n785) );
  NOR2_X1 U879 ( .A1(n980), .A2(n785), .ZN(n786) );
  XNOR2_X1 U880 ( .A(n786), .B(KEYINPUT102), .ZN(n787) );
  NOR2_X1 U881 ( .A1(n986), .A2(n787), .ZN(n788) );
  XOR2_X1 U882 ( .A(n788), .B(KEYINPUT39), .Z(n789) );
  XNOR2_X1 U883 ( .A(KEYINPUT103), .B(n789), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n796), .A2(n790), .ZN(n791) );
  XOR2_X1 U885 ( .A(KEYINPUT104), .B(n791), .Z(n792) );
  NOR2_X1 U886 ( .A1(n981), .A2(n792), .ZN(n794) );
  INV_X1 U887 ( .A(n793), .ZN(n798) );
  NOR2_X1 U888 ( .A1(n794), .A2(n798), .ZN(n795) );
  XOR2_X1 U889 ( .A(n795), .B(KEYINPUT105), .Z(n812) );
  INV_X1 U890 ( .A(n796), .ZN(n800) );
  XNOR2_X1 U891 ( .A(G1986), .B(G290), .ZN(n924) );
  NOR2_X1 U892 ( .A1(n980), .A2(n924), .ZN(n797) );
  NOR2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U895 ( .A1(n812), .A2(n801), .ZN(n804) );
  AND2_X1 U896 ( .A1(n919), .A2(n804), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n819) );
  INV_X1 U898 ( .A(n804), .ZN(n817) );
  NOR2_X1 U899 ( .A1(G2090), .A2(G303), .ZN(n805) );
  NAND2_X1 U900 ( .A1(G8), .A2(n805), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  AND2_X1 U902 ( .A1(n808), .A2(n811), .ZN(n815) );
  NOR2_X1 U903 ( .A1(G1981), .A2(G305), .ZN(n809) );
  XOR2_X1 U904 ( .A(n809), .B(KEYINPUT24), .Z(n810) );
  NOR2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n813) );
  OR2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n816) );
  OR2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U910 ( .A(n820), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U911 ( .A1(n821), .A2(G2106), .ZN(n822) );
  XOR2_X1 U912 ( .A(KEYINPUT107), .B(n822), .Z(G217) );
  NAND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n823) );
  XOR2_X1 U914 ( .A(KEYINPUT108), .B(n823), .Z(n824) );
  NAND2_X1 U915 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U918 ( .A(n827), .ZN(G319) );
  XOR2_X1 U919 ( .A(G2100), .B(G2096), .Z(n829) );
  XNOR2_X1 U920 ( .A(KEYINPUT42), .B(G2678), .ZN(n828) );
  XNOR2_X1 U921 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U922 ( .A(KEYINPUT43), .B(G2090), .Z(n831) );
  XNOR2_X1 U923 ( .A(G2067), .B(G2072), .ZN(n830) );
  XNOR2_X1 U924 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U925 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U926 ( .A(G2084), .B(G2078), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n835), .B(n834), .ZN(G227) );
  XOR2_X1 U928 ( .A(G1986), .B(G1971), .Z(n837) );
  XNOR2_X1 U929 ( .A(G1966), .B(G1961), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U931 ( .A(G1991), .B(G1981), .Z(n839) );
  XNOR2_X1 U932 ( .A(G1996), .B(G1956), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U934 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U935 ( .A(KEYINPUT109), .B(G2474), .ZN(n842) );
  XNOR2_X1 U936 ( .A(n843), .B(n842), .ZN(n845) );
  XOR2_X1 U937 ( .A(G1976), .B(KEYINPUT41), .Z(n844) );
  XNOR2_X1 U938 ( .A(n845), .B(n844), .ZN(G229) );
  NAND2_X1 U939 ( .A1(G124), .A2(n868), .ZN(n846) );
  XNOR2_X1 U940 ( .A(n846), .B(KEYINPUT110), .ZN(n847) );
  XNOR2_X1 U941 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U942 ( .A1(G100), .A2(n874), .ZN(n848) );
  NAND2_X1 U943 ( .A1(n849), .A2(n848), .ZN(n853) );
  NAND2_X1 U944 ( .A1(G112), .A2(n867), .ZN(n851) );
  NAND2_X1 U945 ( .A1(G136), .A2(n865), .ZN(n850) );
  NAND2_X1 U946 ( .A1(n851), .A2(n850), .ZN(n852) );
  NOR2_X1 U947 ( .A1(n853), .A2(n852), .ZN(G162) );
  NAND2_X1 U948 ( .A1(G118), .A2(n867), .ZN(n855) );
  NAND2_X1 U949 ( .A1(G130), .A2(n868), .ZN(n854) );
  NAND2_X1 U950 ( .A1(n855), .A2(n854), .ZN(n860) );
  NAND2_X1 U951 ( .A1(G106), .A2(n874), .ZN(n857) );
  NAND2_X1 U952 ( .A1(G142), .A2(n865), .ZN(n856) );
  NAND2_X1 U953 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U954 ( .A(KEYINPUT45), .B(n858), .Z(n859) );
  NOR2_X1 U955 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U956 ( .A(n988), .B(n861), .ZN(n886) );
  XNOR2_X1 U957 ( .A(KEYINPUT46), .B(KEYINPUT116), .ZN(n864) );
  XNOR2_X1 U958 ( .A(n862), .B(KEYINPUT48), .ZN(n863) );
  XNOR2_X1 U959 ( .A(n864), .B(n863), .ZN(n881) );
  NAND2_X1 U960 ( .A1(n865), .A2(G139), .ZN(n866) );
  XNOR2_X1 U961 ( .A(n866), .B(KEYINPUT112), .ZN(n879) );
  XNOR2_X1 U962 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n873) );
  NAND2_X1 U963 ( .A1(n867), .A2(G115), .ZN(n871) );
  NAND2_X1 U964 ( .A1(n868), .A2(G127), .ZN(n869) );
  XOR2_X1 U965 ( .A(KEYINPUT113), .B(n869), .Z(n870) );
  NAND2_X1 U966 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U967 ( .A(n873), .B(n872), .Z(n877) );
  NAND2_X1 U968 ( .A1(G103), .A2(n874), .ZN(n875) );
  XNOR2_X1 U969 ( .A(KEYINPUT111), .B(n875), .ZN(n876) );
  NOR2_X1 U970 ( .A1(n877), .A2(n876), .ZN(n878) );
  NAND2_X1 U971 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U972 ( .A(n880), .B(KEYINPUT115), .ZN(n974) );
  XOR2_X1 U973 ( .A(n881), .B(n974), .Z(n884) );
  XOR2_X1 U974 ( .A(n882), .B(G162), .Z(n883) );
  XNOR2_X1 U975 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U976 ( .A(n886), .B(n885), .ZN(n890) );
  XNOR2_X1 U977 ( .A(G160), .B(G164), .ZN(n888) );
  XNOR2_X1 U978 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U979 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U980 ( .A1(G37), .A2(n891), .ZN(G395) );
  XOR2_X1 U981 ( .A(KEYINPUT117), .B(G286), .Z(n893) );
  XNOR2_X1 U982 ( .A(G301), .B(n922), .ZN(n892) );
  XNOR2_X1 U983 ( .A(n893), .B(n892), .ZN(n895) );
  XNOR2_X1 U984 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U985 ( .A1(G37), .A2(n896), .ZN(G397) );
  XOR2_X1 U986 ( .A(G2443), .B(G2451), .Z(n898) );
  XNOR2_X1 U987 ( .A(G2446), .B(G2454), .ZN(n897) );
  XNOR2_X1 U988 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U989 ( .A(n899), .B(G2427), .Z(n901) );
  XNOR2_X1 U990 ( .A(G1341), .B(G1348), .ZN(n900) );
  XNOR2_X1 U991 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U992 ( .A(G2435), .B(KEYINPUT106), .Z(n903) );
  XNOR2_X1 U993 ( .A(G2430), .B(G2438), .ZN(n902) );
  XNOR2_X1 U994 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U995 ( .A(n905), .B(n904), .Z(n906) );
  NAND2_X1 U996 ( .A1(G14), .A2(n906), .ZN(n918) );
  NAND2_X1 U997 ( .A1(G319), .A2(n918), .ZN(n909) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U999 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1000 ( .A1(n909), .A2(n908), .ZN(n911) );
  NOR2_X1 U1001 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1002 ( .A1(n911), .A2(n910), .ZN(G225) );
  XOR2_X1 U1003 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  XNOR2_X1 U1005 ( .A(n927), .B(n912), .ZN(n913) );
  NOR2_X1 U1006 ( .A1(G860), .A2(n913), .ZN(n914) );
  XOR2_X1 U1007 ( .A(n915), .B(n914), .Z(G145) );
  INV_X1 U1008 ( .A(G132), .ZN(G219) );
  INV_X1 U1009 ( .A(G120), .ZN(G236) );
  INV_X1 U1010 ( .A(G96), .ZN(G221) );
  INV_X1 U1011 ( .A(G82), .ZN(G220) );
  INV_X1 U1012 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(G325) );
  INV_X1 U1014 ( .A(G325), .ZN(G261) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  INV_X1 U1016 ( .A(n918), .ZN(G401) );
  XNOR2_X1 U1017 ( .A(KEYINPUT56), .B(G16), .ZN(n946) );
  XNOR2_X1 U1018 ( .A(G1966), .B(G168), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n921), .B(KEYINPUT57), .ZN(n944) );
  XNOR2_X1 U1021 ( .A(n922), .B(G1348), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(G1956), .B(G299), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n942) );
  XNOR2_X1 U1025 ( .A(G301), .B(G1961), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n927), .B(G1341), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n940) );
  XOR2_X1 U1028 ( .A(n930), .B(KEYINPUT122), .Z(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(n933), .B(KEYINPUT123), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(G1971), .A2(G303), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(n938), .B(KEYINPUT124), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(n947), .B(KEYINPUT125), .ZN(n973) );
  XNOR2_X1 U1040 ( .A(G5), .B(n948), .ZN(n969) );
  XNOR2_X1 U1041 ( .A(KEYINPUT59), .B(G4), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(n949), .B(KEYINPUT126), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(G1348), .B(n950), .ZN(n954) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G19), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G1981), .B(G6), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(G20), .B(G1956), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1050 ( .A(KEYINPUT60), .B(n957), .Z(n959) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G21), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(KEYINPUT127), .B(n960), .ZN(n967) );
  XNOR2_X1 U1054 ( .A(G1971), .B(G22), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(G23), .B(G1976), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n964) );
  XOR2_X1 U1057 ( .A(G1986), .B(G24), .Z(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(KEYINPUT58), .B(n965), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(KEYINPUT61), .B(n970), .ZN(n971) );
  NOR2_X1 U1063 ( .A1(n971), .A2(G16), .ZN(n972) );
  NOR2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n1002) );
  XNOR2_X1 U1065 ( .A(G2072), .B(n974), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n975), .B(KEYINPUT121), .ZN(n977) );
  XOR2_X1 U1067 ( .A(G2078), .B(G164), .Z(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1069 ( .A(KEYINPUT50), .B(n978), .Z(n997) );
  XOR2_X1 U1070 ( .A(G160), .B(G2084), .Z(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n984) );
  NOR2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n994) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1076 ( .A(KEYINPUT51), .B(n987), .Z(n992) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1078 ( .A(KEYINPUT119), .B(n990), .Z(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1081 ( .A(KEYINPUT120), .B(n995), .Z(n996) );
  NOR2_X1 U1082 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1083 ( .A(KEYINPUT52), .B(n998), .ZN(n999) );
  INV_X1 U1084 ( .A(KEYINPUT55), .ZN(n1020) );
  NAND2_X1 U1085 ( .A1(n999), .A2(n1020), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1000), .A2(G29), .ZN(n1001) );
  NAND2_X1 U1087 ( .A1(n1002), .A2(n1001), .ZN(n1025) );
  XNOR2_X1 U1088 ( .A(G2090), .B(G35), .ZN(n1015) );
  XNOR2_X1 U1089 ( .A(G1996), .B(G32), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(G33), .B(G2072), .ZN(n1003) );
  NOR2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1009) );
  XOR2_X1 U1092 ( .A(G1991), .B(G25), .Z(n1005) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(G28), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G26), .B(G2067), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(G27), .B(n1010), .Z(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(KEYINPUT53), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XOR2_X1 U1101 ( .A(G2084), .B(G34), .Z(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT54), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(n1020), .B(n1019), .ZN(n1022) );
  INV_X1 U1105 ( .A(G29), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(G11), .A2(n1023), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(n1026), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

