//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1244, new_n1245;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AOI22_X1  g0006(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT65), .B(G68), .Z(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n203), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT64), .Z(new_n228));
  INV_X1    g0028(.A(G68), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n214), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n206), .B(new_n224), .C1(new_n228), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G97), .B(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT66), .ZN(new_n249));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(KEYINPUT66), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n258), .B1(new_n215), .B2(new_n261), .C1(new_n216), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n263), .B(new_n264), .C1(G107), .C2(new_n258), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  OAI211_X1 g0071(.A(G1), .B(G13), .C1(new_n254), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n267), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n273), .B2(new_n211), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT70), .ZN(new_n275));
  AOI21_X1  g0075(.A(G169), .B1(new_n265), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT72), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G77), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n225), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(G1), .B2(new_n226), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n210), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G20), .A2(G77), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n226), .A2(G33), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT15), .B(G87), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT71), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n285), .B1(new_n286), .B2(new_n287), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  AOI211_X1 g0091(.A(new_n279), .B(new_n284), .C1(new_n291), .C2(new_n281), .ZN(new_n292));
  OR3_X1    g0092(.A1(new_n276), .A2(new_n277), .A3(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n265), .A2(new_n275), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n277), .B1(new_n276), .B2(new_n292), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G97), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT74), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n261), .A2(new_n209), .B1(new_n215), .B2(new_n262), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n258), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n270), .B1(new_n216), .B2(new_n273), .C1(new_n302), .C2(new_n272), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT13), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(KEYINPUT75), .ZN(new_n307));
  INV_X1    g0107(.A(G13), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(G1), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n218), .A2(KEYINPUT12), .A3(G20), .A4(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n278), .A2(G68), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n310), .B1(KEYINPUT12), .B2(new_n311), .C1(new_n283), .C2(new_n229), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT76), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n217), .A2(new_n226), .B1(new_n210), .B2(new_n286), .ZN(new_n314));
  INV_X1    g0114(.A(new_n288), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n208), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n281), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g0117(.A(new_n317), .B(KEYINPUT11), .Z(new_n318));
  OR2_X1    g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(G200), .B2(new_n304), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n306), .A2(KEYINPUT75), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n307), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT14), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n304), .A2(new_n324), .A3(G169), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n304), .B2(G169), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n304), .A2(new_n295), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n319), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OR3_X1    g0130(.A1(new_n323), .A2(new_n330), .A3(KEYINPUT77), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT77), .B1(new_n330), .B2(new_n323), .ZN(new_n332));
  INV_X1    g0132(.A(new_n278), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(G50), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n283), .B2(G50), .ZN(new_n335));
  XOR2_X1   g0135(.A(new_n335), .B(KEYINPUT69), .Z(new_n336));
  INV_X1    g0136(.A(G150), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n290), .A2(new_n286), .B1(new_n337), .B2(new_n315), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT68), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n208), .A2(new_n214), .A3(new_n229), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(G20), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n336), .B1(new_n282), .B2(new_n342), .ZN(new_n343));
  XOR2_X1   g0143(.A(new_n343), .B(KEYINPUT9), .Z(new_n344));
  INV_X1    g0144(.A(KEYINPUT10), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT67), .B(G1698), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(G222), .B1(G223), .B2(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n258), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n264), .C1(G77), .C2(new_n258), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(new_n270), .C1(new_n209), .C2(new_n273), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n305), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT73), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT73), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n350), .B2(G200), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n352), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  OR3_X1    g0155(.A1(new_n344), .A2(new_n345), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n345), .B1(new_n344), .B2(new_n355), .ZN(new_n357));
  INV_X1    g0157(.A(G169), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n350), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n343), .B(new_n359), .C1(G179), .C2(new_n350), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n356), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  AND4_X1   g0161(.A1(new_n298), .A2(new_n331), .A3(new_n332), .A4(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n254), .A2(new_n220), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AND2_X1   g0164(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n365));
  NOR2_X1   g0165(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n251), .B1(new_n367), .B2(G33), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n209), .A2(new_n262), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(new_n346), .B2(G223), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n364), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n269), .B1(new_n371), .B2(new_n264), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n272), .A2(G232), .A3(new_n267), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT79), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(G223), .B1(new_n259), .B2(new_n260), .ZN(new_n375));
  INV_X1    g0175(.A(new_n369), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT78), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n253), .ZN(new_n379));
  NAND2_X1  g0179(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(G33), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n255), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n363), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n270), .B(new_n373), .C1(new_n383), .C2(new_n272), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT79), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n358), .B1(new_n374), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT80), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n384), .A2(G179), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n290), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n333), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n283), .B2(new_n392), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n217), .A2(G58), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n230), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(G20), .B1(G159), .B2(new_n288), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n379), .A2(new_n380), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(new_n254), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(new_n226), .A3(new_n256), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n252), .A2(new_n257), .A3(new_n226), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n399), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT16), .B1(new_n405), .B2(new_n217), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT7), .B1(new_n382), .B2(G20), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n381), .A2(new_n399), .A3(new_n226), .A4(new_n255), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(G68), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n398), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n398), .A2(new_n406), .B1(new_n410), .B2(KEYINPUT16), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n395), .B1(new_n411), .B2(new_n282), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n384), .A2(new_n385), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n375), .A2(new_n376), .B1(new_n381), .B2(new_n255), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n264), .B1(new_n414), .B2(new_n363), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n415), .A2(KEYINPUT79), .A3(new_n270), .A4(new_n373), .ZN(new_n416));
  AOI21_X1  g0216(.A(G169), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT80), .B1(new_n417), .B2(new_n389), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n391), .A2(new_n412), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n391), .A2(new_n412), .A3(new_n418), .A4(KEYINPUT18), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n413), .A2(new_n416), .ZN(new_n424));
  INV_X1    g0224(.A(G200), .ZN(new_n425));
  INV_X1    g0225(.A(new_n384), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n424), .A2(new_n425), .B1(new_n305), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n406), .A2(new_n398), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n410), .A2(KEYINPUT16), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n394), .B1(new_n431), .B2(new_n281), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(KEYINPUT17), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n412), .B2(new_n427), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n423), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT81), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n294), .A2(G190), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n292), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n294), .A2(new_n425), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n362), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT83), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT5), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n447), .B2(G41), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n271), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n266), .A2(G45), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n447), .B2(G41), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n264), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G264), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G257), .A2(G1698), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n261), .B2(new_n221), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(new_n382), .B1(G33), .B2(G294), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n457), .B2(new_n272), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT84), .ZN(new_n459));
  INV_X1    g0259(.A(new_n451), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n447), .A2(G41), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n448), .A3(new_n461), .A4(new_n449), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n459), .B1(new_n462), .B2(new_n268), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n450), .A2(KEYINPUT84), .A3(new_n452), .A4(G274), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n425), .B1(new_n458), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n456), .A2(new_n382), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G294), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n264), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n471), .A2(new_n305), .A3(new_n465), .A4(new_n454), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n474));
  INV_X1    g0274(.A(G107), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT91), .B1(new_n475), .B2(G20), .ZN(new_n476));
  XOR2_X1   g0276(.A(new_n476), .B(KEYINPUT23), .Z(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  AOI21_X1  g0278(.A(G20), .B1(new_n381), .B2(new_n255), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(G87), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n226), .B(G87), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n252), .B2(new_n257), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n474), .B(new_n477), .C1(new_n480), .C2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT24), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI211_X1 g0287(.A(G20), .B(new_n220), .C1(new_n381), .C2(new_n255), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n252), .A2(new_n257), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n488), .A2(new_n478), .B1(new_n489), .B2(new_n483), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n490), .A2(KEYINPUT24), .A3(new_n474), .A4(new_n477), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(new_n281), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT92), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT25), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n333), .B2(new_n475), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n493), .A2(KEYINPUT25), .ZN(new_n496));
  AND4_X1   g0296(.A1(new_n475), .A2(new_n333), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n281), .B(new_n333), .C1(new_n266), .C2(G33), .ZN(new_n498));
  AOI211_X1 g0298(.A(new_n495), .B(new_n497), .C1(new_n498), .C2(G107), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n473), .A2(new_n492), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n358), .B1(new_n458), .B2(new_n466), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n471), .A2(new_n295), .A3(new_n465), .A4(new_n454), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n499), .B2(new_n492), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT93), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n492), .A2(new_n499), .ZN(new_n506));
  INV_X1    g0306(.A(new_n503), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT93), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n473), .A2(new_n492), .A3(new_n499), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n278), .A2(G97), .ZN(new_n513));
  INV_X1    g0313(.A(new_n498), .ZN(new_n514));
  INV_X1    g0314(.A(G97), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n315), .A2(new_n210), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT6), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n515), .A2(new_n475), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n475), .A2(KEYINPUT6), .A3(G97), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n226), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n399), .B(G20), .C1(new_n400), .C2(new_n254), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(new_n256), .B1(new_n399), .B2(new_n403), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n518), .B(new_n525), .C1(new_n527), .C2(new_n475), .ZN(new_n528));
  AOI211_X1 g0328(.A(new_n513), .B(new_n516), .C1(new_n528), .C2(new_n281), .ZN(new_n529));
  OAI21_X1  g0329(.A(G244), .B1(new_n259), .B2(new_n260), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n382), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n530), .B1(new_n252), .B2(new_n257), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT82), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G283), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n258), .A2(KEYINPUT82), .A3(G250), .A4(G1698), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n535), .A2(new_n538), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n264), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n453), .A2(G257), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n542), .A2(G190), .A3(new_n465), .A4(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n543), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n466), .B(new_n545), .C1(new_n541), .C2(new_n264), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n529), .B(new_n544), .C1(new_n546), .C2(new_n425), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n528), .A2(new_n281), .ZN(new_n548));
  INV_X1    g0348(.A(new_n513), .ZN(new_n549));
  INV_X1    g0349(.A(new_n516), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n542), .A2(new_n295), .A3(new_n465), .A4(new_n543), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n552), .C1(new_n546), .C2(G169), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n382), .A2(new_n226), .A3(G68), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n299), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(G20), .B1(new_n300), .B2(KEYINPUT19), .ZN(new_n557));
  NOR3_X1   g0357(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n554), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(new_n281), .B1(new_n333), .B2(new_n287), .ZN(new_n560));
  INV_X1    g0360(.A(G116), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n264), .B1(new_n254), .B2(new_n561), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n261), .A2(new_n216), .B1(new_n211), .B2(new_n262), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n562), .B1(new_n563), .B2(new_n382), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n451), .A2(KEYINPUT85), .A3(G250), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT85), .ZN(new_n566));
  AOI21_X1  g0366(.A(G274), .B1(new_n566), .B2(G250), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n565), .B(new_n272), .C1(new_n451), .C2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G200), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n498), .A2(G87), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n560), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n570), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G190), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n514), .A2(new_n287), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n560), .A2(new_n577), .B1(new_n358), .B2(new_n570), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n575), .A2(new_n295), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n574), .A2(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n547), .A2(new_n553), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT86), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n346), .A2(G257), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n582), .B1(new_n368), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n489), .A2(G303), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n382), .A2(KEYINPUT86), .A3(G257), .A4(new_n346), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n382), .A2(G264), .A3(G1698), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n264), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n463), .A2(new_n464), .B1(new_n453), .B2(G270), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n498), .A2(G116), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n309), .A2(G20), .A3(new_n561), .ZN(new_n593));
  XNOR2_X1  g0393(.A(new_n593), .B(KEYINPUT87), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n561), .A2(G20), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n281), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT88), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n539), .B(new_n226), .C1(G33), .C2(new_n515), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT20), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n597), .A2(KEYINPUT88), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT88), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n281), .B2(new_n596), .ZN(new_n603));
  OAI211_X1 g0403(.A(KEYINPUT20), .B(new_n599), .C1(new_n601), .C2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n592), .B(new_n595), .C1(new_n600), .C2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n591), .A2(new_n606), .A3(G169), .ZN(new_n607));
  NOR2_X1   g0407(.A1(KEYINPUT89), .A2(KEYINPUT21), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n589), .A2(G179), .A3(new_n590), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n607), .A2(new_n608), .B1(new_n610), .B2(new_n606), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n591), .A2(G200), .ZN(new_n612));
  INV_X1    g0412(.A(new_n606), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n612), .B(new_n613), .C1(new_n305), .C2(new_n591), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n609), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n581), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n445), .A2(new_n512), .A3(new_n616), .ZN(G372));
  AND2_X1   g0417(.A1(new_n547), .A2(new_n553), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT94), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n573), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n560), .A2(KEYINPUT94), .A3(new_n571), .A4(new_n572), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n576), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n578), .A2(new_n579), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n609), .A2(new_n611), .A3(new_n508), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n618), .A2(new_n625), .A3(new_n510), .A4(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n553), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n625), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n580), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT26), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n627), .A2(new_n623), .A3(new_n630), .A4(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n445), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n298), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n322), .B(new_n436), .C1(new_n330), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n423), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n356), .A3(new_n357), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n360), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n634), .A2(new_n640), .ZN(G369));
  NAND2_X1  g0441(.A1(new_n309), .A2(new_n226), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT95), .ZN(new_n643));
  OR3_X1    g0443(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT27), .ZN(new_n644));
  INV_X1    g0444(.A(G213), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n642), .B2(KEYINPUT27), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n643), .B1(new_n642), .B2(KEYINPUT27), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G343), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n506), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n512), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n650), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n508), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n609), .A2(new_n611), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n613), .A2(new_n653), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n615), .B2(new_n657), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n656), .A2(new_n653), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n512), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n504), .B2(new_n653), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n662), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(new_n204), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(G41), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G1), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n558), .A2(new_n561), .ZN(new_n673));
  OAI22_X1  g0473(.A1(new_n672), .A2(new_n673), .B1(new_n231), .B2(new_n671), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT28), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n633), .A2(new_n653), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(KEYINPUT29), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT26), .B1(new_n624), .B2(new_n553), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n628), .A2(new_n629), .A3(new_n580), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n627), .A2(new_n623), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n653), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n677), .B1(KEYINPUT29), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT31), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n542), .A2(new_n465), .A3(new_n543), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n471), .A2(new_n465), .A3(new_n454), .ZN(new_n685));
  AOI21_X1  g0485(.A(G179), .B1(new_n589), .B2(new_n590), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n458), .A2(new_n570), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n542), .A2(new_n465), .A3(new_n688), .A4(new_n543), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n589), .A2(G179), .A3(new_n590), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT30), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n546), .A2(new_n692), .A3(new_n610), .A4(new_n688), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n570), .A2(new_n687), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n650), .B1(new_n694), .B2(KEYINPUT96), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n691), .A2(new_n693), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n684), .A2(new_n685), .A3(new_n570), .A4(new_n686), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(KEYINPUT96), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n683), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n547), .A2(new_n553), .A3(new_n580), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n609), .A2(new_n611), .A3(new_n614), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n512), .A2(new_n701), .A3(new_n702), .A4(new_n653), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT97), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT97), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n616), .A2(new_n705), .A3(new_n512), .A4(new_n653), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n696), .A2(new_n697), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n650), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n700), .A2(new_n704), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n682), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n675), .B1(new_n712), .B2(G1), .ZN(G364));
  NOR2_X1   g0513(.A1(G13), .A2(G33), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n659), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n225), .B1(G20), .B2(new_n358), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT32), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n226), .A2(G190), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G179), .A2(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G159), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(G190), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n720), .A2(new_n725), .B1(new_n728), .B2(new_n515), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n489), .B(new_n729), .C1(new_n720), .C2(new_n725), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n295), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n721), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n226), .A2(new_n305), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n425), .A2(G179), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n730), .B1(new_n210), .B2(new_n732), .C1(new_n220), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n733), .A2(new_n731), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n214), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n295), .A2(new_n425), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n208), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n721), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n721), .A2(new_n734), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n742), .A2(new_n229), .B1(new_n743), .B2(new_n475), .ZN(new_n744));
  NOR4_X1   g0544(.A1(new_n736), .A2(new_n738), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n737), .ZN(new_n746));
  INV_X1    g0546(.A(new_n732), .ZN(new_n747));
  AOI22_X1  g0547(.A1(G322), .A2(new_n746), .B1(new_n747), .B2(G311), .ZN(new_n748));
  INV_X1    g0548(.A(new_n723), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G329), .ZN(new_n750));
  INV_X1    g0550(.A(G326), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n748), .B(new_n750), .C1(new_n751), .C2(new_n740), .ZN(new_n752));
  INV_X1    g0552(.A(G283), .ZN(new_n753));
  XOR2_X1   g0553(.A(KEYINPUT33), .B(G317), .Z(new_n754));
  OAI221_X1 g0554(.A(new_n489), .B1(new_n753), .B2(new_n743), .C1(new_n742), .C2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G294), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n728), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G303), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n735), .A2(new_n758), .ZN(new_n759));
  NOR4_X1   g0559(.A1(new_n752), .A2(new_n755), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n719), .B1(new_n745), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n382), .A2(new_n669), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G45), .B2(new_n231), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT98), .Z(new_n764));
  INV_X1    g0564(.A(G45), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(new_n765), .B2(new_n244), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n258), .A2(G355), .A3(new_n204), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n766), .B(new_n767), .C1(G116), .C2(new_n204), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n716), .A2(new_n719), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n308), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n672), .B1(G45), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n718), .A2(new_n761), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n659), .A2(G330), .ZN(new_n774));
  INV_X1    g0574(.A(new_n772), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n660), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n773), .B1(new_n774), .B2(new_n776), .ZN(G396));
  NOR2_X1   g0577(.A1(new_n292), .A2(new_n653), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n635), .B2(KEYINPUT102), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n298), .A2(new_n442), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT102), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n298), .A2(new_n782), .A3(new_n778), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n714), .ZN(new_n785));
  INV_X1    g0585(.A(new_n743), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G87), .ZN(new_n787));
  INV_X1    g0587(.A(G311), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n788), .B2(new_n723), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n747), .A2(G116), .B1(new_n727), .B2(G97), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n756), .B2(new_n737), .ZN(new_n791));
  INV_X1    g0591(.A(new_n740), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n789), .B(new_n791), .C1(G303), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n735), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n258), .B1(G107), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT99), .B(G283), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n793), .B(new_n795), .C1(new_n742), .C2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT100), .Z(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT101), .B(G143), .Z(new_n800));
  AOI22_X1  g0600(.A1(new_n746), .A2(new_n800), .B1(new_n747), .B2(G159), .ZN(new_n801));
  INV_X1    g0601(.A(G137), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n801), .B1(new_n802), .B2(new_n740), .C1(new_n337), .C2(new_n742), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT34), .Z(new_n804));
  INV_X1    g0604(.A(G132), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n735), .A2(new_n208), .B1(new_n723), .B2(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n368), .B(new_n806), .C1(G68), .C2(new_n786), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n214), .B2(new_n728), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n719), .B1(new_n799), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n719), .A2(new_n714), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n210), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n785), .A2(new_n772), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n784), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n814), .A2(new_n633), .A3(new_n653), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(KEYINPUT103), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n710), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n676), .A2(new_n784), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n817), .B(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n813), .B1(new_n819), .B2(new_n772), .ZN(G384));
  NAND2_X1  g0620(.A1(new_n522), .A2(new_n523), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT104), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n561), .B1(new_n822), .B2(KEYINPUT35), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n823), .B(new_n228), .C1(KEYINPUT35), .C2(new_n822), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT36), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n396), .A2(G77), .A3(new_n232), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(G50), .B2(new_n229), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n827), .A2(G1), .A3(new_n308), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n771), .A2(new_n266), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT16), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n410), .A2(KEYINPUT106), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(KEYINPUT106), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n398), .A2(new_n409), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n281), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n395), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n391), .A2(new_n418), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n428), .A2(new_n432), .ZN(new_n837));
  INV_X1    g0637(.A(new_n648), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT37), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n412), .A2(new_n838), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n419), .A2(new_n837), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n839), .B1(new_n423), .B2(new_n436), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT38), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n839), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n437), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n851), .B2(new_n845), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT39), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n437), .A2(new_n412), .A3(new_n838), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n419), .A2(new_n837), .A3(new_n843), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n844), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT38), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n855), .B1(new_n860), .B2(new_n849), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n330), .A2(new_n653), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n635), .A2(new_n653), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n865), .A2(KEYINPUT105), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(KEYINPUT105), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n815), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n319), .A2(new_n650), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n322), .B(new_n869), .C1(new_n328), .C2(new_n329), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n330), .A2(new_n650), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n873), .A2(new_n853), .B1(new_n423), .B2(new_n838), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n864), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n444), .A2(new_n682), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(new_n639), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n875), .B(new_n877), .Z(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT40), .B1(new_n860), .B2(new_n849), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT96), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n653), .B1(new_n707), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n700), .A2(new_n704), .A3(new_n706), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n784), .B1(new_n870), .B2(new_n871), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n883), .B(new_n884), .C1(new_n849), .C2(new_n852), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT107), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT107), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n887), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n886), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n893), .A2(new_n883), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n879), .A2(new_n885), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n887), .A2(new_n891), .A3(new_n888), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n891), .B1(new_n887), .B2(new_n888), .ZN(new_n897));
  OAI211_X1 g0697(.A(G330), .B(new_n895), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n445), .A2(G330), .A3(new_n883), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n894), .A2(new_n445), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n829), .B1(new_n878), .B2(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT108), .Z(new_n902));
  NOR2_X1   g0702(.A1(new_n878), .A2(new_n900), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT109), .Z(new_n904));
  OAI211_X1 g0704(.A(new_n825), .B(new_n828), .C1(new_n902), .C2(new_n904), .ZN(G367));
  AOI21_X1  g0705(.A(new_n266), .B1(new_n771), .B2(G45), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n666), .B1(new_n655), .B2(new_n663), .ZN(new_n907));
  INV_X1    g0707(.A(new_n660), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n662), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n711), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n618), .B1(new_n529), .B2(new_n653), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n553), .B2(new_n653), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n667), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n914));
  XNOR2_X1  g0714(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n667), .A2(new_n912), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT45), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n712), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n670), .B(KEYINPUT41), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n906), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n665), .A2(new_n911), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT42), .Z(new_n926));
  OAI21_X1  g0726(.A(new_n553), .B1(new_n911), .B2(new_n508), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n927), .A2(new_n653), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n653), .B1(new_n560), .B2(new_n572), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT110), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n625), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n623), .B2(new_n931), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n929), .B1(KEYINPUT43), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT111), .Z(new_n936));
  NAND2_X1  g0736(.A1(new_n661), .A2(new_n912), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n934), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n924), .A2(new_n939), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n792), .A2(new_n800), .B1(new_n794), .B2(G58), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n941), .B1(new_n229), .B2(new_n728), .C1(new_n337), .C2(new_n737), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n742), .A2(new_n724), .B1(new_n743), .B2(new_n210), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n942), .A2(new_n489), .A3(new_n943), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n944), .B1(new_n208), .B2(new_n732), .C1(new_n802), .C2(new_n723), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n794), .A2(G116), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT46), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n382), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(G311), .A2(new_n792), .B1(new_n786), .B2(G97), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(new_n756), .C2(new_n742), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n747), .A2(new_n796), .B1(new_n727), .B2(G107), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT113), .Z(new_n952));
  AOI211_X1 g0752(.A(new_n950), .B(new_n952), .C1(G317), .C2(new_n749), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n758), .B2(new_n737), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n946), .A2(new_n947), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n945), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT47), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n719), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n933), .A2(new_n717), .ZN(new_n959));
  INV_X1    g0759(.A(new_n762), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n769), .B1(new_n204), .B2(new_n287), .C1(new_n236), .C2(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n958), .A2(new_n772), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n940), .A2(new_n962), .ZN(G387));
  AOI21_X1  g0763(.A(new_n671), .B1(new_n711), .B2(new_n909), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n910), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n775), .B1(new_n655), .B2(new_n716), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n368), .B1(new_n561), .B2(new_n743), .ZN(new_n967));
  INV_X1    g0767(.A(new_n742), .ZN(new_n968));
  AOI22_X1  g0768(.A1(G322), .A2(new_n792), .B1(new_n968), .B2(G311), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n969), .B1(new_n758), .B2(new_n732), .C1(new_n970), .C2(new_n737), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT48), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n756), .B2(new_n735), .C1(new_n728), .C2(new_n797), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT49), .Z(new_n974));
  AOI211_X1 g0774(.A(new_n967), .B(new_n974), .C1(G326), .C2(new_n749), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n737), .A2(new_n208), .B1(new_n732), .B2(new_n229), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n728), .A2(new_n287), .ZN(new_n977));
  XOR2_X1   g0777(.A(KEYINPUT115), .B(G150), .Z(new_n978));
  AOI211_X1 g0778(.A(new_n976), .B(new_n977), .C1(new_n749), .C2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n515), .B2(new_n743), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G159), .A2(new_n792), .B1(new_n794), .B2(G77), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n290), .B2(new_n742), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n980), .A2(new_n368), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n719), .B1(new_n975), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n762), .B1(new_n240), .B2(new_n765), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n258), .A2(new_n204), .A3(new_n673), .ZN(new_n986));
  AOI211_X1 g0786(.A(G45), .B(new_n673), .C1(G68), .C2(G77), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n290), .A2(G50), .ZN(new_n988));
  XNOR2_X1  g0788(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n985), .A2(new_n986), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n204), .A2(G107), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n769), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n966), .A2(new_n984), .A3(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n965), .B(new_n994), .C1(new_n906), .C2(new_n909), .ZN(G393));
  XNOR2_X1  g0795(.A(new_n918), .B(new_n662), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(new_n906), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n769), .B1(new_n515), .B2(new_n204), .C1(new_n960), .C2(new_n247), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n912), .A2(new_n717), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n742), .A2(new_n208), .B1(new_n732), .B2(new_n290), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n382), .B1(new_n218), .B2(new_n735), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G77), .C2(new_n727), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n749), .A2(new_n800), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n740), .A2(new_n337), .B1(new_n737), .B2(new_n724), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT51), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n787), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(G322), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n742), .A2(new_n758), .B1(new_n723), .B2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n258), .B(new_n1008), .C1(G294), .C2(new_n747), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n794), .A2(new_n796), .B1(new_n786), .B2(G107), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(new_n561), .C2(new_n728), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n740), .A2(new_n970), .B1(new_n737), .B2(new_n788), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT52), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n1006), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT116), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n775), .B(new_n999), .C1(new_n719), .C2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n997), .B1(new_n998), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n996), .A2(new_n910), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1018), .A2(new_n670), .A3(new_n919), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT117), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT117), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1017), .A2(new_n1022), .A3(new_n1019), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(G390));
  NAND3_X1  g0824(.A1(new_n883), .A2(G330), .A3(new_n884), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n860), .A2(new_n849), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n863), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n814), .A2(new_n653), .A3(new_n680), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(KEYINPUT118), .A3(new_n865), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT118), .B1(new_n1029), .B2(new_n865), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1028), .B1(new_n1033), .B2(new_n872), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n861), .A2(new_n854), .B1(new_n873), .B2(new_n863), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1026), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n709), .A2(G330), .A3(new_n814), .A4(new_n872), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT119), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n873), .A2(new_n863), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n862), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1032), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n1030), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n872), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1041), .B(new_n1043), .C1(new_n1047), .C2(new_n1028), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n906), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1036), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n862), .A2(new_n714), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n811), .A2(new_n290), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n728), .A2(new_n724), .B1(new_n742), .B2(new_n802), .ZN(new_n1053));
  XOR2_X1   g0853(.A(KEYINPUT54), .B(G143), .Z(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT120), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1053), .B1(new_n747), .B2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT121), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1057), .A2(new_n258), .ZN(new_n1058));
  INV_X1    g0858(.A(G125), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n723), .C1(new_n805), .C2(new_n737), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n978), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n1061), .A2(KEYINPUT53), .A3(new_n735), .ZN(new_n1062));
  INV_X1    g0862(.A(G128), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n740), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(KEYINPUT53), .B1(new_n1061), .B2(new_n735), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n208), .B2(new_n743), .ZN(new_n1066));
  NOR4_X1   g0866(.A1(new_n1060), .A2(new_n1062), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n749), .A2(G294), .B1(new_n727), .B2(G77), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n229), .B2(new_n743), .C1(new_n561), .C2(new_n737), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n489), .B1(new_n220), .B2(new_n735), .C1(new_n753), .C2(new_n740), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n742), .A2(new_n475), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n732), .A2(new_n515), .ZN(new_n1072));
  NOR4_X1   g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n719), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1051), .A2(new_n772), .A3(new_n1052), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1050), .A2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT122), .Z(new_n1077));
  NAND3_X1  g0877(.A1(new_n883), .A2(G330), .A3(new_n814), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1039), .A2(new_n1040), .B1(new_n1046), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1046), .B1(new_n710), .B2(new_n784), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n1025), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1079), .A2(new_n1045), .B1(new_n868), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n877), .A2(new_n899), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1036), .A2(new_n1048), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n670), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1077), .A2(new_n1087), .ZN(G378));
  INV_X1    g0888(.A(KEYINPUT124), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n361), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n361), .A2(new_n1091), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n343), .A2(new_n838), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1092), .A2(new_n343), .A3(new_n838), .A4(new_n1093), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n898), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n890), .A2(new_n892), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1101), .A2(G330), .A3(new_n895), .A4(new_n1098), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1100), .A2(new_n1102), .A3(new_n875), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n875), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1089), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n875), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1098), .B1(new_n893), .B2(G330), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n898), .A2(new_n1099), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1100), .A2(new_n1102), .A3(new_n875), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(KEYINPUT124), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1105), .A2(new_n1111), .A3(new_n1049), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1098), .A2(new_n714), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n968), .A2(G97), .B1(new_n727), .B2(G68), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(new_n214), .B2(new_n743), .C1(new_n287), .C2(new_n732), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n723), .A2(new_n753), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n271), .B1(new_n735), .B2(new_n210), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n368), .B1(new_n475), .B2(new_n737), .C1(new_n561), .C2(new_n740), .ZN(new_n1118));
  NOR4_X1   g0918(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT58), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n737), .A2(new_n1063), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n728), .A2(new_n337), .B1(new_n740), .B2(new_n1059), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(new_n794), .C2(new_n1055), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n805), .B2(new_n742), .C1(new_n802), .C2(new_n732), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1124), .A2(KEYINPUT59), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n786), .A2(G159), .ZN(new_n1126));
  AOI21_X1  g0926(.A(G41), .B1(new_n749), .B2(G124), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1125), .A2(new_n254), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1124), .A2(KEYINPUT59), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1120), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n381), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n208), .B1(new_n1131), .B2(G41), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1119), .B2(KEYINPUT58), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT123), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n719), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n775), .B1(new_n208), .B2(new_n811), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1113), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1112), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1083), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1085), .B2(new_n1082), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1105), .A2(new_n1111), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT57), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1140), .A2(new_n1109), .A3(KEYINPUT57), .A4(new_n1110), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1144), .A2(new_n670), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1138), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(G375));
  AOI21_X1  g0947(.A(new_n977), .B1(G294), .B2(new_n792), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n515), .B2(new_n735), .C1(new_n475), .C2(new_n732), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n742), .A2(new_n561), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n737), .A2(new_n753), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n489), .B1(new_n210), .B2(new_n743), .C1(new_n758), .C2(new_n723), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1055), .A2(new_n968), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n727), .A2(G50), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n794), .A2(G159), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G137), .A2(new_n746), .B1(new_n786), .B2(G58), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n740), .A2(new_n805), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n732), .A2(new_n337), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n382), .B1(new_n1063), .B2(new_n723), .ZN(new_n1161));
  NOR4_X1   g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n719), .B1(new_n1153), .B2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n772), .B(new_n1163), .C1(new_n872), .C2(new_n715), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n229), .B2(new_n811), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1082), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n1049), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n922), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1169), .B2(new_n1084), .ZN(G381));
  INV_X1    g0970(.A(new_n1076), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1087), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(G375), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1174), .A2(G384), .A3(G381), .ZN(new_n1175));
  INV_X1    g0975(.A(G387), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1176), .A2(new_n1023), .A3(new_n1021), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1177), .A2(G396), .A3(G393), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1175), .A2(new_n1178), .ZN(G407));
  OAI211_X1 g0979(.A(G407), .B(G213), .C1(G343), .C2(new_n1174), .ZN(G409));
  NAND2_X1  g0980(.A1(G390), .A2(G387), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n1177), .ZN(new_n1182));
  XOR2_X1   g0982(.A(G393), .B(G396), .Z(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1181), .A2(new_n1177), .A3(new_n1183), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1168), .A2(KEYINPUT126), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT60), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1084), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT60), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1168), .A2(KEYINPUT126), .A3(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n670), .A3(new_n1190), .A4(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1167), .ZN(new_n1194));
  INV_X1    g0994(.A(G384), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT127), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1193), .A2(G384), .A3(new_n1167), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n645), .A2(G343), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(G2897), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1198), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G384), .B1(new_n1193), .B2(new_n1167), .ZN(new_n1204));
  OAI21_X1  g1004(.A(KEYINPUT127), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(new_n1201), .A3(new_n1199), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1202), .A2(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1141), .A2(new_n923), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1137), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1210), .B2(new_n1049), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1172), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1138), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(G378), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT125), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1146), .A2(KEYINPUT125), .A3(G378), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1212), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1207), .B1(new_n1219), .B2(new_n1200), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1219), .A2(new_n1200), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT62), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1220), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1212), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT125), .B1(new_n1146), .B2(G378), .ZN(new_n1227));
  AND4_X1   g1027(.A1(KEYINPUT125), .A2(new_n1213), .A3(G378), .A4(new_n1214), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1226), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1200), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n1224), .A3(new_n1230), .A4(new_n1221), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT61), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1187), .B1(new_n1225), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1229), .A2(new_n1230), .A3(new_n1221), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1229), .A2(new_n1230), .B1(new_n1202), .B2(new_n1206), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT63), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1229), .A2(KEYINPUT63), .A3(new_n1230), .A4(new_n1221), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT61), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1234), .A2(new_n1242), .ZN(G405));
  OAI22_X1  g1043(.A1(new_n1227), .A2(new_n1228), .B1(new_n1146), .B2(new_n1172), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(new_n1221), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(new_n1187), .ZN(G402));
endmodule


