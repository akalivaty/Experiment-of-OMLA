//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(G319));
  XNOR2_X1  g035(.A(KEYINPUT68), .B(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n464), .B(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n461), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n461), .A2(new_n462), .A3(G137), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT70), .B1(new_n477), .B2(new_n461), .ZN(new_n478));
  AND2_X1   g053(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n462), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n477), .A2(G2105), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n484), .A2(G124), .B1(G136), .B2(new_n485), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n461), .C2(G112), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n474), .B(new_n476), .C1(new_n479), .C2(new_n480), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT4), .A4(G138), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n474), .A2(new_n476), .A3(G126), .ZN(new_n497));
  NAND2_X1  g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n470), .A2(G102), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT71), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(new_n498), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n462), .B2(G126), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n503), .B(new_n500), .C1(new_n505), .C2(new_n496), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n495), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G62), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n516), .B1(KEYINPUT6), .B2(new_n513), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT72), .B(KEYINPUT6), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(new_n513), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(KEYINPUT72), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n516), .B(G651), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n512), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n515), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(G50), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n509), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G166));
  AOI21_X1  g108(.A(new_n509), .B1(new_n519), .B2(new_n524), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G51), .B1(G63), .B2(new_n514), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n512), .B1(new_n519), .B2(new_n524), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT75), .B(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT74), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n535), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(G168));
  AOI22_X1  g118(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n513), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n536), .A2(G90), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n534), .A2(G52), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n536), .A2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n534), .A2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n512), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT76), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n534), .A2(G43), .B1(G651), .B2(new_n554), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(new_n559), .A3(new_n550), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT77), .Z(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(new_n534), .A2(G53), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(KEYINPUT78), .B(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n512), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n536), .A2(G91), .B1(G651), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n534), .A2(KEYINPUT9), .A3(G53), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n571), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n571), .A2(new_n579), .A3(new_n575), .A4(new_n576), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n542), .B(new_n582), .ZN(G286));
  INV_X1    g158(.A(G166), .ZN(G303));
  OAI21_X1  g159(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT81), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n536), .A2(G87), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n534), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND3_X1  g164(.A1(new_n525), .A2(G48), .A3(G543), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n512), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n536), .A2(G86), .B1(G651), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n534), .A2(KEYINPUT82), .A3(G48), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n592), .A2(new_n596), .A3(KEYINPUT83), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n536), .A2(G85), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n534), .A2(G47), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n603), .B(new_n604), .C1(new_n513), .C2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT10), .B1(new_n527), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n512), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n534), .A2(G54), .B1(G651), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n536), .A2(new_n614), .A3(G92), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n609), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT84), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n609), .A2(new_n618), .A3(new_n613), .A4(new_n615), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n607), .B1(new_n620), .B2(G868), .ZN(G284));
  XOR2_X1   g196(.A(G284), .B(KEYINPUT85), .Z(G321));
  MUX2_X1   g197(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g198(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n620), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n620), .A2(new_n625), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT86), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(KEYINPUT87), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(KEYINPUT87), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n630), .B(new_n631), .C1(G868), .C2(new_n561), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n462), .A2(new_n470), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2100), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n485), .A2(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT88), .Z(new_n640));
  NOR2_X1   g215(.A1(new_n461), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(G123), .B2(new_n484), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2096), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n637), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2435), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2438), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n655), .B(new_n656), .Z(new_n657));
  AND2_X1   g232(.A1(new_n657), .A2(G14), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2067), .B(G2678), .Z(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT18), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT89), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT17), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n660), .B2(new_n661), .ZN(new_n670));
  AOI21_X1  g245(.A(KEYINPUT18), .B1(new_n662), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n668), .B(new_n671), .Z(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT90), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT20), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n682), .A2(new_n674), .A3(new_n677), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n680), .B(new_n683), .C1(new_n674), .C2(new_n682), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  INV_X1    g260(.A(G1981), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n684), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT91), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  NOR2_X1   g268(.A1(G16), .A2(G22), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G166), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT95), .B(G1971), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(G23), .B(G288), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT33), .B(G1976), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(G305), .A2(G16), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT32), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G6), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n703), .B1(new_n600), .B2(new_n601), .ZN(new_n706));
  INV_X1    g281(.A(new_n704), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT32), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n705), .A2(G1981), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(G1981), .B1(new_n705), .B2(new_n708), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n697), .B(new_n700), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n702), .B1(new_n701), .B2(new_n704), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n706), .A2(KEYINPUT32), .A3(new_n707), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n686), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n705), .A2(G1981), .A3(new_n708), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT34), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n717), .A2(new_n718), .A3(new_n700), .A4(new_n697), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(KEYINPUT96), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G25), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n484), .A2(G119), .B1(G131), .B2(new_n485), .ZN(new_n725));
  OAI221_X1 g300(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n461), .C2(G107), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n724), .B1(new_n727), .B2(new_n723), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT92), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT35), .B(G1991), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(G24), .B(G290), .S(G16), .Z(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT93), .B(G1986), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT94), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n732), .B(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n720), .A2(new_n722), .A3(new_n731), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n723), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT25), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(new_n461), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n485), .A2(G139), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n737), .B1(new_n743), .B2(new_n723), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(G2072), .Z(new_n745));
  NAND4_X1  g320(.A1(new_n712), .A2(new_n719), .A3(new_n731), .A4(new_n735), .ZN(new_n746));
  INV_X1    g321(.A(new_n722), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n721), .A2(KEYINPUT96), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(G299), .A2(G16), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n703), .A2(KEYINPUT23), .A3(G20), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT23), .ZN(new_n752));
  INV_X1    g327(.A(G20), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G16), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n750), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G1956), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n750), .A2(G1956), .A3(new_n751), .A4(new_n754), .ZN(new_n758));
  NOR2_X1   g333(.A1(G4), .A2(G16), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n617), .A2(new_n619), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(new_n703), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G1348), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n764), .B(new_n760), .C1(new_n761), .C2(new_n703), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n757), .A2(new_n758), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT26), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n484), .B2(G129), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n470), .A2(G105), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n485), .A2(G141), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G29), .B2(G32), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n703), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n703), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1961), .ZN(new_n781));
  NOR2_X1   g356(.A1(G29), .A2(G35), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G162), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT29), .B(G2090), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n723), .A2(G27), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G164), .B2(new_n723), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2078), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n781), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n766), .A2(new_n777), .A3(new_n778), .A4(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT31), .B(G11), .Z(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G34), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G29), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G160), .B2(G29), .ZN(new_n795));
  INV_X1    g370(.A(G2084), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n798), .A2(G28), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(G28), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n799), .A2(new_n800), .A3(G29), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n643), .B2(G29), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n723), .A2(G26), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n484), .A2(G128), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n485), .A2(G140), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n807));
  NOR2_X1   g382(.A1(G104), .A2(G2105), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT98), .Z(new_n809));
  OAI21_X1  g384(.A(new_n806), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n804), .B1(new_n811), .B2(new_n723), .ZN(new_n812));
  MUX2_X1   g387(.A(new_n804), .B(new_n812), .S(KEYINPUT28), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2067), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n790), .A2(new_n791), .A3(new_n803), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n736), .A2(new_n745), .A3(new_n749), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(G168), .A2(G16), .ZN(new_n817));
  INV_X1    g392(.A(G1966), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT100), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n817), .B(new_n819), .C1(G16), .C2(G21), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n818), .A2(KEYINPUT100), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n820), .B(new_n821), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n703), .A2(G19), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n561), .B2(new_n703), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT97), .Z(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(G1341), .Z(new_n826));
  NOR3_X1   g401(.A1(new_n816), .A2(new_n822), .A3(new_n826), .ZN(G311));
  OAI21_X1  g402(.A(new_n815), .B1(new_n747), .B2(new_n746), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n822), .ZN(new_n831));
  INV_X1    g406(.A(new_n826), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n745), .ZN(G150));
  NAND2_X1  g408(.A1(new_n536), .A2(G93), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n534), .A2(G55), .ZN(new_n835));
  NAND2_X1  g410(.A1(G80), .A2(G543), .ZN(new_n836));
  INV_X1    g411(.A(G67), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n512), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G651), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n834), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G860), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  INV_X1    g417(.A(new_n840), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n557), .B2(new_n560), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n840), .B1(new_n550), .B2(new_n558), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT39), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n620), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n847), .B(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n842), .B1(new_n850), .B2(G860), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT101), .ZN(G145));
  XNOR2_X1  g427(.A(new_n643), .B(G160), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n488), .ZN(new_n854));
  INV_X1    g429(.A(new_n727), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n484), .A2(G130), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT103), .ZN(new_n857));
  OAI221_X1 g432(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n461), .C2(G118), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n485), .A2(G142), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT102), .Z(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n635), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n861), .A2(new_n635), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n855), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n861), .A2(new_n635), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n727), .A3(new_n862), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n811), .A2(new_n772), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n811), .A2(new_n772), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n499), .A2(new_n501), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n493), .A3(new_n494), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  INV_X1    g451(.A(new_n872), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(new_n870), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n743), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n875), .A2(new_n878), .A3(new_n743), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n869), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n869), .A2(new_n883), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n854), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n865), .A2(new_n868), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n881), .A2(new_n865), .A3(new_n868), .A4(new_n882), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n888), .A2(new_n854), .A3(new_n889), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n886), .A2(new_n890), .A3(G37), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT40), .Z(G395));
  NOR2_X1   g467(.A1(new_n840), .A2(G868), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n628), .B(new_n846), .ZN(new_n894));
  INV_X1    g469(.A(new_n616), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(new_n578), .B2(new_n580), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n578), .A2(new_n580), .A3(new_n895), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  INV_X1    g475(.A(new_n898), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n901), .B2(new_n896), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n894), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n905));
  XNOR2_X1  g480(.A(G288), .B(G290), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(G305), .A2(G166), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n600), .A2(G303), .A3(new_n601), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n905), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n901), .A2(new_n896), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n894), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n904), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n915), .A2(new_n916), .A3(new_n905), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n921), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n923), .A2(new_n917), .A3(new_n904), .A4(new_n919), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n893), .B1(new_n925), .B2(G868), .ZN(G295));
  AOI21_X1  g501(.A(new_n893), .B1(new_n925), .B2(G868), .ZN(G331));
  OAI21_X1  g502(.A(KEYINPUT106), .B1(new_n844), .B2(new_n845), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n561), .A2(new_n840), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n930));
  INV_X1    g505(.A(new_n845), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n542), .B(KEYINPUT80), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n933), .A2(G301), .ZN(new_n934));
  NOR2_X1   g509(.A1(G171), .A2(new_n542), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n928), .B(new_n932), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(G286), .B2(G171), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n930), .B1(new_n929), .B2(new_n931), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n844), .A2(KEYINPUT106), .A3(new_n845), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n903), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n936), .A2(new_n940), .A3(new_n918), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n914), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G37), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n936), .A2(new_n940), .A3(new_n918), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n936), .A2(new_n940), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n913), .B(new_n945), .C1(new_n946), .C2(new_n903), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT108), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n951), .A3(KEYINPUT43), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT107), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n941), .B2(new_n942), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n954), .B(new_n945), .C1(new_n946), .C2(new_n903), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n944), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT44), .B1(new_n958), .B2(KEYINPUT43), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n943), .A2(new_n947), .A3(new_n961), .A4(new_n944), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI22_X1  g538(.A1(new_n953), .A2(new_n959), .B1(new_n963), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n493), .A2(new_n494), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n500), .B1(new_n505), .B2(new_n496), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n468), .A2(new_n471), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n463), .A2(new_n466), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n971), .B(G40), .C1(new_n461), .C2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n811), .B(G2067), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n772), .A2(G1996), .ZN(new_n976));
  INV_X1    g551(.A(G1996), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n773), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n730), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n727), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n727), .A2(new_n980), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n979), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G290), .A2(G1986), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(G290), .A2(G1986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n974), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT45), .B(new_n965), .C1(new_n966), .C2(new_n967), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT109), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n874), .A2(new_n991), .A3(KEYINPUT45), .A4(new_n965), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n502), .A2(new_n506), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n965), .B1(new_n994), .B2(new_n966), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n969), .ZN(new_n996));
  INV_X1    g571(.A(G40), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n467), .A2(new_n472), .A3(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT56), .B(G2072), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n993), .A2(new_n996), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n965), .C1(new_n994), .C2(new_n966), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n968), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n998), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n756), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1000), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n577), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n571), .A2(KEYINPUT57), .A3(new_n575), .A4(new_n576), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT120), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1000), .A2(new_n1006), .A3(new_n1011), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT61), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1007), .A2(KEYINPUT120), .A3(new_n1012), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n973), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n968), .A2(new_n1003), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1348), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1384), .B1(new_n495), .B2(new_n873), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(new_n998), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT119), .B1(new_n968), .B2(new_n973), .ZN(new_n1027));
  INV_X1    g602(.A(G2067), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NOR4_X1   g604(.A1(new_n1023), .A2(new_n1029), .A3(KEYINPUT60), .A4(new_n616), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n895), .B1(new_n1023), .B2(new_n1029), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1001), .B1(new_n507), .B2(new_n965), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1033), .A2(new_n973), .A3(new_n1021), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n616), .B(new_n1032), .C1(new_n1034), .C2(G1348), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1030), .B1(new_n1036), .B2(KEYINPUT60), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1011), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1015), .B1(new_n1038), .B2(KEYINPUT121), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1000), .A2(new_n1006), .A3(new_n1011), .A4(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(KEYINPUT61), .A3(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n993), .A2(new_n996), .A3(new_n977), .A4(new_n998), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT58), .B(G1341), .Z(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n561), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT59), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(new_n1050), .A3(new_n561), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1019), .A2(new_n1037), .A3(new_n1042), .A4(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1015), .B(new_n895), .C1(new_n1029), .C2(new_n1023), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1013), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT122), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n993), .A2(new_n996), .A3(new_n998), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT110), .B(G1971), .Z(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(G2090), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G8), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n1063));
  INV_X1    g638(.A(G8), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(G166), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT113), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1067), .B(new_n1063), .C1(G166), .C2(new_n1064), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT55), .B(G8), .C1(new_n529), .C2(new_n532), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1066), .B(new_n1068), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1062), .A2(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1005), .A2(KEYINPUT118), .ZN(new_n1076));
  INV_X1    g651(.A(G2090), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n1005), .B2(KEYINPUT118), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1059), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1073), .B1(new_n1079), .B2(G8), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1064), .B1(new_n1024), .B2(new_n998), .ZN(new_n1082));
  INV_X1    g657(.A(G1976), .ZN(new_n1083));
  NAND3_X1  g658(.A1(G288), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1082), .B(new_n1087), .C1(G288), .C2(new_n1083), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1086), .B(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n598), .A2(G1981), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n592), .A2(new_n596), .A3(new_n686), .A4(new_n597), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT49), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1091), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1097), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(new_n1100), .A3(new_n1082), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1098), .A2(new_n1100), .A3(KEYINPUT116), .A4(new_n1082), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1089), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1034), .A2(G1961), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1057), .A2(G2078), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n1108), .B(G2078), .C1(new_n968), .C2(new_n969), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n972), .B(KEYINPUT124), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n997), .B1(new_n1111), .B2(new_n481), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1110), .A2(new_n993), .A3(new_n971), .A4(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(G301), .B(KEYINPUT54), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1109), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1081), .A2(new_n1105), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n970), .B(new_n998), .C1(new_n995), .C2(new_n969), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n818), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1060), .B2(G2084), .ZN(new_n1123));
  OAI211_X1 g698(.A(G8), .B(new_n1120), .C1(new_n1123), .C2(new_n542), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1120), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n542), .A2(G8), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1034), .A2(new_n796), .B1(new_n1121), .B2(new_n818), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1125), .B(new_n1126), .C1(new_n1127), .C2(new_n1064), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1124), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1123), .A2(G8), .A3(new_n542), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1110), .B(new_n998), .C1(new_n969), .C2(new_n995), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1109), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n1114), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1117), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1053), .A2(new_n1138), .A3(new_n1054), .A4(new_n1013), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1056), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1081), .A2(new_n1105), .ZN(new_n1141));
  AOI21_X1  g716(.A(G301), .B1(new_n1109), .B2(new_n1133), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1132), .A2(KEYINPUT62), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1130), .A2(new_n1144), .A3(new_n1131), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1127), .A2(new_n1064), .A3(G286), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1062), .A2(new_n1074), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1105), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1151), .A2(new_n1080), .B1(new_n1062), .B2(new_n1074), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1149), .A2(KEYINPUT63), .B1(new_n1152), .B2(new_n1105), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1154));
  NOR2_X1   g729(.A1(G288), .A2(G1976), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(KEYINPUT117), .B(new_n1092), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT117), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1092), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(new_n1082), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1146), .A2(new_n1153), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n988), .B1(new_n1140), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n974), .A2(new_n977), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT46), .Z(new_n1166));
  INV_X1    g741(.A(new_n974), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n975), .B2(new_n773), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT47), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n974), .A2(new_n987), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT48), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n984), .B2(new_n1167), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n979), .A2(new_n974), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1174), .A2(new_n982), .B1(new_n1028), .B2(new_n811), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT125), .Z(new_n1176));
  OAI211_X1 g751(.A(new_n1170), .B(new_n1173), .C1(new_n1167), .C2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1164), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g755(.A(new_n891), .B1(new_n960), .B2(new_n962), .ZN(new_n1182));
  INV_X1    g756(.A(G227), .ZN(new_n1183));
  AOI21_X1  g757(.A(KEYINPUT127), .B1(G319), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g758(.A1(G401), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g759(.A1(G319), .A2(KEYINPUT127), .A3(new_n1183), .ZN(new_n1186));
  NAND4_X1  g760(.A1(new_n1182), .A2(new_n692), .A3(new_n1185), .A4(new_n1186), .ZN(G225));
  INV_X1    g761(.A(G225), .ZN(G308));
endmodule


