//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(G211gat), .A2(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207));
  AND2_X1   g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208));
  OAI22_X1  g007(.A1(new_n206), .A2(KEYINPUT22), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT70), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT71), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n209), .B1(new_n212), .B2(KEYINPUT69), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n209), .A2(KEYINPUT69), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(new_n214), .B2(KEYINPUT71), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G226gat), .ZN(new_n217));
  INV_X1    g016(.A(G233gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(KEYINPUT24), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n220), .A2(KEYINPUT24), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n221), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G169gat), .ZN(new_n227));
  INV_X1    g026(.A(G176gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT23), .ZN(new_n229));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n228), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n226), .A2(new_n229), .A3(new_n230), .A4(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n229), .A3(new_n230), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT25), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n237), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n231), .A2(KEYINPUT26), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n230), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n244), .B1(KEYINPUT26), .B2(new_n231), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n243), .A2(new_n245), .B1(G183gat), .B2(G190gat), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT27), .B1(new_n223), .B2(KEYINPUT65), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n223), .A2(KEYINPUT27), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n224), .B(new_n247), .C1(new_n248), .C2(KEYINPUT65), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT27), .B(G183gat), .Z(new_n252));
  NAND2_X1  g051(.A1(new_n224), .A2(KEYINPUT28), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n246), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n219), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n239), .A2(new_n238), .B1(new_n246), .B2(new_n254), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n259), .A2(new_n217), .A3(new_n218), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n216), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT73), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n219), .ZN(new_n263));
  INV_X1    g062(.A(new_n216), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n259), .A2(KEYINPUT29), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n263), .B(new_n264), .C1(new_n265), .C2(new_n219), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n261), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n262), .B1(new_n261), .B2(new_n266), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n205), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n261), .A2(new_n266), .A3(new_n204), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT75), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT30), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n270), .B2(new_n272), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n261), .A2(KEYINPUT30), .A3(new_n266), .A4(new_n204), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT74), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT40), .ZN(new_n280));
  NAND2_X1  g079(.A1(G225gat), .A2(G233gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(G141gat), .B(G148gat), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT2), .B1(new_n282), .B2(KEYINPUT77), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(KEYINPUT77), .B2(new_n282), .ZN(new_n284));
  INV_X1    g083(.A(G155gat), .ZN(new_n285));
  INV_X1    g084(.A(G162gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT76), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT76), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n282), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n290), .B1(new_n287), .B2(KEYINPUT2), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT4), .ZN(new_n298));
  XOR2_X1   g097(.A(G127gat), .B(G134gat), .Z(new_n299));
  XOR2_X1   g098(.A(G113gat), .B(G120gat), .Z(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(KEYINPUT68), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n301), .B(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n297), .A2(new_n298), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT79), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n296), .A3(new_n293), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT4), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT79), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n297), .A2(new_n309), .A3(new_n298), .A4(new_n304), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n304), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT3), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n293), .A2(new_n296), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n293), .A2(KEYINPUT78), .A3(new_n296), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n312), .B(new_n314), .C1(new_n319), .C2(new_n313), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n281), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT39), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT0), .ZN(new_n325));
  XNOR2_X1  g124(.A(G57gat), .B(G85gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n325), .B(new_n326), .Z(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n317), .A2(new_n318), .A3(new_n312), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n307), .ZN(new_n330));
  INV_X1    g129(.A(new_n281), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT39), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n321), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n280), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n327), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n321), .B2(new_n322), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n336), .B(KEYINPUT40), .C1(new_n321), .C2(new_n332), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n331), .B1(new_n308), .B2(new_n305), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n320), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT5), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n330), .B2(new_n331), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n311), .A2(new_n320), .A3(new_n340), .A4(new_n281), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT83), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n335), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n343), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(KEYINPUT83), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n334), .B(new_n337), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT84), .B1(new_n279), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n270), .A2(new_n272), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT75), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n276), .B(KEYINPUT74), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n269), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n328), .A2(new_n333), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n344), .A2(new_n345), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n327), .B1(new_n347), .B2(KEYINPUT83), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n357), .A2(KEYINPUT40), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n356), .A2(new_n360), .A3(new_n361), .A4(new_n334), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n264), .B1(new_n258), .B2(new_n260), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n263), .B(new_n216), .C1(new_n265), .C2(new_n219), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(KEYINPUT37), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT37), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n261), .A2(new_n366), .A3(new_n266), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT85), .B(KEYINPUT38), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n365), .A2(new_n367), .A3(new_n205), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n270), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT37), .B1(new_n267), .B2(new_n268), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n367), .A2(new_n205), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n368), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n327), .B1(new_n342), .B2(new_n343), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT6), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n376), .B2(KEYINPUT6), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT6), .B1(new_n344), .B2(new_n327), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(new_n346), .B2(new_n348), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n375), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n385));
  INV_X1    g184(.A(G228gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(new_n218), .ZN(new_n387));
  INV_X1    g186(.A(new_n257), .ZN(new_n388));
  INV_X1    g187(.A(new_n211), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(new_n209), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n389), .B2(new_n209), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n313), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n315), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n315), .A2(KEYINPUT3), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n216), .B1(new_n394), .B2(new_n388), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n387), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n387), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n213), .A2(new_n399), .A3(new_n215), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n319), .B1(new_n313), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n397), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n313), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n317), .A3(new_n318), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n404), .A2(KEYINPUT81), .A3(new_n387), .A4(new_n395), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n396), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G22gat), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n385), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT31), .B(G50gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n406), .A2(new_n407), .ZN(new_n413));
  AOI211_X1 g212(.A(G22gat), .B(new_n396), .C1(new_n402), .C2(new_n405), .ZN(new_n414));
  OAI22_X1  g213(.A1(new_n408), .A2(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n402), .A2(new_n405), .ZN(new_n416));
  OAI21_X1  g215(.A(G22gat), .B1(new_n416), .B2(new_n396), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n406), .A2(new_n407), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n417), .A2(new_n385), .A3(new_n418), .A4(new_n411), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n350), .A2(new_n362), .A3(new_n384), .A4(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n376), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n382), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n380), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n378), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n279), .ZN(new_n426));
  INV_X1    g225(.A(new_n420), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n256), .A2(new_n304), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n259), .A2(new_n312), .ZN(new_n429));
  INV_X1    g228(.A(G227gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(new_n218), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT32), .ZN(new_n433));
  XOR2_X1   g232(.A(G15gat), .B(G43gat), .Z(new_n434));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT34), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n428), .A2(new_n429), .ZN(new_n441));
  INV_X1    g240(.A(new_n431), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI211_X1 g242(.A(KEYINPUT34), .B(new_n431), .C1(new_n428), .C2(new_n429), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n439), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n439), .A2(new_n443), .A3(new_n444), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n433), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OR3_X1    g247(.A1(new_n439), .A2(new_n443), .A3(new_n444), .ZN(new_n449));
  INV_X1    g248(.A(new_n433), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n445), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT36), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n451), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT36), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n426), .A2(new_n427), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n420), .A2(new_n425), .A3(new_n279), .A4(new_n452), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT35), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n454), .B1(new_n419), .B2(new_n415), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT35), .B1(new_n381), .B2(new_n383), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n279), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n421), .A2(new_n457), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT15), .ZN(new_n465));
  XNOR2_X1  g264(.A(G43gat), .B(G50gat), .ZN(new_n466));
  INV_X1    g265(.A(G36gat), .ZN(new_n467));
  AND2_X1   g266(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G29gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n472));
  AOI211_X1 g271(.A(new_n465), .B(new_n466), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n465), .A3(new_n472), .ZN(new_n474));
  INV_X1    g273(.A(new_n466), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n470), .A2(new_n472), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(KEYINPUT15), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n479));
  INV_X1    g278(.A(G8gat), .ZN(new_n480));
  INV_X1    g279(.A(G15gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G22gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n407), .A2(G15gat), .ZN(new_n483));
  INV_X1    g282(.A(G1gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT16), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(G1gat), .B1(new_n482), .B2(new_n483), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n479), .B(new_n480), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n482), .A2(new_n483), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n484), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n479), .A2(new_n480), .ZN(new_n492));
  NAND2_X1  g291(.A1(KEYINPUT87), .A2(G8gat), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n464), .B1(new_n478), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT14), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n471), .ZN(new_n498));
  NAND2_X1  g297(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n499));
  AOI21_X1  g298(.A(G36gat), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n472), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT15), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(new_n474), .A3(new_n466), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n476), .A2(KEYINPUT15), .A3(new_n475), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n488), .A2(new_n494), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT88), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n496), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G229gat), .A2(G233gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n503), .A2(new_n510), .A3(new_n504), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n503), .B2(new_n504), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n495), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n508), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT18), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT88), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT88), .B1(new_n505), .B2(new_n506), .ZN(new_n518));
  OAI22_X1  g317(.A1(new_n517), .A2(new_n518), .B1(new_n506), .B2(new_n505), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n509), .B(KEYINPUT13), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n508), .A2(KEYINPUT18), .A3(new_n509), .A4(new_n513), .ZN(new_n522));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(G169gat), .B(G197gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT12), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n516), .A2(new_n521), .A3(new_n522), .A4(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n528), .B1(new_n514), .B2(new_n515), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(KEYINPUT90), .A3(new_n521), .A4(new_n522), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT89), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n522), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n516), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n536), .B1(new_n521), .B2(new_n522), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n528), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT21), .ZN(new_n543));
  XNOR2_X1  g342(.A(G57gat), .B(G64gat), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n547), .B(new_n546), .C1(new_n544), .C2(new_n549), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n495), .B1(new_n543), .B2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT92), .Z(new_n555));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT91), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n555), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n553), .A2(new_n543), .ZN(new_n561));
  XOR2_X1   g360(.A(G127gat), .B(G155gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G99gat), .B(G106gat), .Z(new_n569));
  NAND2_X1  g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT8), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(G99gat), .B2(G106gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(G85gat), .A2(G92gat), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT93), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT8), .ZN(new_n580));
  OR2_X1    g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI211_X1 g382(.A(new_n569), .B(new_n574), .C1(new_n578), .C2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n569), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n578), .A2(new_n583), .ZN(new_n586));
  INV_X1    g385(.A(new_n574), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI22_X1  g387(.A1(new_n511), .A2(new_n512), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n584), .ZN(new_n590));
  AND2_X1   g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n590), .A2(new_n505), .B1(KEYINPUT41), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT94), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n593), .A2(new_n595), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n599));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n598), .A2(new_n601), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n568), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G120gat), .B(G148gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n553), .B1(new_n588), .B2(new_n584), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n580), .A2(new_n582), .A3(new_n581), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n582), .B1(new_n580), .B2(new_n581), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n587), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n569), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n551), .A2(new_n552), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n586), .A2(new_n585), .A3(new_n587), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n610), .A2(new_n611), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n610), .B2(new_n618), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n609), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n625), .A2(KEYINPUT95), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(KEYINPUT95), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n623), .A2(new_n627), .A3(new_n608), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NOR4_X1   g429(.A1(new_n463), .A2(new_n542), .A3(new_n605), .A4(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n631), .A2(KEYINPUT96), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(KEYINPUT96), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n425), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g436(.A(KEYINPUT16), .B(G8gat), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI211_X1 g438(.A(new_n279), .B(new_n639), .C1(new_n632), .C2(new_n633), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n640), .A2(KEYINPUT42), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n480), .B1(new_n634), .B2(new_n356), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT42), .B1(new_n642), .B2(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(G1325gat));
  NAND3_X1  g443(.A1(new_n634), .A2(new_n481), .A3(new_n452), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n453), .A2(new_n456), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n634), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n647), .B2(new_n481), .ZN(G1326gat));
  NAND2_X1  g447(.A1(new_n634), .A2(new_n427), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT97), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n651), .A3(new_n427), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT43), .B(G22gat), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n651), .B1(new_n634), .B2(new_n427), .ZN(new_n656));
  AOI211_X1 g455(.A(KEYINPUT97), .B(new_n420), .C1(new_n632), .C2(new_n633), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(G1327gat));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n604), .A2(KEYINPUT101), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n602), .B2(new_n603), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT100), .B(KEYINPUT44), .Z(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n660), .B1(new_n463), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT44), .B1(new_n463), .B2(new_n604), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n421), .A2(new_n457), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n420), .A2(new_n452), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n356), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n673), .A2(new_n461), .B1(new_n458), .B2(KEYINPUT35), .ZN(new_n674));
  OAI211_X1 g473(.A(KEYINPUT102), .B(new_n667), .C1(new_n671), .C2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n669), .A2(new_n670), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n535), .A2(new_n677), .A3(new_n540), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n535), .B2(new_n540), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n568), .ZN(new_n682));
  INV_X1    g481(.A(new_n630), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT99), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n676), .A2(new_n635), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n471), .B1(new_n687), .B2(KEYINPUT103), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(KEYINPUT103), .B2(new_n687), .ZN(new_n689));
  NOR4_X1   g488(.A1(new_n463), .A2(new_n542), .A3(new_n604), .A4(new_n684), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n471), .A3(new_n635), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT45), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(G1328gat));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n694));
  AOI21_X1  g493(.A(G36gat), .B1(new_n694), .B2(KEYINPUT46), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n690), .A2(new_n356), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n694), .A2(KEYINPUT46), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n676), .A2(new_n356), .A3(new_n686), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n467), .B2(new_n699), .ZN(G1329gat));
  NAND3_X1  g499(.A1(new_n676), .A2(new_n646), .A3(new_n686), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n676), .A2(KEYINPUT106), .A3(new_n646), .A4(new_n686), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(G43gat), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n454), .A2(G43gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n705), .A2(KEYINPUT47), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n701), .A2(G43gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n707), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n709), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n701), .A2(G43gat), .B1(new_n690), .B2(new_n706), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(KEYINPUT105), .A3(KEYINPUT47), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n708), .B1(new_n713), .B2(new_n715), .ZN(G1330gat));
  NAND4_X1  g515(.A1(new_n676), .A2(G50gat), .A3(new_n427), .A4(new_n686), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n690), .A2(new_n427), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(G50gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g519(.A1(new_n680), .A2(new_n605), .A3(new_n683), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT107), .Z(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n463), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n635), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G57gat), .ZN(G1332gat));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n726));
  INV_X1    g525(.A(G64gat), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n723), .B(new_n356), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1333gat));
  INV_X1    g529(.A(G71gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n723), .A2(new_n731), .A3(new_n452), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n723), .A2(new_n646), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(new_n731), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g534(.A1(new_n723), .A2(new_n427), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g536(.A1(new_n680), .A2(new_n568), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n630), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n676), .A2(new_n635), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(G85gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n463), .A2(new_n604), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n743), .A2(KEYINPUT51), .A3(new_n738), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT51), .B1(new_n743), .B2(new_n738), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n630), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n635), .A2(new_n742), .ZN(new_n747));
  OAI22_X1  g546(.A1(new_n741), .A2(new_n742), .B1(new_n746), .B2(new_n747), .ZN(G1336gat));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n279), .A2(G92gat), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n630), .B(new_n750), .C1(new_n744), .C2(new_n745), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n676), .A2(new_n356), .A3(new_n740), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n753), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n749), .B(new_n751), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n752), .A2(G92gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n751), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT52), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(G1337gat));
  NAND3_X1  g560(.A1(new_n676), .A2(new_n646), .A3(new_n740), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G99gat), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n454), .A2(G99gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n746), .B2(new_n764), .ZN(G1338gat));
  NAND3_X1  g564(.A1(new_n676), .A2(new_n427), .A3(new_n740), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G106gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n420), .A2(G106gat), .A3(new_n683), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT109), .Z(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n744), .B2(new_n745), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n621), .B2(new_n622), .ZN(new_n776));
  INV_X1    g575(.A(new_n622), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n619), .A2(new_n777), .A3(new_n620), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n774), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  AOI211_X1 g578(.A(KEYINPUT54), .B(new_n777), .C1(new_n619), .C2(new_n620), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n780), .A2(KEYINPUT110), .A3(new_n608), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n621), .A2(new_n775), .A3(new_n622), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n609), .ZN(new_n784));
  OAI211_X1 g583(.A(KEYINPUT111), .B(new_n779), .C1(new_n781), .C2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT110), .B1(new_n780), .B2(new_n608), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n782), .A3(new_n609), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT111), .B1(new_n789), .B2(new_n779), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n787), .A2(new_n788), .B1(new_n778), .B2(new_n776), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n629), .B1(new_n792), .B2(KEYINPUT55), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n773), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n789), .A2(new_n779), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n785), .ZN(new_n798));
  INV_X1    g597(.A(new_n629), .ZN(new_n799));
  INV_X1    g598(.A(new_n792), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(new_n774), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n801), .A3(KEYINPUT112), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n680), .A2(new_n794), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n519), .A2(new_n520), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n509), .B1(new_n508), .B2(new_n513), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n527), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT113), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n535), .A3(new_n630), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n664), .B1(new_n803), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n808), .A2(new_n535), .ZN(new_n811));
  AND4_X1   g610(.A1(new_n664), .A2(new_n794), .A3(new_n802), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n682), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n605), .A2(new_n630), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n681), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n425), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n673), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n680), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n427), .B1(new_n813), .B2(new_n815), .ZN(new_n820));
  AND4_X1   g619(.A1(new_n635), .A2(new_n820), .A3(new_n279), .A4(new_n452), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n541), .A2(G113gat), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(G1340gat));
  AOI21_X1  g622(.A(G120gat), .B1(new_n818), .B2(new_n630), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n630), .A2(G120gat), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n821), .B2(new_n825), .ZN(G1341gat));
  NOR3_X1   g625(.A1(new_n817), .A2(G127gat), .A3(new_n682), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n821), .A2(new_n568), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(G127gat), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT114), .ZN(G1342gat));
  INV_X1    g629(.A(new_n604), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n821), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G134gat), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n356), .A2(new_n604), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT115), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(G134gat), .A3(new_n672), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n816), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g636(.A(new_n837), .B(KEYINPUT56), .Z(new_n838));
  NAND2_X1  g637(.A1(new_n833), .A2(new_n838), .ZN(G1343gat));
  NAND3_X1  g638(.A1(new_n798), .A2(new_n801), .A3(new_n541), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n831), .B1(new_n840), .B2(new_n809), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n682), .B1(new_n812), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n815), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(KEYINPUT57), .A3(new_n427), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n420), .B1(new_n813), .B2(new_n815), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(KEYINPUT57), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n646), .A2(new_n425), .A3(new_n356), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G141gat), .B1(new_n848), .B2(new_n681), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n646), .A2(new_n420), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n542), .A2(G141gat), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n816), .A2(new_n279), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT58), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(G141gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n813), .A2(new_n815), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT57), .B1(new_n859), .B2(new_n427), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n843), .A2(KEYINPUT57), .A3(new_n427), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n541), .B(new_n847), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n858), .B1(new_n862), .B2(KEYINPUT116), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n846), .A2(new_n864), .A3(new_n541), .A4(new_n847), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n855), .B(new_n857), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n862), .A2(KEYINPUT116), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(G141gat), .A3(new_n865), .ZN(new_n868));
  INV_X1    g667(.A(new_n857), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT117), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n854), .B1(new_n866), .B2(new_n870), .ZN(G1344gat));
  INV_X1    g670(.A(G148gat), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(KEYINPUT59), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n873), .B1(new_n848), .B2(new_n683), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(KEYINPUT118), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(KEYINPUT118), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n845), .A2(KEYINPUT57), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879));
  AND4_X1   g678(.A1(new_n831), .A2(new_n811), .A3(new_n798), .A4(new_n801), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n682), .B1(new_n880), .B2(new_n841), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n814), .A2(new_n542), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n420), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n879), .B1(new_n883), .B2(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n845), .A2(new_n879), .A3(KEYINPUT57), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n847), .A2(new_n630), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n872), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI22_X1  g688(.A1(new_n875), .A2(new_n876), .B1(new_n877), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n816), .A2(new_n850), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(new_n279), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n872), .A3(new_n630), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(G1345gat));
  NAND3_X1  g693(.A1(new_n892), .A2(new_n285), .A3(new_n568), .ZN(new_n895));
  OAI21_X1  g694(.A(G155gat), .B1(new_n848), .B2(new_n682), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n897), .B(new_n898), .ZN(G1346gat));
  NOR2_X1   g698(.A1(new_n835), .A2(G162gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n891), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT121), .Z(new_n902));
  OAI21_X1  g701(.A(G162gat), .B1(new_n848), .B2(new_n665), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n635), .A2(new_n279), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n454), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n820), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(new_n227), .A3(new_n542), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT122), .B1(new_n859), .B2(new_n425), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  AOI211_X1 g710(.A(new_n911), .B(new_n635), .C1(new_n813), .C2(new_n815), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n460), .A2(new_n356), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT123), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n913), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n917), .A2(new_n680), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n909), .B1(new_n920), .B2(new_n227), .ZN(G1348gat));
  OAI21_X1  g720(.A(G176gat), .B1(new_n908), .B2(new_n683), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n917), .A2(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n630), .A2(new_n228), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(G1349gat));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(KEYINPUT60), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n682), .A2(new_n252), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n915), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G183gat), .B1(new_n908), .B2(new_n682), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n926), .A2(KEYINPUT60), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT125), .Z(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n931), .B(new_n934), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n908), .B2(new_n604), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n664), .A2(new_n224), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n923), .B2(new_n938), .ZN(G1351gat));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n906), .A2(new_n646), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n887), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n940), .B1(new_n942), .B2(new_n542), .ZN(new_n943));
  INV_X1    g742(.A(new_n941), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n944), .B1(new_n885), .B2(new_n886), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(KEYINPUT126), .A3(new_n541), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n943), .A2(G197gat), .A3(new_n946), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n646), .A2(new_n279), .A3(new_n420), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n913), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n681), .A2(G197gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1352gat));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n683), .A2(G204gat), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n948), .B(new_n953), .C1(new_n910), .C2(new_n912), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT62), .ZN(new_n955));
  INV_X1    g754(.A(G204gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n956), .B1(new_n945), .B2(new_n630), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n952), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n942), .B2(new_n683), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n954), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n961), .A3(KEYINPUT127), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n958), .A2(new_n962), .ZN(G1353gat));
  OR3_X1    g762(.A1(new_n949), .A2(G211gat), .A3(new_n682), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n945), .A2(new_n568), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  OAI21_X1  g767(.A(G218gat), .B1(new_n942), .B2(new_n604), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n665), .A2(G218gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n949), .B2(new_n970), .ZN(G1355gat));
endmodule


