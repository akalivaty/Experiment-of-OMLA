

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593;

  XNOR2_X1 U324 ( .A(n404), .B(n403), .ZN(n405) );
  NOR2_X1 U325 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U326 ( .A(KEYINPUT124), .B(n457), .ZN(n574) );
  XNOR2_X1 U327 ( .A(n387), .B(n585), .ZN(n556) );
  XOR2_X1 U328 ( .A(G92GAT), .B(G218GAT), .Z(n292) );
  AND2_X1 U329 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U330 ( .A(G50GAT), .B(n509), .Z(n294) );
  NOR2_X1 U331 ( .A1(n589), .A2(n389), .ZN(n390) );
  XNOR2_X1 U332 ( .A(G71GAT), .B(G57GAT), .ZN(n337) );
  XNOR2_X1 U333 ( .A(n414), .B(n353), .ZN(n354) );
  OR2_X1 U334 ( .A1(n537), .A2(n529), .ZN(n477) );
  INV_X1 U335 ( .A(KEYINPUT95), .ZN(n403) );
  XNOR2_X1 U336 ( .A(n375), .B(n293), .ZN(n376) );
  AND2_X1 U337 ( .A1(n577), .A2(n454), .ZN(n455) );
  NOR2_X1 U338 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U339 ( .A(n377), .B(n376), .ZN(n381) );
  XNOR2_X1 U340 ( .A(n406), .B(n405), .ZN(n409) );
  AND2_X1 U341 ( .A1(n497), .A2(n522), .ZN(n498) );
  NOR2_X1 U342 ( .A1(n541), .A2(n456), .ZN(n457) );
  XNOR2_X1 U343 ( .A(n383), .B(n382), .ZN(n585) );
  INV_X1 U344 ( .A(G190GAT), .ZN(n459) );
  XNOR2_X1 U345 ( .A(n411), .B(n410), .ZN(n527) );
  XNOR2_X1 U346 ( .A(KEYINPUT38), .B(n499), .ZN(n508) );
  XNOR2_X1 U347 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U348 ( .A(n462), .B(n461), .ZN(G1351GAT) );
  XOR2_X1 U349 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n296) );
  XNOR2_X1 U350 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U352 ( .A(G169GAT), .B(n297), .Z(n400) );
  XOR2_X1 U353 ( .A(KEYINPUT80), .B(G134GAT), .Z(n299) );
  XNOR2_X1 U354 ( .A(G127GAT), .B(G120GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U356 ( .A(KEYINPUT0), .B(n300), .ZN(n452) );
  XOR2_X1 U357 ( .A(n400), .B(n452), .Z(n313) );
  XOR2_X1 U358 ( .A(G190GAT), .B(G99GAT), .Z(n302) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(G15GAT), .ZN(n301) );
  XNOR2_X1 U360 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U361 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n304) );
  XNOR2_X1 U362 ( .A(G71GAT), .B(KEYINPUT83), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U364 ( .A(n306), .B(n305), .Z(n311) );
  XOR2_X1 U365 ( .A(G183GAT), .B(G176GAT), .Z(n308) );
  NAND2_X1 U366 ( .A1(G227GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U368 ( .A(G113GAT), .B(n309), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n541) );
  XNOR2_X1 U371 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n314), .B(G29GAT), .ZN(n315) );
  XOR2_X1 U373 ( .A(n315), .B(KEYINPUT69), .Z(n317) );
  XNOR2_X1 U374 ( .A(KEYINPUT68), .B(KEYINPUT7), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n351) );
  XOR2_X1 U376 ( .A(G8GAT), .B(G15GAT), .Z(n319) );
  XNOR2_X1 U377 ( .A(G169GAT), .B(G197GAT), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n351), .B(n320), .ZN(n330) );
  XOR2_X1 U380 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n322) );
  XNOR2_X1 U381 ( .A(KEYINPUT67), .B(KEYINPUT66), .ZN(n321) );
  XOR2_X1 U382 ( .A(n322), .B(n321), .Z(n326) );
  XOR2_X1 U383 ( .A(G36GAT), .B(G50GAT), .Z(n324) );
  XOR2_X1 U384 ( .A(G141GAT), .B(G22GAT), .Z(n415) );
  XOR2_X1 U385 ( .A(G113GAT), .B(G1GAT), .Z(n436) );
  XNOR2_X1 U386 ( .A(n415), .B(n436), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n326), .B(n325), .ZN(n328) );
  NAND2_X1 U389 ( .A1(G229GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n580) );
  XOR2_X1 U392 ( .A(G8GAT), .B(G183GAT), .Z(n402) );
  XOR2_X1 U393 ( .A(G155GAT), .B(G78GAT), .Z(n332) );
  XNOR2_X1 U394 ( .A(G22GAT), .B(G211GAT), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U396 ( .A(n402), .B(n333), .Z(n335) );
  NAND2_X1 U397 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U399 ( .A(n336), .B(KEYINPUT79), .Z(n339) );
  XNOR2_X1 U400 ( .A(n337), .B(KEYINPUT13), .ZN(n369) );
  XNOR2_X1 U401 ( .A(n369), .B(KEYINPUT78), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n347) );
  XOR2_X1 U403 ( .A(G64GAT), .B(G127GAT), .Z(n341) );
  XNOR2_X1 U404 ( .A(G15GAT), .B(G1GAT), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U406 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n343) );
  XNOR2_X1 U407 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U409 ( .A(n345), .B(n344), .Z(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n589) );
  INV_X1 U411 ( .A(n589), .ZN(n561) );
  XOR2_X1 U412 ( .A(KEYINPUT10), .B(KEYINPUT74), .Z(n349) );
  XNOR2_X1 U413 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n361) );
  XNOR2_X1 U416 ( .A(G36GAT), .B(G190GAT), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n292), .B(n352), .ZN(n401) );
  XOR2_X1 U418 ( .A(G50GAT), .B(G162GAT), .Z(n414) );
  AND2_X1 U419 ( .A1(G232GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n401), .B(n354), .ZN(n355) );
  XOR2_X1 U421 ( .A(n355), .B(KEYINPUT75), .Z(n359) );
  XOR2_X1 U422 ( .A(KEYINPUT71), .B(G85GAT), .Z(n357) );
  XNOR2_X1 U423 ( .A(G99GAT), .B(G106GAT), .ZN(n356) );
  XNOR2_X1 U424 ( .A(n357), .B(n356), .ZN(n379) );
  XNOR2_X1 U425 ( .A(n379), .B(KEYINPUT9), .ZN(n358) );
  XNOR2_X1 U426 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n564) );
  XNOR2_X1 U428 ( .A(n564), .B(KEYINPUT76), .ZN(n458) );
  INV_X1 U429 ( .A(KEYINPUT36), .ZN(n362) );
  XNOR2_X1 U430 ( .A(n458), .B(n362), .ZN(n492) );
  NOR2_X1 U431 ( .A1(n561), .A2(n492), .ZN(n365) );
  XOR2_X1 U432 ( .A(KEYINPUT117), .B(KEYINPUT45), .Z(n363) );
  XNOR2_X1 U433 ( .A(KEYINPUT64), .B(n363), .ZN(n364) );
  XNOR2_X1 U434 ( .A(n365), .B(n364), .ZN(n384) );
  XOR2_X1 U435 ( .A(KEYINPUT32), .B(G92GAT), .Z(n367) );
  XNOR2_X1 U436 ( .A(G120GAT), .B(G204GAT), .ZN(n366) );
  XOR2_X1 U437 ( .A(n367), .B(n366), .Z(n383) );
  XOR2_X1 U438 ( .A(G176GAT), .B(G64GAT), .Z(n407) );
  INV_X1 U439 ( .A(n407), .ZN(n368) );
  NAND2_X1 U440 ( .A1(n369), .A2(n368), .ZN(n372) );
  INV_X1 U441 ( .A(n369), .ZN(n370) );
  NAND2_X1 U442 ( .A1(n370), .A2(n407), .ZN(n371) );
  NAND2_X1 U443 ( .A1(n372), .A2(n371), .ZN(n377) );
  XOR2_X1 U444 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n374) );
  XNOR2_X1 U445 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n373) );
  XNOR2_X1 U446 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U447 ( .A(G78GAT), .B(KEYINPUT70), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n378), .B(G148GAT), .ZN(n426) );
  XNOR2_X1 U449 ( .A(n426), .B(n379), .ZN(n380) );
  XNOR2_X1 U450 ( .A(n381), .B(n380), .ZN(n382) );
  NAND2_X1 U451 ( .A1(n384), .A2(n585), .ZN(n385) );
  NOR2_X1 U452 ( .A1(n580), .A2(n385), .ZN(n386) );
  XNOR2_X1 U453 ( .A(KEYINPUT118), .B(n386), .ZN(n395) );
  INV_X1 U454 ( .A(KEYINPUT116), .ZN(n391) );
  INV_X1 U455 ( .A(KEYINPUT41), .ZN(n387) );
  INV_X1 U456 ( .A(n580), .ZN(n553) );
  NOR2_X1 U457 ( .A1(n556), .A2(n553), .ZN(n388) );
  XNOR2_X1 U458 ( .A(n388), .B(KEYINPUT46), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n391), .B(n390), .ZN(n392) );
  NOR2_X1 U460 ( .A1(n564), .A2(n392), .ZN(n393) );
  XOR2_X1 U461 ( .A(KEYINPUT47), .B(n393), .Z(n394) );
  XNOR2_X1 U462 ( .A(n396), .B(KEYINPUT48), .ZN(n538) );
  XOR2_X1 U463 ( .A(KEYINPUT21), .B(G211GAT), .Z(n398) );
  XNOR2_X1 U464 ( .A(KEYINPUT84), .B(G204GAT), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U466 ( .A(G197GAT), .B(n399), .Z(n434) );
  XNOR2_X1 U467 ( .A(n400), .B(n434), .ZN(n411) );
  XOR2_X1 U468 ( .A(n402), .B(n401), .Z(n406) );
  NAND2_X1 U469 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n407), .B(KEYINPUT94), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n527), .B(KEYINPUT123), .ZN(n412) );
  NOR2_X1 U473 ( .A1(n538), .A2(n412), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n413), .B(KEYINPUT54), .ZN(n577) );
  XOR2_X1 U475 ( .A(G106GAT), .B(G218GAT), .Z(n417) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U477 ( .A(n417), .B(n416), .ZN(n430) );
  XOR2_X1 U478 ( .A(KEYINPUT22), .B(KEYINPUT90), .Z(n419) );
  XNOR2_X1 U479 ( .A(KEYINPUT88), .B(KEYINPUT24), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U481 ( .A(KEYINPUT89), .B(KEYINPUT86), .Z(n421) );
  XNOR2_X1 U482 ( .A(KEYINPUT23), .B(KEYINPUT87), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U484 ( .A(n423), .B(n422), .Z(n428) );
  XOR2_X1 U485 ( .A(G155GAT), .B(KEYINPUT2), .Z(n425) );
  XNOR2_X1 U486 ( .A(KEYINPUT3), .B(KEYINPUT85), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n426), .B(n435), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U490 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U493 ( .A(n434), .B(n433), .Z(n473) );
  XOR2_X1 U494 ( .A(G162GAT), .B(n435), .Z(n438) );
  XNOR2_X1 U495 ( .A(G29GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n451) );
  XOR2_X1 U497 ( .A(KEYINPUT1), .B(G85GAT), .Z(n440) );
  XNOR2_X1 U498 ( .A(G141GAT), .B(G148GAT), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U500 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n442) );
  XNOR2_X1 U501 ( .A(G57GAT), .B(KEYINPUT6), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U503 ( .A(n444), .B(n443), .Z(n449) );
  XOR2_X1 U504 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n446) );
  NAND2_X1 U505 ( .A1(G225GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U506 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U507 ( .A(KEYINPUT91), .B(n447), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n576) );
  INV_X1 U511 ( .A(n576), .ZN(n525) );
  NOR2_X1 U512 ( .A1(n473), .A2(n525), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n455), .B(KEYINPUT55), .ZN(n456) );
  NAND2_X1 U514 ( .A1(n574), .A2(n458), .ZN(n462) );
  XOR2_X1 U515 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n460) );
  AND2_X1 U516 ( .A1(n580), .A2(n585), .ZN(n497) );
  INV_X1 U517 ( .A(n541), .ZN(n529) );
  NAND2_X1 U518 ( .A1(n527), .A2(n529), .ZN(n463) );
  XOR2_X1 U519 ( .A(KEYINPUT98), .B(n463), .Z(n464) );
  NOR2_X1 U520 ( .A1(n473), .A2(n464), .ZN(n466) );
  XNOR2_X1 U521 ( .A(KEYINPUT25), .B(KEYINPUT99), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(n470) );
  NAND2_X1 U523 ( .A1(n473), .A2(n541), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n467), .B(KEYINPUT26), .ZN(n579) );
  XOR2_X1 U525 ( .A(n527), .B(KEYINPUT96), .Z(n468) );
  XNOR2_X1 U526 ( .A(KEYINPUT27), .B(n468), .ZN(n475) );
  NOR2_X1 U527 ( .A1(n579), .A2(n475), .ZN(n469) );
  NOR2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n525), .A2(n471), .ZN(n472) );
  XNOR2_X1 U530 ( .A(KEYINPUT100), .B(n472), .ZN(n479) );
  XOR2_X1 U531 ( .A(n473), .B(KEYINPUT28), .Z(n474) );
  XNOR2_X1 U532 ( .A(KEYINPUT65), .B(n474), .ZN(n532) );
  NOR2_X1 U533 ( .A1(n576), .A2(n475), .ZN(n476) );
  XNOR2_X1 U534 ( .A(KEYINPUT97), .B(n476), .ZN(n537) );
  NOR2_X1 U535 ( .A1(n532), .A2(n477), .ZN(n478) );
  NOR2_X1 U536 ( .A1(n479), .A2(n478), .ZN(n493) );
  NOR2_X1 U537 ( .A1(n561), .A2(n458), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n480), .Z(n481) );
  NOR2_X1 U539 ( .A1(n493), .A2(n481), .ZN(n482) );
  XOR2_X1 U540 ( .A(KEYINPUT101), .B(n482), .Z(n510) );
  NAND2_X1 U541 ( .A1(n497), .A2(n510), .ZN(n490) );
  NOR2_X1 U542 ( .A1(n576), .A2(n490), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U545 ( .A(G1GAT), .B(n485), .Z(G1324GAT) );
  INV_X1 U546 ( .A(n527), .ZN(n502) );
  NOR2_X1 U547 ( .A1(n502), .A2(n490), .ZN(n486) );
  XOR2_X1 U548 ( .A(G8GAT), .B(n486), .Z(G1325GAT) );
  NOR2_X1 U549 ( .A1(n541), .A2(n490), .ZN(n488) );
  XNOR2_X1 U550 ( .A(KEYINPUT35), .B(KEYINPUT103), .ZN(n487) );
  XNOR2_X1 U551 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U552 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  INV_X1 U553 ( .A(n532), .ZN(n539) );
  NOR2_X1 U554 ( .A1(n539), .A2(n490), .ZN(n491) );
  XOR2_X1 U555 ( .A(G22GAT), .B(n491), .Z(G1327GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT37), .B(KEYINPUT104), .Z(n496) );
  NAND2_X1 U557 ( .A1(n494), .A2(n561), .ZN(n495) );
  XOR2_X1 U558 ( .A(n496), .B(n495), .Z(n522) );
  XNOR2_X1 U559 ( .A(n498), .B(KEYINPUT105), .ZN(n499) );
  NOR2_X1 U560 ( .A1(n508), .A2(n576), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NOR2_X1 U563 ( .A1(n508), .A2(n502), .ZN(n503) );
  XOR2_X1 U564 ( .A(KEYINPUT106), .B(n503), .Z(n504) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(n504), .ZN(G1329GAT) );
  XNOR2_X1 U566 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n506) );
  NOR2_X1 U567 ( .A1(n541), .A2(n508), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NOR2_X1 U570 ( .A1(n539), .A2(n508), .ZN(n509) );
  XNOR2_X1 U571 ( .A(KEYINPUT108), .B(n294), .ZN(G1331GAT) );
  NOR2_X1 U572 ( .A1(n580), .A2(n556), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n510), .A2(n523), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(KEYINPUT109), .ZN(n517) );
  NAND2_X1 U575 ( .A1(n517), .A2(n525), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(KEYINPUT42), .ZN(n513) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n513), .ZN(G1332GAT) );
  NAND2_X1 U578 ( .A1(n517), .A2(n527), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(KEYINPUT110), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n529), .A2(n517), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U584 ( .A1(n517), .A2(n532), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n521) );
  XOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT112), .Z(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(KEYINPUT113), .B(n524), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n533), .A2(n525), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n526), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n533), .A2(n527), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n529), .A2(n533), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(KEYINPUT114), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT115), .B(KEYINPUT44), .Z(n535) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  NOR2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n552) );
  NAND2_X1 U602 ( .A1(n539), .A2(n552), .ZN(n540) );
  NOR2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n580), .A2(n548), .ZN(n542) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n544) );
  INV_X1 U607 ( .A(n556), .ZN(n569) );
  NAND2_X1 U608 ( .A1(n548), .A2(n569), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U610 ( .A(G120GAT), .B(n545), .Z(G1341GAT) );
  NAND2_X1 U611 ( .A1(n589), .A2(n548), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT50), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U615 ( .A1(n548), .A2(n458), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  INV_X1 U617 ( .A(n579), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n565) );
  NOR2_X1 U619 ( .A1(n553), .A2(n565), .ZN(n554) );
  XOR2_X1 U620 ( .A(G141GAT), .B(n554), .Z(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT120), .B(n555), .ZN(G1344GAT) );
  NOR2_X1 U622 ( .A1(n565), .A2(n556), .ZN(n560) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n565), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT122), .B(n562), .Z(n563) );
  XNOR2_X1 U629 ( .A(G155GAT), .B(n563), .ZN(G1346GAT) );
  INV_X1 U630 ( .A(n564), .ZN(n566) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  NAND2_X1 U633 ( .A1(n580), .A2(n574), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G169GAT), .B(n568), .ZN(G1348GAT) );
  XOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT56), .Z(n571) );
  NAND2_X1 U636 ( .A1(n574), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  NAND2_X1 U640 ( .A1(n574), .A2(n589), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT127), .Z(n582) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n588) );
  NAND2_X1 U645 ( .A1(n588), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n584) );
  XOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n587) );
  INV_X1 U650 ( .A(n588), .ZN(n591) );
  OR2_X1 U651 ( .A1(n591), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n492), .A2(n591), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

