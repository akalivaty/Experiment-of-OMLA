//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n188), .A2(G952), .ZN(new_n189));
  NAND2_X1  g003(.A1(G234), .A2(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT21), .B(G898), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n192), .B(KEYINPUT94), .Z(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(G902), .A3(G953), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G110), .B(G122), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n196), .B(KEYINPUT78), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n198));
  INV_X1    g012(.A(G113), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(KEYINPUT71), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT71), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(KEYINPUT2), .B2(G113), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n200), .A2(new_n202), .B1(KEYINPUT2), .B2(G113), .ZN(new_n203));
  XNOR2_X1  g017(.A(G116), .B(G119), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(new_n202), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT2), .A2(G113), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(new_n204), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT72), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n203), .A2(KEYINPUT72), .A3(new_n204), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n205), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G104), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G101), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n214), .A2(new_n217), .A3(new_n221), .A4(new_n218), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(new_n224), .A3(G101), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(KEYINPUT76), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT76), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n220), .A2(new_n227), .A3(KEYINPUT4), .A4(new_n222), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n212), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n210), .A2(new_n211), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n216), .A2(G104), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n213), .A2(G107), .ZN(new_n232));
  OAI21_X1  g046(.A(G101), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n222), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G116), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n237), .A2(KEYINPUT5), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G119), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n240), .A3(KEYINPUT5), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(G113), .A3(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n230), .A2(new_n235), .A3(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n197), .B1(new_n229), .B2(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n225), .A2(KEYINPUT76), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n228), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n212), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n230), .A2(new_n235), .A3(new_n242), .ZN(new_n250));
  INV_X1    g064(.A(new_n197), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n244), .A2(new_n252), .A3(new_n253), .A4(KEYINPUT6), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n244), .A2(new_n252), .A3(KEYINPUT6), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(new_n197), .C1(new_n229), .C2(new_n243), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT79), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n254), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n262), .A2(KEYINPUT65), .A3(G146), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT65), .B1(new_n262), .B2(G146), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT64), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT0), .A3(G128), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT0), .ZN(new_n270));
  INV_X1    g084(.A(G128), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n267), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n262), .A2(G146), .ZN(new_n274));
  INV_X1    g088(.A(new_n266), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(G143), .B2(new_n260), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n262), .A2(KEYINPUT66), .A3(G146), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n274), .B(new_n275), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G125), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n262), .A2(G146), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n283));
  OAI21_X1  g097(.A(G128), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n265), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G125), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT66), .B1(new_n262), .B2(G146), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n276), .A2(new_n260), .A3(G143), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n289), .A2(new_n283), .A3(G128), .A4(new_n274), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n285), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n281), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G224), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(G953), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n292), .B(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n259), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G210), .B1(G237), .B2(G902), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n291), .A2(KEYINPUT80), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT80), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n285), .A2(new_n290), .A3(new_n300), .A4(new_n286), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n281), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT7), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n303), .B2(new_n294), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n294), .A2(KEYINPUT81), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n303), .B1(new_n294), .B2(KEYINPUT81), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n292), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(new_n197), .B(KEYINPUT8), .Z(new_n308));
  AOI21_X1  g122(.A(new_n235), .B1(new_n230), .B2(new_n242), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n243), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n304), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT82), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n304), .A2(new_n307), .A3(new_n310), .A4(KEYINPUT82), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n252), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n297), .A2(new_n298), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n298), .B1(new_n297), .B2(new_n315), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n187), .B(new_n195), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G469), .ZN(new_n319));
  INV_X1    g133(.A(G902), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G140), .ZN(new_n322));
  INV_X1    g136(.A(G227), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G953), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n322), .B(new_n324), .Z(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n271), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n287), .A2(new_n288), .B1(new_n262), .B2(G146), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n290), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT10), .B1(new_n329), .B2(new_n235), .ZN(new_n330));
  INV_X1    g144(.A(new_n280), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n247), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n285), .A2(new_n290), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(KEYINPUT10), .A3(new_n235), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n333), .A2(KEYINPUT77), .A3(KEYINPUT10), .A4(new_n235), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G131), .ZN(new_n339));
  INV_X1    g153(.A(G137), .ZN(new_n340));
  INV_X1    g154(.A(G134), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT68), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G134), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n340), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT11), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n344), .A3(new_n340), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(KEYINPUT11), .A2(G134), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT69), .B1(new_n349), .B2(G137), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT69), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n351), .A2(new_n340), .A3(KEYINPUT11), .A4(G134), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n339), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT68), .B(G134), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT11), .B1(new_n356), .B2(new_n340), .ZN(new_n357));
  XOR2_X1   g171(.A(KEYINPUT70), .B(G131), .Z(new_n358));
  NOR4_X1   g172(.A1(new_n357), .A2(new_n353), .A3(new_n345), .A4(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n332), .A2(new_n338), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n332), .B2(new_n338), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n326), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n332), .A2(new_n338), .A3(new_n360), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n347), .A2(new_n346), .ZN(new_n365));
  INV_X1    g179(.A(new_n358), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n342), .A2(new_n344), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G137), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n354), .A2(new_n365), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n357), .A2(new_n345), .A3(new_n353), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(new_n339), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT12), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n328), .A2(new_n327), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n234), .B1(new_n373), .B2(new_n290), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n285), .A2(new_n290), .A3(new_n234), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n371), .B(new_n372), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT12), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n364), .A2(new_n376), .A3(new_n325), .A4(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(G902), .B1(new_n363), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n321), .B1(new_n380), .B2(new_n319), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n361), .A2(new_n362), .A3(new_n326), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n378), .A2(new_n376), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n325), .B1(new_n383), .B2(new_n364), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n381), .B1(new_n319), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G221), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT9), .B(G234), .Z(new_n389));
  AOI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(new_n320), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G116), .B(G122), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n216), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n262), .A2(G128), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n271), .A2(G143), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n397), .A2(new_n356), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n356), .ZN(new_n399));
  XOR2_X1   g213(.A(G116), .B(G122), .Z(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT14), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n239), .A2(KEYINPUT14), .A3(G122), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G107), .ZN(new_n403));
  OAI221_X1 g217(.A(new_n394), .B1(new_n398), .B2(new_n399), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(G107), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n399), .B1(new_n394), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT91), .ZN(new_n407));
  INV_X1    g221(.A(new_n395), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n408), .A2(KEYINPUT13), .B1(KEYINPUT90), .B2(new_n396), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT13), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n395), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n262), .A2(KEYINPUT90), .A3(KEYINPUT13), .A4(G128), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G134), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n406), .A2(new_n407), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n407), .B1(new_n406), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n404), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n389), .A2(G217), .A3(new_n188), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n418), .B(KEYINPUT92), .Z(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n405), .A2(new_n394), .ZN(new_n422));
  INV_X1    g236(.A(new_n399), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n413), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n396), .A2(KEYINPUT90), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n426), .B1(new_n410), .B2(new_n395), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n341), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT91), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n406), .A2(new_n407), .A3(new_n414), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n404), .A3(new_n419), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n421), .A2(new_n320), .A3(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT93), .ZN(new_n434));
  INV_X1    g248(.A(G478), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(KEYINPUT15), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n433), .B2(KEYINPUT93), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G475), .ZN(new_n441));
  NAND2_X1  g255(.A1(G125), .A2(G140), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(G125), .A2(G140), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G140), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n286), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT84), .B1(new_n448), .B2(new_n442), .ZN(new_n449));
  OAI21_X1  g263(.A(G146), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT85), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n442), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n260), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT85), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n454), .B(G146), .C1(new_n446), .C2(new_n449), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(KEYINPUT18), .A2(G131), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G237), .A2(G953), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(G143), .A3(G214), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(G143), .B1(new_n459), .B2(G214), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n458), .B1(new_n463), .B2(KEYINPUT83), .ZN(new_n464));
  INV_X1    g278(.A(G237), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n188), .A3(G214), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n262), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n460), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT83), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n457), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n463), .A2(KEYINPUT83), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n456), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n286), .A2(KEYINPUT16), .A3(G140), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n452), .B2(KEYINPUT16), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(new_n260), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n463), .A2(new_n366), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT17), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n468), .A2(new_n358), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n468), .A2(KEYINPUT17), .A3(new_n358), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n476), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n473), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(G113), .B(G122), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n213), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT89), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(G902), .B1(new_n483), .B2(new_n488), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n441), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n487), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n483), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n477), .A2(new_n479), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n475), .A2(G146), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT19), .B1(new_n446), .B2(new_n449), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT19), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n452), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT86), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT86), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n452), .A2(new_n501), .A3(new_n498), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n495), .B(new_n496), .C1(new_n503), .C2(G146), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n473), .A2(new_n487), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n493), .A2(new_n494), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n493), .A2(new_n505), .A3(new_n441), .A4(new_n320), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n473), .A2(new_n487), .A3(new_n504), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n487), .B1(new_n473), .B2(new_n482), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n511), .A2(new_n512), .A3(G475), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n513), .A2(new_n506), .A3(new_n507), .A4(new_n320), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n491), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR4_X1   g330(.A1(new_n318), .A2(new_n392), .A3(new_n440), .A4(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G472), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n347), .B1(G134), .B2(new_n340), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n285), .A2(new_n290), .B1(new_n519), .B2(G131), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n369), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n280), .A2(KEYINPUT67), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT67), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT65), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n274), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n262), .A2(KEYINPUT65), .A3(G146), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n282), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n267), .A2(new_n269), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n270), .A2(new_n271), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n279), .B(new_n523), .C1(new_n527), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n522), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n521), .B1(new_n532), .B2(new_n360), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n248), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT28), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n371), .A2(new_n331), .B1(new_n369), .B2(new_n520), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(new_n212), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n331), .B1(new_n355), .B2(new_n359), .ZN(new_n538));
  AND4_X1   g352(.A1(new_n535), .A2(new_n538), .A3(new_n212), .A4(new_n521), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n534), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  XOR2_X1   g354(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n541));
  NAND2_X1  g355(.A1(new_n459), .A2(G210), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT26), .B(G101), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n538), .A2(KEYINPUT30), .A3(new_n521), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n519), .A2(G131), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n333), .A2(new_n369), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n531), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n523), .B1(new_n273), .B2(new_n279), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n549), .B1(new_n552), .B2(new_n371), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n248), .B(new_n547), .C1(new_n553), .C2(KEYINPUT30), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n536), .A2(new_n212), .ZN(new_n555));
  INV_X1    g369(.A(new_n545), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n546), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT29), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n537), .A2(new_n539), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n536), .A2(new_n212), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n556), .A2(new_n559), .ZN(new_n565));
  AOI21_X1  g379(.A(G902), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n518), .B1(new_n560), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n554), .A2(new_n555), .A3(new_n545), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n568), .A2(KEYINPUT74), .A3(KEYINPUT31), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT74), .B1(new_n568), .B2(KEYINPUT31), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n540), .A2(new_n556), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT31), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n554), .A2(new_n572), .A3(new_n555), .A4(new_n545), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n569), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT32), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n571), .A2(new_n573), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n568), .A2(KEYINPUT31), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT74), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n568), .A2(KEYINPUT74), .A3(KEYINPUT31), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT32), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(new_n576), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n567), .B1(new_n578), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT75), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT25), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT23), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n236), .B2(G128), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n271), .A2(KEYINPUT23), .A3(G119), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n592), .B(new_n593), .C1(G119), .C2(new_n271), .ZN(new_n594));
  XNOR2_X1  g408(.A(G119), .B(G128), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT24), .B(G110), .Z(new_n596));
  OAI22_X1  g410(.A1(new_n594), .A2(G110), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n496), .A3(new_n453), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(G110), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n595), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n598), .B1(new_n476), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT22), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(new_n340), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n602), .A2(new_n605), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n590), .B1(new_n609), .B2(G902), .ZN(new_n610));
  INV_X1    g424(.A(G217), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(G234), .B2(new_n320), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n608), .A2(new_n588), .A3(new_n589), .A4(new_n320), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n612), .A2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n587), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n517), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT95), .B(G101), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G3));
  AOI21_X1  g435(.A(new_n518), .B1(new_n584), .B2(new_n320), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n576), .B2(new_n584), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n617), .A2(new_n390), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n623), .A2(new_n387), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT96), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT97), .B(G478), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n433), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n417), .A2(new_n420), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n419), .B1(new_n431), .B2(new_n404), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n421), .A2(KEYINPUT33), .A3(new_n432), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n629), .B1(new_n635), .B2(G478), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n516), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n318), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n626), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  XNOR2_X1  g456(.A(new_n491), .B(KEYINPUT98), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n509), .B(KEYINPUT20), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n440), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n318), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n626), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n605), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n602), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n615), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n614), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n517), .A2(new_n623), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT37), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G110), .ZN(G12));
  OAI211_X1 g472(.A(new_n655), .B(new_n187), .C1(new_n316), .C2(new_n317), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n587), .A2(new_n392), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n191), .B(KEYINPUT99), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(G900), .B2(new_n194), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n646), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n663), .B(KEYINPUT39), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n387), .A2(new_n391), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n259), .A2(new_n296), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n320), .A3(new_n315), .ZN(new_n674));
  INV_X1    g488(.A(new_n298), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n297), .A2(new_n298), .A3(new_n315), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT38), .ZN(new_n679));
  INV_X1    g493(.A(new_n187), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n655), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n672), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n584), .A2(new_n585), .A3(new_n576), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n585), .B1(new_n584), .B2(new_n576), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n555), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n556), .B1(new_n563), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(G472), .A3(new_n568), .ZN(new_n688));
  NAND2_X1  g502(.A1(G472), .A2(G902), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n690), .B(KEYINPUT100), .Z(new_n691));
  NOR2_X1   g505(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n439), .A2(new_n515), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n668), .B1(new_n682), .B2(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n692), .A2(new_n439), .A3(new_n515), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n679), .A2(new_n681), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n697), .A2(new_n698), .A3(KEYINPUT101), .A4(new_n672), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n262), .ZN(G45));
  INV_X1    g515(.A(new_n567), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n702), .B1(new_n683), .B2(new_n684), .ZN(new_n703));
  AOI211_X1 g517(.A(new_n680), .B(new_n654), .C1(new_n676), .C2(new_n677), .ZN(new_n704));
  INV_X1    g518(.A(new_n392), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n515), .A2(new_n636), .A3(new_n664), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n578), .A2(new_n586), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n392), .B1(new_n709), .B2(new_n702), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n704), .A4(new_n706), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  INV_X1    g528(.A(new_n617), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n380), .A2(new_n319), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n380), .A2(new_n319), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n391), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n639), .A2(new_n703), .A3(new_n715), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  NAND3_X1  g536(.A1(new_n618), .A2(new_n647), .A3(new_n719), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G116), .ZN(G18));
  NAND2_X1  g538(.A1(new_n655), .A2(new_n195), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n709), .B2(new_n702), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n440), .A2(new_n516), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n187), .B1(new_n316), .B2(new_n317), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n728), .A2(new_n729), .A3(new_n718), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n680), .B1(new_n676), .B2(new_n677), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT103), .B1(new_n731), .B2(new_n719), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n726), .B(new_n727), .C1(new_n730), .C2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  AND3_X1   g548(.A1(new_n731), .A2(new_n694), .A3(new_n719), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n580), .B(new_n573), .C1(new_n545), .C2(new_n564), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n576), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(KEYINPUT104), .A3(new_n576), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n622), .A3(new_n617), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n735), .A2(new_n742), .A3(new_n195), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  INV_X1    g558(.A(new_n706), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n729), .B1(new_n728), .B2(new_n718), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n731), .A2(KEYINPUT103), .A3(new_n719), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n741), .A2(new_n622), .A3(new_n654), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  OAI21_X1  g565(.A(KEYINPUT105), .B1(new_n382), .B2(new_n384), .ZN(new_n752));
  INV_X1    g566(.A(new_n362), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n364), .A3(new_n325), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(G469), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n381), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n706), .A2(new_n758), .A3(new_n391), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n676), .A2(new_n187), .A3(new_n677), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n703), .A3(new_n715), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n761), .A2(new_n703), .A3(KEYINPUT106), .A4(new_n715), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n709), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n578), .A2(KEYINPUT107), .A3(new_n586), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n702), .A3(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(KEYINPUT42), .A3(new_n715), .A4(new_n761), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  NOR3_X1   g588(.A1(new_n587), .A2(new_n617), .A3(new_n760), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n390), .B1(new_n757), .B2(new_n381), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n775), .A2(new_n665), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n341), .ZN(G36));
  NAND2_X1  g592(.A1(new_n637), .A2(new_n515), .ZN(new_n779));
  AND2_X1   g593(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n780));
  NOR2_X1   g594(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n780), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n623), .B1(new_n785), .B2(KEYINPUT110), .ZN(new_n786));
  INV_X1    g600(.A(new_n784), .ZN(new_n787));
  OR3_X1    g601(.A1(new_n787), .A2(new_n782), .A3(KEYINPUT110), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n655), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n760), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n752), .A2(KEYINPUT45), .A3(new_n756), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n792), .B(G469), .C1(KEYINPUT45), .C2(new_n385), .ZN(new_n793));
  INV_X1    g607(.A(new_n321), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT46), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(KEYINPUT46), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n717), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n391), .A3(new_n669), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT108), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n786), .A2(KEYINPUT44), .A3(new_n655), .A4(new_n788), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT108), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n798), .A2(new_n802), .A3(new_n391), .A4(new_n669), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n791), .A2(new_n800), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT111), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n340), .ZN(G39));
  NOR3_X1   g620(.A1(new_n703), .A2(new_n715), .A3(new_n760), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n798), .A2(KEYINPUT47), .A3(new_n391), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT47), .B1(new_n798), .B2(new_n391), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n706), .B(new_n807), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  NOR2_X1   g626(.A1(new_n693), .A2(new_n191), .ZN(new_n813));
  INV_X1    g627(.A(new_n760), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n715), .A3(new_n719), .A4(new_n814), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n815), .A2(new_n516), .A3(new_n637), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n785), .A2(new_n662), .A3(new_n718), .A4(new_n760), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT115), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n749), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n661), .A2(new_n742), .A3(new_n784), .A4(new_n783), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n719), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n187), .A3(new_n679), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT50), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n821), .A2(new_n814), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n809), .A2(new_n810), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n716), .A2(new_n390), .A3(new_n717), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT51), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n827), .A2(KEYINPUT113), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n809), .B2(new_n810), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n833), .A3(new_n828), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n835));
  INV_X1    g649(.A(new_n826), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n824), .A4(new_n820), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n835), .B1(new_n834), .B2(new_n836), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n830), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n821), .B1(new_n732), .B2(new_n730), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n703), .A2(new_n705), .A3(new_n439), .A4(new_n663), .ZN(new_n843));
  INV_X1    g657(.A(new_n645), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n741), .A2(new_n759), .A3(new_n622), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n655), .B(new_n814), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n777), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n773), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n733), .A2(new_n723), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n656), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n515), .A2(new_n636), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n440), .B2(new_n515), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n318), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n625), .A2(new_n855), .B1(new_n517), .B2(new_n618), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n743), .A2(new_n720), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n851), .A2(new_n852), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n849), .A2(new_n859), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n748), .A2(new_n749), .B1(new_n660), .B2(new_n665), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n731), .A2(new_n694), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n654), .A2(new_n663), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT112), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n693), .A2(new_n863), .A3(new_n776), .A4(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n861), .A2(new_n713), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT52), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n861), .A2(new_n713), .A3(new_n866), .A4(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n870), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n850), .A2(new_n656), .A3(new_n857), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n777), .B1(new_n767), .B2(new_n772), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n856), .A4(new_n847), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n872), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n871), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n871), .A2(new_n877), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT54), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n841), .A2(new_n842), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n771), .A2(new_n715), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n818), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT48), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n885), .B(new_n189), .C1(new_n638), .C2(new_n815), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n882), .A2(new_n886), .B1(G952), .B2(G953), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n716), .A2(new_n717), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n779), .B(new_n693), .C1(KEYINPUT49), .C2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n624), .B1(new_n888), .B2(KEYINPUT49), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n679), .A2(new_n680), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n892), .ZN(G75));
  NOR2_X1   g707(.A1(new_n188), .A2(G952), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n871), .A2(new_n877), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n320), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT56), .B1(new_n897), .B2(G210), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n259), .B(new_n295), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT55), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n895), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  XOR2_X1   g715(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n897), .B2(G210), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(G51));
  NAND2_X1  g719(.A1(new_n363), .A2(new_n379), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT117), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n880), .B2(KEYINPUT54), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n881), .A2(new_n879), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n907), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n321), .B(KEYINPUT57), .Z(new_n911));
  OAI21_X1  g725(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n896), .A2(new_n320), .A3(new_n793), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n894), .B1(new_n912), .B2(new_n913), .ZN(G54));
  NAND3_X1  g728(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n493), .A2(new_n505), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n917), .A2(new_n918), .A3(new_n894), .ZN(G60));
  NAND2_X1  g733(.A1(new_n633), .A2(new_n634), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT59), .Z(new_n923));
  NOR3_X1   g737(.A1(new_n910), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n881), .B2(new_n879), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n920), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n895), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n926), .A2(new_n925), .A3(new_n920), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n924), .A2(new_n928), .A3(new_n929), .ZN(G63));
  XNOR2_X1  g744(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT119), .B1(new_n880), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n936));
  AOI211_X1 g750(.A(new_n936), .B(new_n933), .C1(new_n871), .C2(new_n877), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n894), .B1(new_n938), .B2(new_n609), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n652), .B1(new_n935), .B2(new_n937), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n931), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n936), .B1(new_n896), .B2(new_n933), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n880), .A2(KEYINPUT119), .A3(new_n934), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n609), .A3(new_n943), .ZN(new_n944));
  AND4_X1   g758(.A1(new_n895), .A2(new_n944), .A3(new_n940), .A4(new_n931), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n941), .A2(new_n945), .ZN(G66));
  INV_X1    g760(.A(new_n193), .ZN(new_n947));
  OAI21_X1  g761(.A(G953), .B1(new_n947), .B2(new_n293), .ZN(new_n948));
  INV_X1    g762(.A(new_n859), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(G953), .ZN(new_n950));
  INV_X1    g764(.A(new_n259), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(G898), .B2(new_n188), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n950), .B(new_n952), .ZN(G69));
  OAI21_X1  g767(.A(new_n547), .B1(new_n553), .B2(KEYINPUT30), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n503), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n861), .A2(new_n713), .ZN(new_n956));
  NOR2_X1   g770(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n957));
  OR3_X1    g771(.A1(new_n700), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n700), .B2(new_n956), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n804), .A2(new_n811), .A3(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n854), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n775), .A2(new_n705), .A3(new_n669), .A4(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n960), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT122), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT122), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n960), .A2(new_n962), .A3(new_n967), .A4(new_n964), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n955), .B1(new_n969), .B2(new_n188), .ZN(new_n970));
  INV_X1    g784(.A(new_n955), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n804), .A2(new_n811), .ZN(new_n972));
  INV_X1    g786(.A(new_n875), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n973), .A2(KEYINPUT124), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n972), .A2(new_n974), .A3(new_n956), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n800), .A2(new_n863), .A3(new_n883), .A4(new_n803), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n973), .A2(KEYINPUT124), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n188), .ZN(new_n979));
  INV_X1    g793(.A(G900), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(G953), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n971), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n970), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(G953), .B1(new_n323), .B2(new_n980), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT123), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n970), .B2(new_n982), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(G72));
  NAND2_X1  g803(.A1(new_n554), .A2(new_n555), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n545), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n689), .B(KEYINPUT63), .Z(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n557), .A3(new_n992), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT126), .Z(new_n994));
  NOR2_X1   g808(.A1(new_n896), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT127), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n966), .A2(new_n949), .A3(new_n968), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n992), .B(KEYINPUT125), .Z(new_n998));
  AOI21_X1  g812(.A(new_n991), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n975), .A2(new_n949), .A3(new_n976), .A4(new_n977), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n557), .B1(new_n1000), .B2(new_n998), .ZN(new_n1001));
  NOR4_X1   g815(.A1(new_n996), .A2(new_n999), .A3(new_n894), .A4(new_n1001), .ZN(G57));
endmodule


