//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G141gat), .B(G148gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n202), .B(new_n205), .C1(new_n206), .C2(KEYINPUT2), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(new_n202), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n207), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(KEYINPUT73), .A2(G204gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT73), .A2(G204gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(G197gat), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G197gat), .ZN(new_n220));
  AND2_X1   g019(.A1(KEYINPUT73), .A2(G204gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT73), .A2(G204gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G211gat), .A2(G218gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT22), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n219), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G211gat), .ZN(new_n228));
  INV_X1    g027(.A(G218gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(new_n224), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n219), .A2(new_n223), .A3(new_n232), .A4(new_n226), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT29), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n237), .B1(new_n236), .B2(new_n238), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n216), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n207), .A2(new_n240), .A3(new_n215), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT76), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n207), .A2(new_n215), .A3(KEYINPUT76), .A4(new_n240), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n238), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT83), .ZN(new_n250));
  INV_X1    g049(.A(new_n236), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G228gat), .ZN(new_n253));
  INV_X1    g052(.A(G233gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT29), .B1(new_n246), .B2(new_n247), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT83), .B1(new_n256), .B2(new_n236), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n243), .A2(new_n252), .A3(new_n255), .A4(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n216), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n230), .A2(new_n224), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n227), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n260), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n262), .A2(new_n219), .A3(new_n223), .A4(new_n226), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n238), .A3(new_n263), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n264), .A2(KEYINPUT81), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT3), .B1(new_n264), .B2(KEYINPUT81), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n259), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n256), .A2(new_n236), .ZN(new_n268));
  OAI22_X1  g067(.A1(new_n267), .A2(new_n268), .B1(new_n253), .B2(new_n254), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n258), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT84), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT84), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n258), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(G22gat), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT85), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n271), .A2(KEYINPUT85), .A3(G22gat), .A4(new_n273), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(G50gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(G78gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(G106gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT86), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n270), .B2(G22gat), .ZN(new_n283));
  INV_X1    g082(.A(G22gat), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n258), .A2(new_n269), .A3(KEYINPUT86), .A4(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n281), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n276), .A2(new_n277), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n270), .A2(G22gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n284), .B1(new_n258), .B2(new_n269), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n281), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n287), .A2(KEYINPUT87), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT87), .B1(new_n287), .B2(new_n290), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT70), .B(G127gat), .ZN(new_n293));
  INV_X1    g092(.A(G134gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G113gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT69), .B(G113gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(new_n297), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n295), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT67), .B(G134gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G127gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT68), .B(G127gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G134gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G113gat), .B(G120gat), .Z(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n296), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n301), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT4), .B1(new_n310), .B2(new_n216), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n300), .A2(new_n296), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n312), .A2(new_n295), .B1(new_n306), .B2(new_n308), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT4), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n314), .A3(new_n259), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(KEYINPUT79), .A3(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n248), .B(new_n310), .C1(new_n240), .C2(new_n259), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT79), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n318), .B(KEYINPUT4), .C1(new_n310), .C2(new_n216), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OR3_X1    g121(.A1(new_n320), .A2(KEYINPUT5), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n313), .B(new_n216), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n324), .B1(new_n325), .B2(new_n321), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n315), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(new_n321), .A3(new_n317), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n313), .B(new_n259), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT77), .A3(new_n322), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n326), .A2(new_n328), .A3(new_n330), .A4(KEYINPUT5), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(G1gat), .B(G29gat), .Z(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G57gat), .B(G85gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT6), .ZN(new_n339));
  INV_X1    g138(.A(new_n337), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n331), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n332), .A2(KEYINPUT6), .A3(new_n337), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n345));
  INV_X1    g144(.A(G169gat), .ZN(new_n346));
  INV_X1    g145(.A(G176gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n348), .A2(new_n349), .B1(G169gat), .B2(G176gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n351), .B(KEYINPUT64), .Z(new_n352));
  NAND2_X1  g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT24), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n344), .B(new_n350), .C1(new_n352), .C2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n350), .B1(new_n355), .B2(new_n351), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT25), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT26), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n346), .A2(new_n347), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G183gat), .ZN(new_n364));
  OAI211_X1 g163(.A(KEYINPUT65), .B(KEYINPUT27), .C1(new_n364), .C2(KEYINPUT66), .ZN(new_n365));
  NAND2_X1  g164(.A1(KEYINPUT65), .A2(KEYINPUT27), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT66), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(G183gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT65), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n369), .B1(new_n370), .B2(G183gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n365), .A2(new_n368), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n363), .B(new_n353), .C1(G190gat), .C2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT27), .B(G183gat), .ZN(new_n375));
  INV_X1    g174(.A(G190gat), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n359), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(KEYINPUT29), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(G226gat), .B2(G233gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT75), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n236), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n383), .ZN(new_n386));
  OAI221_X1 g185(.A(new_n251), .B1(new_n382), .B2(new_n379), .C1(new_n380), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390));
  INV_X1    g189(.A(G64gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G92gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n388), .A2(new_n389), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n388), .A2(new_n395), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n385), .A2(new_n387), .A3(new_n394), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(KEYINPUT30), .A3(new_n398), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n342), .A2(new_n343), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n291), .A2(new_n292), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G15gat), .B(G43gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(G71gat), .B(G99gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  INV_X1    g203(.A(G227gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n405), .A2(new_n254), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n310), .B1(new_n359), .B2(new_n378), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n373), .A2(G190gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n377), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n409), .A2(new_n353), .A3(new_n410), .A4(new_n363), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n313), .A2(new_n411), .A3(new_n358), .A4(new_n356), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n407), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n404), .B1(new_n413), .B2(KEYINPUT33), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT32), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n408), .A2(new_n412), .A3(new_n407), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT34), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n408), .A2(new_n412), .ZN(new_n421));
  AOI221_X4 g220(.A(new_n415), .B1(KEYINPUT33), .B2(new_n404), .C1(new_n421), .C2(new_n406), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n417), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n414), .A2(new_n416), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n419), .B1(new_n425), .B2(new_n422), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT71), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT36), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n417), .A2(new_n420), .A3(KEYINPUT71), .A4(new_n423), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT72), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n424), .A2(new_n426), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT36), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n428), .A2(KEYINPUT72), .A3(new_n429), .A4(new_n430), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT88), .B1(new_n401), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n342), .A2(new_n343), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT37), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n395), .B1(new_n388), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT38), .ZN(new_n445));
  OAI22_X1  g244(.A1(new_n380), .A2(new_n386), .B1(new_n382), .B2(new_n379), .ZN(new_n446));
  OR3_X1    g245(.A1(new_n446), .A2(KEYINPUT92), .A3(new_n251), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n251), .B1(new_n381), .B2(new_n384), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT92), .B1(new_n446), .B2(new_n251), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n444), .B(new_n445), .C1(new_n450), .C2(new_n443), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n444), .B1(new_n443), .B2(new_n388), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT38), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n442), .A2(new_n397), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n287), .A2(new_n290), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n287), .A2(KEYINPUT87), .A3(new_n290), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n320), .A2(new_n322), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n325), .A2(new_n321), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT39), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT89), .B(KEYINPUT39), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n320), .A2(new_n322), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n340), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT40), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n462), .A2(KEYINPUT90), .A3(new_n340), .A4(new_n464), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT91), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n399), .A2(new_n396), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n465), .A2(new_n468), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n471), .A2(new_n338), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n470), .A2(KEYINPUT91), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n454), .B(new_n459), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n441), .A2(new_n472), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n457), .A2(new_n478), .A3(new_n458), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(new_n438), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n440), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n400), .B(new_n435), .C1(new_n291), .C2(new_n292), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT35), .ZN(new_n484));
  NAND2_X1  g283(.A1(KEYINPUT93), .A2(KEYINPUT35), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n428), .A2(new_n430), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n459), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n400), .B1(KEYINPUT93), .B2(KEYINPUT35), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT16), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(G1gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(G1gat), .B2(new_n491), .ZN(new_n494));
  INV_X1    g293(.A(G8gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(G71gat), .A2(G78gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT9), .ZN(new_n498));
  NAND2_X1  g297(.A1(G71gat), .A2(G78gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n391), .A2(G57gat), .ZN(new_n500));
  INV_X1    g299(.A(G57gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(G64gat), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n498), .A2(new_n499), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n502), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT97), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT97), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n500), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(KEYINPUT9), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n499), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(new_n497), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n503), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT21), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(new_n364), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT98), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT19), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n511), .A2(KEYINPUT21), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n517), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT99), .B(G211gat), .Z(new_n520));
  NAND2_X1  g319(.A1(G231gat), .A2(G233gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G127gat), .B(G155gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT20), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n522), .B(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n525), .B1(new_n518), .B2(new_n519), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT94), .B(G36gat), .Z(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G29gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT14), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(G29gat), .B2(G36gat), .ZN(new_n532));
  OR3_X1    g331(.A1(new_n531), .A2(G29gat), .A3(G36gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537));
  INV_X1    g336(.A(G43gat), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT95), .B1(new_n538), .B2(G50gat), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n539), .A2(new_n535), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n536), .B(new_n537), .C1(new_n540), .C2(new_n534), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n534), .A2(new_n540), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT17), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n496), .B(KEYINPUT96), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n496), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT18), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n543), .B(new_n547), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n549), .B(KEYINPUT13), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n546), .A2(KEYINPUT18), .A3(new_n548), .A4(new_n549), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT11), .B(G169gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G197gat), .ZN(new_n559));
  XOR2_X1   g358(.A(G113gat), .B(G141gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT12), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n552), .A2(new_n562), .A3(new_n555), .A4(new_n556), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n568), .B1(new_n569), .B2(new_n393), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n569), .B2(new_n393), .ZN(new_n572));
  NAND3_X1  g371(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n568), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n568), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n570), .A2(new_n577), .A3(new_n572), .A4(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n510), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n500), .A2(new_n502), .A3(new_n506), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n506), .B1(new_n500), .B2(new_n502), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n580), .B1(new_n583), .B2(KEYINPUT9), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n579), .B1(new_n584), .B2(new_n503), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT10), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n508), .A2(new_n510), .ZN(new_n587));
  INV_X1    g386(.A(new_n503), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n587), .A2(new_n578), .A3(new_n576), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT102), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n579), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(KEYINPUT10), .A3(new_n511), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n585), .A2(new_n589), .A3(KEYINPUT102), .A4(new_n586), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT103), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT103), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n592), .A2(new_n598), .A3(new_n594), .A4(new_n595), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n589), .ZN(new_n603));
  INV_X1    g402(.A(new_n601), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G120gat), .B(G148gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n347), .ZN(new_n607));
  INV_X1    g406(.A(G204gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n602), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n601), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n612), .A2(new_n605), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n613), .B2(new_n610), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n614), .A2(KEYINPUT104), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(KEYINPUT104), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n567), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n544), .A2(new_n579), .ZN(new_n619));
  AND2_X1   g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n543), .A2(new_n593), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n622), .A2(new_n623), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n627));
  XNOR2_X1  g426(.A(G190gat), .B(G218gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G134gat), .B(G162gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n625), .A2(new_n626), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n625), .B2(new_n626), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n528), .A2(new_n618), .A3(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n490), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n442), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT105), .B(G1gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(G1324gat));
  INV_X1    g439(.A(KEYINPUT42), .ZN(new_n641));
  INV_X1    g440(.A(new_n637), .ZN(new_n642));
  OAI21_X1  g441(.A(G8gat), .B1(new_n642), .B2(new_n472), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT106), .B(G8gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(new_n492), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n637), .A2(new_n473), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n641), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n641), .B2(new_n646), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT107), .ZN(G1325gat));
  AOI21_X1  g448(.A(G15gat), .B1(new_n637), .B2(new_n486), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n637), .A2(G15gat), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT108), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n438), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n433), .A2(KEYINPUT108), .A3(new_n436), .A4(new_n437), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n650), .B1(new_n651), .B2(new_n656), .ZN(G1326gat));
  INV_X1    g456(.A(new_n459), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n637), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT43), .B(G22gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  INV_X1    g460(.A(new_n528), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n618), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n490), .A2(new_n635), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(G29gat), .A3(new_n441), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT45), .Z(new_n667));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n490), .B2(new_n635), .ZN(new_n669));
  INV_X1    g468(.A(new_n635), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n457), .A2(new_n478), .A3(KEYINPUT109), .A4(new_n458), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n479), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n477), .A2(new_n655), .A3(new_n673), .A4(new_n675), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n670), .B(new_n672), .C1(new_n676), .C2(new_n489), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n678), .A2(new_n663), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n442), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(G29gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n667), .A2(new_n681), .ZN(G1328gat));
  NOR3_X1   g481(.A1(new_n665), .A2(new_n472), .A3(new_n529), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT46), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n679), .A2(new_n473), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n529), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(G1329gat));
  NAND3_X1  g486(.A1(new_n679), .A2(G43gat), .A3(new_n656), .ZN(new_n688));
  INV_X1    g487(.A(new_n486), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n538), .B1(new_n665), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g491(.A1(new_n678), .A2(new_n658), .A3(new_n663), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT111), .B1(new_n693), .B2(G50gat), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n665), .A2(G50gat), .A3(new_n459), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n697), .B1(new_n693), .B2(G50gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n696), .B(new_n698), .ZN(G1331gat));
  OAI211_X1 g498(.A(new_n566), .B(new_n670), .C1(new_n526), .C2(new_n527), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n676), .B2(new_n489), .ZN(new_n701));
  INV_X1    g500(.A(new_n617), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n441), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(new_n501), .ZN(G1332gat));
  NOR2_X1   g504(.A1(new_n703), .A2(new_n472), .ZN(new_n706));
  NOR2_X1   g505(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n707));
  AND2_X1   g506(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n706), .B2(new_n707), .ZN(G1333gat));
  INV_X1    g509(.A(new_n703), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(G71gat), .A3(new_n656), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n703), .A2(new_n689), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(G71gat), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n658), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g516(.A1(new_n676), .A2(new_n489), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n662), .A2(new_n567), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(new_n635), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(new_n442), .A3(new_n702), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n662), .A2(new_n567), .A3(new_n617), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n678), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n441), .A2(new_n569), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n723), .A2(new_n569), .B1(new_n725), .B2(new_n726), .ZN(G1336gat));
  NAND4_X1  g526(.A1(new_n722), .A2(new_n393), .A3(new_n473), .A4(new_n702), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n473), .B(new_n724), .C1(new_n669), .C2(new_n677), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G92gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(KEYINPUT112), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n730), .A2(new_n734), .A3(G92gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n728), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT52), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n736), .B2(KEYINPUT52), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n732), .B1(new_n738), .B2(new_n739), .ZN(G1337gat));
  INV_X1    g539(.A(G99gat), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n722), .A2(new_n741), .A3(new_n486), .A4(new_n702), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n725), .A2(new_n656), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(new_n741), .ZN(G1338gat));
  NAND2_X1  g543(.A1(new_n725), .A2(new_n658), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G106gat), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n459), .A2(G106gat), .A3(new_n617), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT53), .B1(new_n722), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT114), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n722), .A2(new_n751), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n747), .A2(new_n750), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n745), .A2(G106gat), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n749), .B1(new_n754), .B2(new_n755), .ZN(G1339gat));
  NOR2_X1   g555(.A1(new_n700), .A2(new_n702), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n604), .B1(new_n597), .B2(new_n599), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n596), .A2(new_n601), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n609), .B1(new_n612), .B2(KEYINPUT54), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n761), .A2(KEYINPUT55), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764));
  INV_X1    g563(.A(new_n760), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n602), .A2(KEYINPUT54), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n762), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n611), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n549), .B1(new_n546), .B2(new_n548), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n553), .A2(new_n554), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n561), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n565), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n633), .B2(new_n634), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT55), .B1(new_n761), .B2(new_n762), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n766), .A2(new_n764), .A3(new_n767), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(KEYINPUT115), .A3(new_n611), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n771), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT116), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n771), .A2(new_n776), .A3(new_n783), .A4(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT115), .B1(new_n779), .B2(new_n611), .ZN(new_n786));
  INV_X1    g585(.A(new_n611), .ZN(new_n787));
  AOI211_X1 g586(.A(new_n770), .B(new_n787), .C1(new_n777), .C2(new_n778), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n786), .A2(new_n788), .A3(new_n566), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n617), .A2(new_n775), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n670), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n757), .B1(new_n792), .B2(new_n528), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n793), .A2(new_n658), .A3(new_n689), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n473), .A2(new_n441), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT117), .ZN(new_n797));
  OAI21_X1  g596(.A(G113gat), .B1(new_n797), .B2(new_n566), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n793), .A2(new_n658), .A3(new_n434), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n566), .A2(new_n299), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1340gat));
  OAI21_X1  g601(.A(G120gat), .B1(new_n797), .B2(new_n617), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(new_n297), .A3(new_n795), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n617), .B2(new_n804), .ZN(G1341gat));
  NOR3_X1   g604(.A1(new_n797), .A2(new_n304), .A3(new_n528), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n799), .A2(new_n662), .A3(new_n795), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n304), .B2(new_n807), .ZN(G1342gat));
  OAI21_X1  g607(.A(G134gat), .B1(new_n797), .B2(new_n670), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n799), .A2(new_n302), .A3(new_n635), .A4(new_n795), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT56), .Z(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1343gat));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n793), .B2(new_n459), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT118), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n662), .B1(new_n785), .B2(new_n791), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n658), .B1(new_n816), .B2(new_n757), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n818), .A3(new_n813), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n617), .A2(new_n775), .B1(new_n566), .B2(new_n769), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n670), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n820), .A2(new_n822), .B1(new_n782), .B2(new_n784), .ZN(new_n823));
  INV_X1    g622(.A(new_n822), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT119), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n662), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT57), .B(new_n658), .C1(new_n826), .C2(new_n757), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n815), .A2(new_n819), .A3(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n655), .A2(new_n795), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n567), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G141gat), .ZN(new_n831));
  INV_X1    g630(.A(new_n817), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n829), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n208), .A3(new_n567), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT58), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n831), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(G1344gat));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n828), .A2(new_n829), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n841), .B(G148gat), .C1(new_n842), .C2(new_n617), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n817), .A2(KEYINPUT57), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n670), .A2(new_n775), .A3(new_n769), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n662), .B1(new_n822), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n813), .B(new_n658), .C1(new_n847), .C2(new_n757), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n844), .A2(new_n702), .A3(new_n829), .A4(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(new_n210), .ZN(new_n853));
  XNOR2_X1  g652(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n843), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n834), .A2(new_n210), .A3(new_n702), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1345gat));
  NOR3_X1   g656(.A1(new_n842), .A2(new_n203), .A3(new_n528), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n834), .A2(new_n662), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT122), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n858), .B1(new_n860), .B2(new_n203), .ZN(G1346gat));
  NOR3_X1   g660(.A1(new_n842), .A2(new_n204), .A3(new_n670), .ZN(new_n862));
  AOI21_X1  g661(.A(G162gat), .B1(new_n834), .B2(new_n635), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(G1347gat));
  NOR2_X1   g663(.A1(new_n442), .A2(new_n472), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n799), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n346), .A3(new_n567), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n794), .A2(new_n865), .ZN(new_n869));
  OAI21_X1  g668(.A(G169gat), .B1(new_n869), .B2(new_n566), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1348gat));
  NOR3_X1   g670(.A1(new_n869), .A2(new_n347), .A3(new_n617), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n867), .A2(new_n702), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n347), .B2(new_n873), .ZN(G1349gat));
  OAI21_X1  g673(.A(G183gat), .B1(new_n869), .B2(new_n528), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n662), .A2(new_n375), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n866), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g677(.A(G190gat), .B1(new_n869), .B2(new_n670), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT61), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n867), .A2(new_n376), .A3(new_n635), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1351gat));
  AND2_X1   g681(.A1(new_n655), .A2(new_n865), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n832), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(G197gat), .B1(new_n885), .B2(new_n567), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n844), .A2(new_n848), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n883), .B(KEYINPUT123), .Z(new_n888));
  AND2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n566), .A2(new_n220), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G1352gat));
  NOR3_X1   g690(.A1(new_n884), .A2(G204gat), .A3(new_n617), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT62), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n887), .A2(new_n702), .A3(new_n888), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n608), .B2(new_n894), .ZN(G1353gat));
  NAND4_X1  g694(.A1(new_n885), .A2(KEYINPUT124), .A3(new_n228), .A4(new_n662), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n832), .A2(new_n228), .A3(new_n883), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n528), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n844), .A2(new_n662), .A3(new_n848), .A4(new_n883), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n902), .A3(G211gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(G211gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT63), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n900), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n900), .A2(new_n905), .A3(KEYINPUT125), .A4(new_n903), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1354gat));
  NAND2_X1  g709(.A1(new_n635), .A2(G218gat), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT126), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n887), .A2(new_n888), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n229), .B1(new_n884), .B2(new_n670), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n915), .B(KEYINPUT127), .Z(G1355gat));
endmodule


