//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT3), .A3(G104), .ZN(new_n192));
  AOI22_X1  g006(.A1(new_n190), .A2(new_n192), .B1(new_n189), .B2(G107), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n187), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(G107), .ZN(new_n196));
  INV_X1    g010(.A(new_n192), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT3), .B1(new_n191), .B2(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n196), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT2), .B(G113), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G116), .ZN(new_n204));
  INV_X1    g018(.A(G116), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT72), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n204), .B2(new_n206), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n202), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(new_n206), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n211), .A2(new_n202), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n199), .A2(new_n187), .A3(G101), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n201), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n194), .B(new_n196), .C1(new_n197), .C2(new_n198), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT83), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n191), .B2(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n191), .A2(G104), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n189), .A2(KEYINPUT83), .A3(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G101), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n205), .A2(G119), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n203), .A2(G116), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT72), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(KEYINPUT5), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G113), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT5), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n229), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n223), .A2(new_n232), .A3(new_n212), .ZN(new_n233));
  XOR2_X1   g047(.A(G110), .B(G122), .Z(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n215), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n215), .B2(new_n233), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n238), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT86), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G146), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  INV_X1    g060(.A(G146), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n246), .A2(new_n247), .A3(G143), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT64), .B1(new_n243), .B2(G146), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT65), .B1(new_n247), .B2(G143), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n243), .A3(G146), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n244), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n250), .A2(new_n254), .B1(new_n258), .B2(new_n252), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  OR2_X1    g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n255), .A2(new_n257), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT70), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n262), .A2(G128), .A3(new_n245), .A4(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n258), .A2(KEYINPUT71), .A3(G128), .A4(new_n267), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G128), .B1(new_n267), .B2(new_n244), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n250), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n261), .B1(new_n275), .B2(G125), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G224), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(KEYINPUT87), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n276), .B(new_n279), .Z(new_n280));
  NAND2_X1  g094(.A1(new_n215), .A2(new_n233), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n234), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n215), .A2(new_n233), .A3(new_n235), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(KEYINPUT6), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT86), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n242), .A2(new_n280), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n279), .A2(KEYINPUT7), .ZN(new_n289));
  OR2_X1    g103(.A1(new_n276), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n223), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n212), .A3(new_n232), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n234), .B(KEYINPUT8), .Z(new_n293));
  OAI21_X1  g107(.A(new_n231), .B1(new_n230), .B2(new_n211), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(new_n212), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n292), .B(new_n293), .C1(new_n291), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n276), .A2(new_n289), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n290), .A2(new_n283), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n287), .A2(new_n288), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G210), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT88), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT88), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n299), .A2(new_n304), .A3(new_n301), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n287), .A2(new_n288), .A3(new_n300), .A4(new_n298), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT89), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n285), .B1(new_n284), .B2(new_n240), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n236), .A2(new_n237), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT86), .B1(new_n309), .B2(KEYINPUT6), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(G902), .B1(new_n311), .B2(new_n280), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT89), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n300), .A4(new_n298), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n303), .A2(new_n305), .B1(new_n307), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n277), .A2(G952), .ZN(new_n316));
  INV_X1    g130(.A(G234), .ZN(new_n317));
  INV_X1    g131(.A(G237), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI211_X1 g134(.A(new_n288), .B(new_n277), .C1(G234), .C2(G237), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT21), .B(G898), .Z(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G214), .B1(G237), .B2(G902), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n326), .B(KEYINPUT85), .Z(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G237), .A2(G953), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G214), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT90), .A3(new_n243), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n243), .A2(KEYINPUT90), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(G214), .A3(new_n329), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G131), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT17), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n333), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G131), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT16), .ZN(new_n341));
  NAND2_X1  g155(.A1(KEYINPUT77), .A2(G125), .ZN(new_n342));
  INV_X1    g156(.A(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(KEYINPUT77), .A2(G125), .A3(G140), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n341), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n260), .A2(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n341), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT78), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n348), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G146), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n348), .B(new_n247), .C1(new_n346), .C2(new_n351), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n338), .A2(KEYINPUT17), .A3(G131), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n340), .A2(new_n353), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT92), .ZN(new_n357));
  INV_X1    g171(.A(new_n345), .ZN(new_n358));
  AOI21_X1  g172(.A(G140), .B1(KEYINPUT77), .B2(G125), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n344), .A2(KEYINPUT92), .A3(new_n345), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G146), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT93), .ZN(new_n364));
  XNOR2_X1  g178(.A(G125), .B(G140), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n343), .A2(G125), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT80), .B1(new_n349), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n247), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT93), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n362), .A2(new_n372), .A3(G146), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n364), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT18), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n375), .A2(new_n335), .A3(KEYINPUT91), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n334), .B(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n356), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G113), .B(G122), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(new_n189), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n379), .B(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G475), .B1(new_n382), .B2(G902), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n356), .A2(new_n378), .A3(new_n381), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT19), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n367), .A2(new_n369), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT19), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n247), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT94), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n336), .A2(new_n339), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(KEYINPUT94), .A3(new_n247), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n392), .A2(new_n353), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n395), .A2(new_n378), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n385), .B1(new_n396), .B2(new_n381), .ZN(new_n397));
  NOR2_X1   g211(.A1(G475), .A2(G902), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n384), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n381), .B1(new_n395), .B2(new_n378), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n356), .A2(new_n378), .A3(new_n381), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n384), .B(new_n398), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n383), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n205), .A2(G122), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n205), .A2(G122), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n406), .A2(KEYINPUT95), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(KEYINPUT95), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(G107), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n409), .A2(new_n191), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT96), .B1(new_n243), .B2(G128), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT96), .ZN(new_n414));
  INV_X1    g228(.A(G128), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(G143), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT13), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G134), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n413), .A2(new_n416), .B1(G128), .B2(new_n243), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  OAI22_X1  g236(.A1(new_n411), .A2(new_n412), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n405), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n191), .B1(new_n424), .B2(KEYINPUT14), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n410), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n424), .A2(KEYINPUT14), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n409), .B1(new_n191), .B2(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n420), .A2(new_n418), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n420), .A2(new_n418), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n426), .B(new_n428), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT9), .B(G234), .Z(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(G217), .A3(new_n277), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n423), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n423), .B2(new_n431), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n288), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G478), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(KEYINPUT15), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n438), .B(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n404), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n315), .A2(new_n328), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G119), .B(G128), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT76), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT24), .B(G110), .Z(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n203), .A2(G128), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n449), .A2(KEYINPUT23), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n203), .A2(G128), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(KEYINPUT23), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(G110), .ZN(new_n454));
  OR3_X1    g268(.A1(new_n448), .A2(new_n454), .A3(KEYINPUT79), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT79), .B1(new_n448), .B2(new_n454), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n353), .A4(new_n371), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n353), .A2(new_n354), .B1(new_n446), .B2(new_n447), .ZN(new_n458));
  INV_X1    g272(.A(G110), .ZN(new_n459));
  INV_X1    g273(.A(new_n453), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT22), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(G137), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n457), .A2(new_n461), .A3(new_n465), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n288), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT81), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT25), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G217), .B1(new_n317), .B2(G902), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT75), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n467), .A2(new_n468), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n474), .A2(G902), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(KEYINPUT67), .A2(G137), .ZN(new_n481));
  NOR2_X1   g295(.A1(KEYINPUT67), .A2(G137), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n481), .A2(new_n482), .A3(G134), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(new_n418), .B2(G137), .ZN(new_n485));
  INV_X1    g299(.A(G137), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(KEYINPUT68), .A3(G134), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(KEYINPUT69), .B(G131), .C1(new_n483), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT11), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n418), .B2(G137), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT66), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(KEYINPUT11), .A2(G134), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n495), .B1(new_n481), .B2(new_n482), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n486), .A2(G134), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(KEYINPUT66), .B(new_n491), .C1(new_n418), .C2(G137), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n494), .A2(new_n496), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT69), .B1(new_n500), .B2(G131), .ZN(new_n501));
  OR3_X1    g315(.A1(new_n481), .A2(new_n482), .A3(G134), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n485), .A2(new_n487), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n335), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n490), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n275), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n500), .A2(G131), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT67), .B(G137), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n497), .B1(new_n509), .B2(new_n495), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n510), .A2(new_n335), .A3(new_n494), .A4(new_n499), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n259), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n507), .A2(KEYINPUT30), .A3(new_n513), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n213), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n329), .A2(G210), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n519), .B(KEYINPUT27), .Z(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT26), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(new_n194), .ZN(new_n522));
  INV_X1    g336(.A(new_n213), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n507), .A2(new_n513), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT31), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT28), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n270), .A2(new_n271), .B1(new_n250), .B2(new_n273), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n504), .B1(new_n511), .B2(KEYINPUT69), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n529), .A2(new_n530), .A3(new_n490), .ZN(new_n531));
  INV_X1    g345(.A(new_n513), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n213), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n507), .A2(KEYINPUT28), .A3(new_n513), .A4(new_n523), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n528), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n522), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT31), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n518), .A2(new_n538), .A3(new_n522), .A4(new_n524), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n526), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(G472), .A2(G902), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n540), .A2(KEYINPUT32), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT32), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT73), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n533), .A2(new_n545), .A3(new_n524), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n514), .A2(KEYINPUT73), .A3(new_n213), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(KEYINPUT28), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT74), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n528), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n546), .A2(new_n549), .A3(KEYINPUT28), .A4(new_n547), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n551), .A2(KEYINPUT29), .A3(new_n522), .A4(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n528), .A2(new_n522), .A3(new_n533), .A4(new_n534), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT29), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n507), .A2(KEYINPUT30), .A3(new_n513), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT30), .B1(new_n507), .B2(new_n513), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n557), .A2(new_n558), .A3(new_n523), .ZN(new_n559));
  INV_X1    g373(.A(new_n524), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n536), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(G902), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n553), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G472), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n480), .B1(new_n544), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n432), .ZN(new_n566));
  OAI21_X1  g380(.A(G221), .B1(new_n566), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G469), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n275), .A2(KEYINPUT10), .A3(new_n223), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT10), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n258), .B1(G128), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n270), .B2(new_n271), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n571), .B1(new_n574), .B2(new_n291), .ZN(new_n575));
  INV_X1    g389(.A(new_n512), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n201), .A2(new_n259), .A3(new_n214), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n570), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(G110), .B(G140), .ZN(new_n579));
  INV_X1    g393(.A(G227), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G953), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n579), .B(new_n581), .Z(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n275), .A2(new_n223), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n574), .A2(new_n291), .ZN(new_n585));
  OAI211_X1 g399(.A(KEYINPUT12), .B(new_n512), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n512), .B1(new_n584), .B2(new_n585), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT12), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n583), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n570), .A2(new_n575), .A3(new_n577), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n512), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n582), .B1(new_n592), .B2(new_n578), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n569), .B(new_n288), .C1(new_n590), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT84), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n578), .ZN(new_n596));
  INV_X1    g410(.A(new_n582), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n586), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n529), .A2(new_n291), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n291), .B2(new_n574), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT12), .B1(new_n601), .B2(new_n512), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n578), .B(new_n582), .C1(new_n599), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT84), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n569), .A4(new_n288), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n595), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n578), .B1(new_n599), .B2(new_n602), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n582), .B(KEYINPUT82), .Z(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n583), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n608), .A2(new_n610), .B1(new_n611), .B2(new_n592), .ZN(new_n612));
  OAI21_X1  g426(.A(G469), .B1(new_n612), .B2(G902), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n568), .B1(new_n607), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n444), .A2(new_n565), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n617));
  INV_X1    g431(.A(G472), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n540), .A2(new_n288), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n620), .B1(new_n540), .B2(new_n288), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n476), .A2(new_n479), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n624), .A2(new_n625), .A3(new_n614), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT98), .ZN(new_n627));
  INV_X1    g441(.A(new_n326), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n302), .B2(new_n306), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n438), .A2(new_n439), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n436), .B2(new_n437), .ZN(new_n632));
  INV_X1    g446(.A(new_n437), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(KEYINPUT33), .A3(new_n435), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n288), .A2(G478), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n630), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n404), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n629), .A2(new_n325), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  NOR2_X1   g456(.A1(new_n400), .A2(new_n401), .ZN(new_n643));
  INV_X1    g457(.A(new_n398), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT20), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n402), .ZN(new_n647));
  OAI211_X1 g461(.A(KEYINPUT99), .B(KEYINPUT20), .C1(new_n643), .C2(new_n644), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n647), .A2(new_n441), .A3(new_n383), .A4(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n629), .A2(new_n325), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n627), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  INV_X1    g468(.A(new_n623), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n466), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT100), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(new_n462), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n478), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n476), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n655), .A2(new_n660), .A3(new_n621), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n624), .A2(KEYINPUT101), .A3(new_n660), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n444), .A2(new_n663), .A3(new_n664), .A4(new_n614), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT37), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n459), .ZN(G12));
  AND2_X1   g481(.A1(new_n476), .A2(new_n659), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n544), .B2(new_n564), .ZN(new_n669));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n321), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n319), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n649), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n629), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n629), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT102), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n669), .A2(new_n614), .A3(new_n676), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  NAND2_X1  g494(.A1(new_n303), .A2(new_n305), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n314), .A2(new_n307), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT103), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n315), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n684), .A2(KEYINPUT38), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT38), .B1(new_n684), .B2(new_n686), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n540), .A2(new_n541), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT32), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n540), .A2(KEYINPUT32), .A3(new_n541), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n518), .A2(new_n524), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n522), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n546), .A2(new_n547), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n695), .B(new_n288), .C1(new_n522), .C2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(G472), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n692), .A2(new_n693), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n404), .ZN(new_n700));
  INV_X1    g514(.A(new_n441), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n476), .A2(new_n326), .A3(new_n659), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n689), .A2(KEYINPUT104), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n704), .B1(new_n687), .B2(new_n688), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n672), .B(KEYINPUT39), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n614), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n710), .B(KEYINPUT40), .Z(new_n711));
  NAND3_X1  g525(.A1(new_n705), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NAND3_X1  g527(.A1(new_n404), .A2(new_n637), .A3(new_n672), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n404), .A2(KEYINPUT105), .A3(new_n637), .A4(new_n672), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n629), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT106), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n716), .A2(new_n629), .A3(new_n720), .A4(new_n717), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n669), .A2(new_n719), .A3(new_n614), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  NAND2_X1  g537(.A1(new_n604), .A2(new_n288), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n595), .A2(new_n606), .B1(G469), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n567), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n564), .A2(new_n692), .A3(new_n693), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n639), .A2(new_n727), .A3(new_n728), .A4(new_n625), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND4_X1  g545(.A1(new_n651), .A2(new_n727), .A3(new_n728), .A4(new_n625), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  AND4_X1   g547(.A1(new_n567), .A2(new_n629), .A3(new_n725), .A4(new_n325), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n669), .A2(new_n442), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  INV_X1    g550(.A(new_n541), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n551), .A2(new_n552), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n536), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n526), .A2(new_n539), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n540), .A2(new_n288), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G472), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n742), .A2(KEYINPUT107), .A3(G472), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n741), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n629), .A2(new_n702), .A3(new_n325), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n625), .A3(new_n727), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT108), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n739), .A2(new_n740), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n541), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT107), .B1(new_n742), .B2(G472), .ZN(new_n753));
  AOI211_X1 g567(.A(new_n744), .B(new_n618), .C1(new_n540), .C2(new_n288), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n625), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n726), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n748), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  NAND2_X1  g574(.A1(new_n716), .A2(new_n717), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n629), .A2(new_n725), .A3(new_n567), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n747), .A2(new_n660), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G125), .ZN(G27));
  NAND3_X1  g579(.A1(new_n681), .A2(new_n326), .A3(new_n682), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n607), .A2(new_n613), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n567), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n770));
  NOR2_X1   g584(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n769), .A2(new_n565), .A3(new_n762), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n728), .A2(new_n625), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n614), .A2(new_n326), .A3(new_n681), .A4(new_n682), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n775), .A2(new_n776), .A3(new_n761), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n774), .B1(new_n777), .B2(new_n770), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G131), .ZN(G33));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n674), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT110), .B1(new_n649), .B2(new_n673), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n769), .A2(new_n565), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND2_X1  g598(.A1(new_n700), .A2(new_n637), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT43), .Z(new_n786));
  OAI211_X1 g600(.A(new_n786), .B(new_n660), .C1(new_n622), .C2(new_n623), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n766), .B1(new_n788), .B2(KEYINPUT44), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n612), .A2(KEYINPUT45), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n611), .A2(new_n592), .ZN(new_n791));
  INV_X1    g605(.A(new_n578), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n589), .B2(new_n586), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n791), .B1(new_n793), .B2(new_n609), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n790), .A2(new_n796), .A3(G469), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT111), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n790), .A2(new_n796), .A3(new_n799), .A4(G469), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(G469), .A2(G902), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n798), .A2(new_n800), .B1(G469), .B2(G902), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT46), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n607), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n567), .A3(new_n709), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n789), .B(new_n810), .C1(KEYINPUT44), .C2(new_n788), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G137), .ZN(G39));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  INV_X1    g627(.A(new_n807), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n607), .B1(new_n806), .B2(KEYINPUT46), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n813), .B(new_n567), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n813), .B1(new_n808), .B2(new_n567), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n766), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n728), .A2(new_n625), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n819), .A2(new_n762), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G140), .ZN(G42));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n786), .A2(new_n320), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n756), .A3(new_n628), .ZN(new_n827));
  OR3_X1    g641(.A1(new_n689), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n825), .B1(new_n689), .B2(new_n827), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n828), .A2(KEYINPUT118), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n755), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n826), .A2(new_n820), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n725), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n567), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n835), .B(new_n837), .C1(new_n819), .C2(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n660), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n841));
  OR3_X1    g655(.A1(new_n836), .A2(new_n726), .A3(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n766), .A2(new_n699), .A3(new_n726), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n625), .A3(new_n320), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n844), .A2(new_n404), .A3(new_n637), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n840), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n824), .B1(new_n834), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n840), .A2(new_n842), .A3(new_n845), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(KEYINPUT119), .A3(KEYINPUT51), .A4(new_n830), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n840), .A2(KEYINPUT51), .A3(new_n842), .A4(new_n845), .ZN(new_n851));
  INV_X1    g665(.A(new_n830), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n836), .A2(new_n775), .A3(new_n726), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(KEYINPUT48), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n826), .A2(new_n756), .A3(new_n629), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(KEYINPUT48), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n316), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n847), .A2(new_n849), .A3(new_n853), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n735), .A2(new_n729), .A3(new_n732), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n759), .A2(new_n778), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n328), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n299), .A2(new_n304), .A3(new_n301), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n304), .B1(new_n299), .B2(new_n301), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n306), .B(new_n313), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n863), .B(new_n638), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT112), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT112), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n683), .A2(new_n870), .A3(new_n863), .A4(new_n638), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n626), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n404), .A2(new_n701), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n315), .A2(new_n328), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n626), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n872), .A2(new_n665), .A3(new_n615), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n441), .A2(new_n673), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n383), .A2(new_n878), .A3(new_n648), .A4(new_n647), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n728), .A2(new_n660), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n841), .B2(new_n761), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n769), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n783), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n862), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n735), .A2(new_n729), .A3(new_n732), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n758), .B2(new_n750), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n860), .B1(new_n887), .B2(new_n778), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT113), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n302), .A2(new_n306), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n614), .A2(new_n672), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n704), .A2(new_n891), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n699), .A2(new_n703), .A3(new_n892), .A4(new_n702), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT113), .B1(new_n896), .B2(new_n893), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n722), .A2(new_n679), .A3(new_n764), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT52), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT52), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n895), .A2(new_n897), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n722), .A2(new_n679), .A3(new_n764), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n900), .A2(KEYINPUT114), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT114), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n906), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n759), .A2(new_n778), .A3(new_n861), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n909), .A2(new_n877), .A3(new_n883), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n900), .A2(new_n904), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g726(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n890), .A2(new_n908), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n912), .A2(new_n914), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n910), .A2(new_n907), .A3(new_n905), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n889), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT116), .B1(new_n920), .B2(new_n916), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n889), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n912), .B2(new_n914), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT116), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT54), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n859), .A2(new_n917), .A3(new_n921), .A4(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n638), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n844), .A2(new_n927), .ZN(new_n928));
  OAI22_X1  g742(.A1(new_n926), .A2(new_n928), .B1(G952), .B2(G953), .ZN(new_n929));
  INV_X1    g743(.A(new_n689), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n725), .B(KEYINPUT49), .Z(new_n931));
  NOR4_X1   g745(.A1(new_n931), .A2(new_n480), .A3(new_n699), .A4(new_n785), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n930), .A2(new_n567), .A3(new_n327), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n929), .A2(new_n933), .ZN(G75));
  XOR2_X1   g748(.A(new_n311), .B(new_n280), .Z(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT120), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n915), .A2(new_n288), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(G210), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n277), .A2(G952), .ZN(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n939), .A2(new_n937), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n939), .A2(KEYINPUT122), .A3(new_n937), .A4(new_n943), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n941), .B(new_n942), .C1(new_n946), .C2(new_n947), .ZN(G51));
  AND2_X1   g762(.A1(new_n862), .A2(new_n884), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n889), .B1(new_n909), .B2(KEYINPUT117), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(new_n907), .A3(new_n950), .A4(new_n905), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT52), .B1(new_n898), .B2(new_n899), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n902), .A2(new_n903), .A3(new_n901), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n877), .ZN(new_n955));
  INV_X1    g769(.A(new_n883), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n887), .A2(new_n955), .A3(new_n956), .A4(new_n778), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n914), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n951), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n916), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n802), .B(KEYINPUT57), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n604), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n938), .A2(new_n800), .A3(new_n798), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n942), .B1(new_n962), .B2(new_n963), .ZN(G54));
  NAND3_X1  g778(.A1(new_n938), .A2(KEYINPUT58), .A3(G475), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n965), .A2(new_n643), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n643), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n942), .ZN(G60));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT59), .Z(new_n970));
  NOR3_X1   g784(.A1(new_n960), .A2(new_n635), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n921), .A2(new_n917), .A3(new_n925), .ZN(new_n972));
  INV_X1    g786(.A(new_n970), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n942), .B(new_n971), .C1(new_n974), .C2(new_n635), .ZN(G63));
  INV_X1    g789(.A(new_n477), .ZN(new_n976));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT60), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n976), .B1(new_n915), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n942), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n978), .B1(new_n951), .B2(new_n958), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n658), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n979), .A2(KEYINPUT61), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n984));
  AOI21_X1  g798(.A(KEYINPUT123), .B1(new_n979), .B2(new_n980), .ZN(new_n985));
  OAI211_X1 g799(.A(KEYINPUT123), .B(new_n980), .C1(new_n981), .C2(new_n477), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n982), .ZN(new_n987));
  OAI211_X1 g801(.A(KEYINPUT124), .B(new_n984), .C1(new_n985), .C2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n980), .B1(new_n981), .B2(new_n477), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT123), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n986), .A3(new_n982), .ZN(new_n993));
  AOI21_X1  g807(.A(KEYINPUT124), .B1(new_n993), .B2(new_n984), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n983), .B1(new_n989), .B2(new_n994), .ZN(G66));
  AOI21_X1  g809(.A(new_n277), .B1(new_n322), .B2(G224), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n955), .A2(new_n887), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(new_n277), .ZN(new_n998));
  OAI22_X1  g812(.A1(new_n308), .A2(new_n310), .B1(G898), .B2(new_n277), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n998), .B(new_n999), .Z(G69));
  NAND2_X1  g814(.A1(new_n516), .A2(new_n517), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(new_n389), .Z(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n822), .A2(new_n899), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n810), .A2(new_n565), .A3(new_n629), .A4(new_n702), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n811), .A2(new_n1005), .A3(new_n778), .A4(new_n783), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n1004), .A2(new_n1006), .A3(G953), .ZN(new_n1007));
  AOI211_X1 g821(.A(new_n1003), .B(new_n1007), .C1(G900), .C2(G953), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1002), .B(KEYINPUT125), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n903), .B1(new_n1010), .B2(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n712), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  AOI211_X1 g828(.A(new_n766), .B(new_n710), .C1(new_n927), .C2(new_n874), .ZN(new_n1015));
  AOI22_X1  g829(.A1(new_n1012), .A2(new_n1014), .B1(new_n565), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n712), .A2(new_n1013), .A3(new_n1011), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1016), .A2(new_n811), .A3(new_n822), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1009), .B1(new_n1018), .B2(new_n277), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1008), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(G953), .B1(new_n580), .B2(new_n670), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1020), .B(new_n1021), .ZN(G72));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n1018), .B2(new_n997), .ZN(new_n1025));
  INV_X1    g839(.A(new_n695), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n942), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n694), .A2(new_n522), .ZN(new_n1028));
  NOR3_X1   g842(.A1(new_n1004), .A2(new_n1006), .A3(new_n997), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1024), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n1026), .A2(new_n1030), .A3(new_n1028), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n923), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1027), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(KEYINPUT127), .ZN(new_n1035));
  INV_X1    g849(.A(KEYINPUT127), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n1027), .A2(new_n1036), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1035), .A2(new_n1037), .ZN(G57));
endmodule


