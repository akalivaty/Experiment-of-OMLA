//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G107), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT68), .B(G116), .ZN(new_n189));
  INV_X1    g003(.A(G122), .ZN(new_n190));
  NOR3_X1   g004(.A1(new_n189), .A2(KEYINPUT14), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT94), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n189), .B2(new_n190), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G116), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(KEYINPUT94), .A3(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n191), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT95), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT66), .A2(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT93), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n201), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(new_n202), .B2(new_n203), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT93), .B1(new_n211), .B2(new_n207), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n209), .A2(G134), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(G134), .B1(new_n209), .B2(new_n212), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n193), .B(KEYINPUT95), .C1(new_n191), .C2(new_n196), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n195), .B1(new_n189), .B2(new_n190), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n217), .A2(G107), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n199), .A2(new_n215), .A3(new_n216), .A4(new_n218), .ZN(new_n219));
  XOR2_X1   g033(.A(KEYINPUT9), .B(G234), .Z(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G217), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n205), .A2(new_n208), .ZN(new_n224));
  OAI21_X1  g038(.A(G134), .B1(new_n211), .B2(KEYINPUT13), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n217), .B(G107), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n219), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n223), .B1(new_n219), .B2(new_n228), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n187), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT96), .ZN(new_n232));
  INV_X1    g046(.A(G478), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(KEYINPUT15), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT96), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n235), .B(new_n187), .C1(new_n229), .C2(new_n230), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT97), .B1(new_n231), .B2(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n232), .A2(KEYINPUT97), .A3(new_n234), .A4(new_n236), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G952), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G953), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(G234), .B2(G237), .ZN(new_n246));
  AOI211_X1 g060(.A(new_n187), .B(new_n221), .C1(G234), .C2(G237), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT21), .B(G898), .Z(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n246), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(G214), .B1(G237), .B2(G902), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT2), .B(G113), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G119), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(KEYINPUT68), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n262), .B2(G119), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n256), .B1(new_n263), .B2(KEYINPUT67), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n265));
  INV_X1    g079(.A(G119), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n259), .B2(new_n261), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n265), .B(new_n255), .C1(new_n267), .C2(new_n258), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G104), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G107), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT80), .ZN(new_n272));
  OAI22_X1  g086(.A1(new_n272), .A2(KEYINPUT3), .B1(new_n270), .B2(G107), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n188), .A2(G104), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n271), .B(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G101), .ZN(new_n277));
  INV_X1    g091(.A(new_n275), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(KEYINPUT80), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G101), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n271), .A4(new_n273), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n277), .A2(new_n284), .A3(KEYINPUT4), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n276), .A2(new_n286), .A3(G101), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n269), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n271), .A2(new_n275), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G101), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n276), .B2(G101), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n263), .A2(new_n256), .ZN(new_n293));
  INV_X1    g107(.A(G113), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(new_n258), .ZN(new_n296));
  INV_X1    g110(.A(new_n258), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n189), .B2(new_n266), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n296), .B1(new_n298), .B2(new_n295), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n292), .A2(new_n293), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(G110), .B(G122), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n288), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT87), .ZN(new_n303));
  INV_X1    g117(.A(G224), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n303), .B1(new_n304), .B2(G953), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n221), .A2(KEYINPUT87), .A3(G224), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(KEYINPUT7), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n308));
  INV_X1    g122(.A(G146), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G143), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n210), .A2(G146), .ZN(new_n311));
  AND4_X1   g125(.A1(new_n308), .A2(new_n310), .A3(new_n311), .A4(G128), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT64), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n313), .B1(new_n210), .B2(G146), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n309), .A2(KEYINPUT64), .A3(G143), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT65), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n210), .B2(G146), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n309), .A2(KEYINPUT65), .A3(G143), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n314), .B(new_n315), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT1), .B1(new_n210), .B2(G146), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n202), .A3(new_n203), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n312), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AND4_X1   g139(.A1(KEYINPUT0), .A2(new_n310), .A3(new_n311), .A4(G128), .ZN(new_n326));
  XOR2_X1   g140(.A(KEYINPUT0), .B(G128), .Z(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n319), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(new_n323), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n307), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n291), .A2(new_n293), .A3(new_n299), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n301), .B(KEYINPUT8), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n333), .A2(new_n296), .B1(new_n263), .B2(new_n256), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n331), .B(new_n332), .C1(new_n334), .C2(new_n291), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n328), .A2(new_n323), .ZN(new_n336));
  INV_X1    g150(.A(new_n307), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(new_n324), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n302), .A2(new_n330), .A3(new_n335), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n187), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT88), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n288), .A2(new_n300), .ZN(new_n342));
  INV_X1    g156(.A(new_n301), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(KEYINPUT6), .A3(new_n302), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n346), .A3(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n336), .A2(new_n324), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n305), .A2(new_n306), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT86), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n348), .B(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT88), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n339), .A2(new_n353), .A3(new_n187), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT89), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(G210), .B1(G237), .B2(G902), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT90), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n341), .A2(new_n352), .A3(KEYINPUT89), .A4(new_n354), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n341), .A2(new_n352), .A3(new_n358), .A4(new_n354), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n254), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G140), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT16), .B1(new_n365), .B2(G125), .ZN(new_n366));
  AND2_X1   g180(.A1(KEYINPUT74), .A2(G140), .ZN(new_n367));
  NOR2_X1   g181(.A1(KEYINPUT74), .A2(G140), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT75), .B(G125), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  OR2_X1    g183(.A1(KEYINPUT74), .A2(G140), .ZN(new_n370));
  NAND2_X1  g184(.A1(KEYINPUT74), .A2(G140), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n323), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT75), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n323), .B2(G140), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n369), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n366), .B1(new_n375), .B2(KEYINPUT16), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n309), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT16), .ZN(new_n378));
  OAI21_X1  g192(.A(G125), .B1(new_n367), .B2(new_n368), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n323), .A2(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT75), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n378), .B1(new_n382), .B2(new_n369), .ZN(new_n383));
  OAI21_X1  g197(.A(G146), .B1(new_n383), .B2(new_n366), .ZN(new_n384));
  INV_X1    g198(.A(G237), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n221), .A3(G214), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n210), .ZN(new_n387));
  NOR2_X1   g201(.A1(G237), .A2(G953), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(G143), .A3(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT17), .A3(G131), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(G131), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT17), .ZN(new_n393));
  INV_X1    g207(.A(G131), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n387), .A2(new_n394), .A3(new_n389), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n377), .A2(new_n384), .A3(new_n391), .A4(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G113), .B(G122), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT92), .B(G104), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT18), .A2(G131), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n390), .B(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n309), .B1(new_n382), .B2(new_n369), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n365), .A2(G125), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n380), .A2(new_n405), .A3(new_n309), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n403), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n397), .A2(new_n401), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n401), .B1(new_n397), .B2(new_n408), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n187), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G475), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G475), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n392), .A2(new_n395), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n375), .A2(KEYINPUT19), .ZN(new_n416));
  OR2_X1    g230(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n417));
  NAND2_X1  g231(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n417), .A2(new_n380), .A3(new_n405), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n384), .B(new_n415), .C1(new_n420), .C2(G146), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n401), .B1(new_n421), .B2(new_n408), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n414), .B(new_n187), .C1(new_n409), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT20), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n415), .B1(new_n376), .B2(new_n309), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n416), .A2(new_n309), .A3(new_n419), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n408), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n400), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n397), .A2(new_n401), .A3(new_n408), .ZN(new_n429));
  AOI21_X1  g243(.A(G475), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n431), .A3(new_n187), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n413), .B1(new_n424), .B2(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n242), .A2(new_n364), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT69), .ZN(new_n435));
  INV_X1    g249(.A(new_n268), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n255), .B1(new_n298), .B2(new_n265), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT11), .ZN(new_n439));
  INV_X1    g253(.A(G134), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(G137), .ZN(new_n441));
  INV_X1    g255(.A(G137), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(KEYINPUT11), .A3(G134), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(G137), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G131), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n441), .A2(new_n443), .A3(new_n394), .A4(new_n444), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n328), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n440), .A2(G137), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n442), .A2(G134), .ZN(new_n451));
  OAI21_X1  g265(.A(G131), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n314), .A2(new_n315), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT65), .B1(new_n309), .B2(G143), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n316), .A2(new_n210), .A3(G146), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n204), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n455), .A2(new_n458), .B1(new_n459), .B2(new_n320), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n453), .B1(new_n460), .B2(new_n312), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n268), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n438), .A2(new_n449), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT70), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n456), .A2(new_n457), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n321), .B1(new_n466), .B2(new_n454), .ZN(new_n467));
  INV_X1    g281(.A(new_n312), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n469), .A2(new_n453), .B1(new_n328), .B2(new_n448), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n470), .A2(KEYINPUT70), .A3(new_n462), .A4(new_n438), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n268), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT69), .B1(new_n264), .B2(new_n268), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n472), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT28), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT28), .B1(new_n475), .B2(new_n470), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n388), .A2(G210), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(new_n283), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n481), .B(new_n482), .Z(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT29), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n477), .A2(new_n479), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n470), .B1(new_n268), .B2(new_n264), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT70), .B1(new_n475), .B2(new_n470), .ZN(new_n490));
  AND4_X1   g304(.A1(KEYINPUT70), .A2(new_n470), .A3(new_n462), .A4(new_n438), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT71), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT28), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n478), .A2(new_n493), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n488), .B1(new_n465), .B2(new_n471), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT28), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n484), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n461), .A2(new_n449), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n470), .A2(KEYINPUT30), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(new_n269), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n472), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n484), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n485), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n187), .B(new_n487), .C1(new_n499), .C2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT72), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n508), .A2(new_n509), .A3(G472), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n508), .B2(G472), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT32), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n494), .A2(new_n498), .A3(new_n484), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n472), .A2(new_n483), .A3(new_n504), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT31), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n472), .A2(KEYINPUT31), .A3(new_n483), .A4(new_n504), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(G902), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G472), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n512), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n513), .A2(new_n518), .ZN(new_n522));
  AND4_X1   g336(.A1(new_n512), .A2(new_n522), .A3(new_n520), .A4(new_n187), .ZN(new_n523));
  OAI22_X1  g337(.A1(new_n510), .A2(new_n511), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT25), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT22), .B(G137), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n526), .B(new_n527), .Z(new_n528));
  AOI21_X1  g342(.A(new_n266), .B1(new_n202), .B2(new_n203), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n201), .A2(G119), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g345(.A(KEYINPUT24), .B(G110), .Z(new_n532));
  OAI21_X1  g346(.A(KEYINPUT76), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n534));
  AND2_X1   g348(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n535));
  NOR2_X1   g349(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n536));
  OAI22_X1  g350(.A1(new_n535), .A2(new_n536), .B1(new_n266), .B2(G128), .ZN(new_n537));
  INV_X1    g351(.A(G110), .ZN(new_n538));
  INV_X1    g352(.A(new_n530), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n534), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n532), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT76), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n541), .B(new_n542), .C1(new_n530), .C2(new_n529), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n533), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n384), .A3(new_n406), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n534), .A2(new_n537), .A3(new_n539), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G110), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n531), .A2(new_n532), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n377), .B2(new_n384), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT77), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n377), .A2(new_n384), .ZN(new_n553));
  INV_X1    g367(.A(new_n550), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT77), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n545), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n528), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n528), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n546), .A2(new_n551), .A3(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n558), .A2(G902), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n525), .B1(new_n561), .B2(KEYINPUT78), .ZN(new_n562));
  INV_X1    g376(.A(G217), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(G234), .B2(new_n187), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n546), .A2(new_n551), .A3(KEYINPUT77), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n556), .B1(new_n555), .B2(new_n545), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n559), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n560), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n187), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT78), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT25), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n562), .A2(new_n564), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n558), .A2(new_n560), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n564), .A2(G902), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT84), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n291), .A2(new_n322), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT82), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n310), .A2(new_n311), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n201), .B1(new_n310), .B2(KEYINPUT1), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n468), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n292), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT82), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n291), .A2(new_n322), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n580), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n588), .A2(KEYINPUT12), .A3(new_n448), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT12), .B1(new_n588), .B2(new_n448), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n578), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n448), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT12), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n588), .A2(KEYINPUT12), .A3(new_n448), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(KEYINPUT84), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n585), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n285), .A2(new_n328), .A3(new_n287), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n292), .A2(KEYINPUT10), .A3(new_n469), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n448), .B(KEYINPUT81), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n221), .A2(G227), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT79), .ZN(new_n604));
  XNOR2_X1  g418(.A(G110), .B(G140), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n591), .A2(new_n596), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n448), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n602), .ZN(new_n611));
  INV_X1    g425(.A(new_n606), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G469), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n615), .A3(new_n187), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n602), .B1(new_n589), .B2(new_n590), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT83), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(KEYINPUT83), .B(new_n602), .C1(new_n589), .C2(new_n590), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n612), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n607), .A2(new_n610), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(G469), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(G469), .A2(G902), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n616), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(G221), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n220), .B2(new_n187), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n434), .A2(new_n524), .A3(new_n577), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  INV_X1    g444(.A(new_n358), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n355), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n363), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n251), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT99), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n633), .A2(new_n636), .A3(new_n251), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n433), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n232), .A2(new_n233), .A3(new_n236), .ZN(new_n640));
  INV_X1    g454(.A(new_n230), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n219), .A2(new_n228), .A3(new_n223), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(KEYINPUT33), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n229), .B2(new_n230), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n643), .A2(new_n645), .A3(G478), .A4(new_n187), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n639), .A2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n638), .A2(new_n250), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(KEYINPUT98), .A2(G472), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n519), .B(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n627), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n572), .A2(new_n575), .A3(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n651), .A2(new_n625), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  NOR2_X1   g471(.A1(new_n638), .A2(new_n250), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n423), .A2(KEYINPUT20), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n431), .B1(new_n430), .B2(new_n187), .ZN(new_n660));
  OAI21_X1  g474(.A(KEYINPUT100), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n424), .A2(new_n432), .A3(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n661), .A2(new_n412), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n658), .A2(new_n654), .A3(new_n241), .A4(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NAND2_X1  g481(.A1(new_n552), .A2(new_n557), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n574), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n572), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n651), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n434), .A2(new_n673), .A3(new_n628), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n524), .A2(new_n628), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n636), .B1(new_n633), .B2(new_n251), .ZN(new_n679));
  AOI211_X1 g493(.A(KEYINPUT99), .B(new_n252), .C1(new_n632), .C2(new_n363), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n572), .A2(new_n671), .ZN(new_n682));
  INV_X1    g496(.A(new_n246), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n247), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n661), .A2(new_n412), .A3(new_n663), .A4(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n239), .B2(new_n240), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n681), .A2(new_n682), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n677), .B1(new_n678), .B2(new_n689), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n637), .A2(new_n688), .A3(new_n635), .A4(new_n682), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(KEYINPUT101), .A3(new_n524), .A4(new_n628), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  XOR2_X1   g508(.A(new_n686), .B(KEYINPUT39), .Z(new_n695));
  NOR3_X1   g509(.A1(new_n625), .A2(new_n627), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n514), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n484), .B2(new_n476), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n187), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  OAI21_X1  g518(.A(G472), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n523), .B2(new_n521), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n362), .A2(new_n363), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT38), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n362), .A2(KEYINPUT38), .A3(new_n363), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n241), .A2(new_n639), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n713), .A2(new_n252), .A3(new_n682), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n698), .A2(new_n706), .A3(new_n712), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  NOR3_X1   g530(.A1(new_n672), .A2(new_n679), .A3(new_n680), .ZN(new_n717));
  INV_X1    g531(.A(new_n686), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n648), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n717), .A2(new_n524), .A3(new_n628), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT104), .B(G146), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G48));
  INV_X1    g536(.A(new_n511), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n508), .A2(new_n509), .A3(G472), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n523), .A2(new_n521), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n576), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n614), .A2(new_n187), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n652), .A3(new_n616), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT105), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n615), .B1(new_n614), .B2(new_n187), .ZN(new_n732));
  AOI211_X1 g546(.A(G469), .B(G902), .C1(new_n608), .C2(new_n613), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n652), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n727), .A2(new_n649), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT41), .B(G113), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G15));
  INV_X1    g554(.A(new_n250), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n681), .A2(new_n241), .A3(new_n741), .A4(new_n664), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n743), .A2(new_n727), .A3(new_n737), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n257), .ZN(G18));
  NAND3_X1  g559(.A1(new_n524), .A2(new_n433), .A3(new_n242), .ZN(new_n746));
  INV_X1    g560(.A(new_n730), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n681), .A2(new_n747), .A3(new_n741), .A4(new_n682), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n266), .ZN(G21));
  AOI21_X1  g564(.A(new_n478), .B1(new_n476), .B2(KEYINPUT28), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n518), .B1(new_n751), .B2(new_n483), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n520), .A3(new_n187), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT106), .B(G472), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n753), .B1(new_n519), .B2(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n713), .A2(new_n755), .A3(new_n576), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n658), .A2(new_n756), .A3(new_n737), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  NOR3_X1   g572(.A1(new_n755), .A2(new_n648), .A3(new_n718), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n681), .A3(new_n682), .A4(new_n747), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  NAND3_X1  g575(.A1(new_n362), .A2(new_n363), .A3(new_n251), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n625), .A2(new_n762), .A3(new_n627), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n524), .A2(new_n763), .A3(new_n577), .A4(new_n719), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(KEYINPUT42), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n765), .A2(KEYINPUT42), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n766), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n727), .A2(new_n719), .A3(new_n763), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n727), .A2(new_n773), .A3(new_n688), .A4(new_n763), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n524), .A2(new_n763), .A3(new_n577), .A4(new_n688), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT108), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n647), .A2(new_n779), .A3(new_n433), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n779), .B1(new_n647), .B2(new_n433), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n651), .A3(new_n682), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT109), .Z(new_n786));
  INV_X1    g600(.A(new_n762), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n783), .A2(new_n784), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n621), .A2(new_n622), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n621), .A2(KEYINPUT45), .A3(new_n622), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(G469), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(KEYINPUT46), .A3(new_n624), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n616), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT46), .B1(new_n793), .B2(new_n624), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n652), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n695), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  NOR2_X1   g614(.A1(new_n797), .A2(KEYINPUT47), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT47), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT46), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n791), .A2(new_n792), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n803), .B(G469), .C1(new_n804), .C2(G902), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n616), .A3(new_n794), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n802), .B1(new_n806), .B2(new_n652), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n524), .A2(new_n762), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n576), .A3(new_n719), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n720), .A2(new_n760), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n690), .B2(new_n692), .ZN(new_n814));
  INV_X1    g628(.A(new_n706), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n682), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n638), .A2(new_n713), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n628), .A3(new_n817), .A4(new_n686), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n812), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n720), .A2(new_n760), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n812), .A2(new_n693), .A3(new_n820), .A4(new_n818), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT112), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n768), .A2(new_n770), .B1(new_n774), .B2(new_n776), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n639), .B1(new_n239), .B2(new_n240), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n824), .A2(new_n825), .A3(new_n364), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n825), .B1(new_n824), .B2(new_n364), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n654), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n757), .A2(new_n828), .A3(new_n629), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n744), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n648), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n654), .A2(new_n364), .A3(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n832), .B(new_n674), .C1(new_n748), .C2(new_n746), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n738), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n241), .B(new_n687), .C1(new_n725), .C2(new_n726), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n682), .B(new_n763), .C1(new_n835), .C2(new_n759), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n823), .A2(new_n830), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n693), .A2(new_n820), .A3(new_n818), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT52), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n693), .A2(new_n820), .A3(new_n818), .A4(new_n812), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n822), .A2(KEYINPUT53), .A3(new_n838), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  XNOR2_X1  g659(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n840), .A2(new_n842), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n847), .B2(new_n837), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n847), .A2(new_n837), .A3(new_n846), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n822), .A2(new_n838), .A3(new_n843), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(KEYINPUT114), .B(new_n849), .C1(new_n853), .C2(new_n845), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n755), .A2(new_n576), .A3(new_n683), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n252), .A3(new_n711), .A4(new_n782), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT50), .B1(new_n860), .B2(new_n730), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n734), .A2(new_n652), .A3(new_n246), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n706), .A2(new_n862), .A3(new_n762), .ZN(new_n863));
  INV_X1    g677(.A(new_n647), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n577), .A3(new_n433), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n862), .A2(new_n762), .ZN(new_n866));
  INV_X1    g680(.A(new_n755), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n682), .A3(new_n867), .A4(new_n782), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n861), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  OR3_X1    g683(.A1(new_n860), .A2(KEYINPUT50), .A3(new_n730), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n797), .A2(KEYINPUT47), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n806), .A2(new_n802), .A3(new_n652), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n729), .A2(new_n616), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT115), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n871), .A2(new_n872), .B1(new_n627), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n859), .A2(new_n782), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n787), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n869), .B(new_n870), .C1(new_n875), .C2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n874), .A2(new_n627), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n801), .B2(new_n807), .ZN(new_n882));
  INV_X1    g696(.A(new_n877), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(KEYINPUT51), .A3(new_n870), .A4(new_n869), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n876), .A2(new_n681), .A3(new_n747), .ZN(new_n886));
  AND4_X1   g700(.A1(new_n244), .A2(new_n880), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n727), .A2(new_n782), .A3(new_n866), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT48), .Z(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n863), .A2(new_n577), .A3(new_n831), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n887), .A2(new_n888), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n245), .B1(new_n878), .B2(new_n879), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(new_n892), .A3(new_n886), .A4(new_n885), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT116), .B1(new_n895), .B2(new_n890), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n858), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT117), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n243), .A2(new_n221), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n858), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NOR4_X1   g717(.A1(new_n653), .A2(new_n639), .A3(new_n864), .A4(new_n252), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT110), .Z(new_n905));
  AOI21_X1  g719(.A(new_n712), .B1(KEYINPUT49), .B2(new_n873), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n873), .A2(KEYINPUT49), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n905), .A2(new_n815), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n903), .A2(new_n908), .ZN(G75));
  NOR2_X1   g723(.A1(new_n221), .A2(G952), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n844), .A2(new_n848), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(G210), .A3(G902), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n345), .A2(new_n347), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(new_n351), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT55), .Z(new_n917));
  AOI21_X1  g731(.A(new_n910), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n187), .B1(new_n844), .B2(new_n848), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n360), .ZN(new_n921));
  INV_X1    g735(.A(new_n917), .ZN(new_n922));
  XOR2_X1   g736(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n923));
  AND4_X1   g737(.A1(new_n919), .A2(new_n921), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n917), .B1(new_n920), .B2(new_n360), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n919), .B1(new_n925), .B2(new_n923), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n918), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT120), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n929), .B(new_n918), .C1(new_n924), .C2(new_n926), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(G51));
  NAND2_X1  g745(.A1(new_n624), .A2(KEYINPUT57), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n624), .A2(KEYINPUT57), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n845), .B1(new_n844), .B2(new_n848), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n932), .B(new_n933), .C1(new_n855), .C2(new_n934), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n935), .A2(KEYINPUT121), .A3(new_n614), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT121), .B1(new_n935), .B2(new_n614), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n920), .A2(G469), .A3(new_n804), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n910), .B1(new_n938), .B2(new_n939), .ZN(G54));
  NAND3_X1  g754(.A1(new_n920), .A2(KEYINPUT58), .A3(G475), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n409), .A2(new_n422), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(new_n910), .ZN(G60));
  NAND2_X1  g758(.A1(new_n643), .A2(new_n645), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT122), .ZN(new_n946));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT59), .Z(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n858), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n910), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n855), .A2(new_n934), .ZN(new_n951));
  OR3_X1    g765(.A1(new_n951), .A2(new_n948), .A3(new_n946), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(G63));
  XNOR2_X1  g767(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n954));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n844), .B2(new_n848), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n910), .B1(new_n957), .B2(new_n670), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n573), .B2(new_n957), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g774(.A(G953), .B1(new_n249), .B2(new_n304), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n830), .A2(new_n834), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n961), .B1(new_n962), .B2(G953), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n915), .B1(G898), .B2(new_n221), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT124), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n963), .B(new_n965), .ZN(G69));
  XOR2_X1   g780(.A(new_n814), .B(KEYINPUT126), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n715), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT62), .Z(new_n969));
  AND2_X1   g783(.A1(new_n799), .A2(new_n810), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n831), .A2(new_n824), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n695), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n727), .A2(new_n763), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n969), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n502), .A2(new_n503), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT125), .Z(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(new_n420), .Z(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n974), .A2(new_n221), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(G227), .A2(G900), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(G953), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n798), .A2(new_n727), .A3(new_n817), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n970), .A2(new_n982), .ZN(new_n983));
  AND4_X1   g797(.A1(new_n221), .A2(new_n983), .A3(new_n823), .A4(new_n967), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n684), .A2(new_n221), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n977), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n979), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n984), .A2(new_n985), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n988), .A2(G953), .A3(new_n980), .A4(new_n977), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n987), .A2(new_n989), .ZN(G72));
  INV_X1    g804(.A(new_n853), .ZN(new_n991));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  XOR2_X1   g807(.A(new_n506), .B(KEYINPUT127), .Z(new_n994));
  OAI211_X1 g808(.A(new_n991), .B(new_n993), .C1(new_n699), .C2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n983), .A2(new_n962), .A3(new_n823), .A4(new_n967), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n996), .A2(new_n993), .ZN(new_n997));
  INV_X1    g811(.A(new_n505), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n484), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n950), .B(new_n995), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n969), .A2(new_n962), .A3(new_n970), .A4(new_n973), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n998), .B1(new_n1001), .B2(new_n993), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1000), .B1(new_n1002), .B2(new_n483), .ZN(G57));
endmodule


