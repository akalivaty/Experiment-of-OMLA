//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G952), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n188), .B1(G234), .B2(G237), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT72), .B(G902), .Z(new_n191));
  AOI211_X1 g005(.A(new_n187), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT21), .B(G898), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n190), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G214), .B1(G237), .B2(G902), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT67), .B1(new_n200), .B2(G116), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n198), .A3(G119), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n199), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT5), .ZN(new_n205));
  INV_X1    g019(.A(new_n199), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n205), .B(G113), .C1(KEYINPUT5), .C2(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT2), .A2(G113), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n210));
  INV_X1    g024(.A(G113), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n208), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n204), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(new_n216), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G104), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(G107), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n217), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n216), .A2(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n219), .A2(G104), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n207), .A2(new_n215), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n217), .A2(new_n220), .A3(new_n222), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n230), .A2(KEYINPUT79), .A3(G101), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT79), .B1(new_n230), .B2(G101), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n223), .A2(KEYINPUT4), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n230), .A2(G101), .A3(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n204), .A2(new_n214), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n204), .A2(new_n214), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n234), .A2(new_n239), .A3(KEYINPUT81), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n230), .A2(G101), .A3(new_n235), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n201), .A2(new_n203), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n206), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n212), .A2(new_n213), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT2), .A2(G113), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n242), .B1(new_n248), .B2(new_n215), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n230), .A2(G101), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT79), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n230), .A2(KEYINPUT79), .A3(G101), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n253), .A4(new_n223), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n241), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n229), .B1(new_n240), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G110), .B(G122), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT81), .B1(new_n234), .B2(new_n239), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n249), .A2(new_n254), .A3(new_n241), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n228), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n257), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(KEYINPUT6), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G146), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G143), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(G143), .B(G146), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT0), .B(G128), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n270), .B(G125), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(KEYINPUT1), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n275), .A2(new_n266), .A3(new_n268), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n266), .A2(new_n268), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(KEYINPUT65), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G128), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT1), .B1(new_n267), .B2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n276), .B1(new_n277), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n273), .B1(new_n284), .B2(G125), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n187), .A2(G224), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n287), .B(KEYINPUT82), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n256), .A2(new_n289), .A3(new_n258), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n264), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n286), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT85), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n285), .A2(new_n294), .A3(KEYINPUT7), .A4(new_n286), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n257), .B(KEYINPUT8), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n227), .A2(new_n215), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n205), .A2(KEYINPUT83), .ZN(new_n299));
  OAI21_X1  g113(.A(G113), .B1(new_n206), .B2(KEYINPUT5), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n205), .B2(KEYINPUT83), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n298), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n227), .B1(new_n207), .B2(new_n215), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n297), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT7), .ZN(new_n305));
  AOI22_X1  g119(.A1(KEYINPUT84), .A2(new_n305), .B1(new_n187), .B2(G224), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(KEYINPUT84), .B2(new_n305), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n273), .B(new_n307), .C1(new_n284), .C2(G125), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n296), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(G902), .B1(new_n309), .B2(new_n263), .ZN(new_n310));
  OAI21_X1  g124(.A(G210), .B1(G237), .B2(G902), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n291), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n311), .B1(new_n291), .B2(new_n310), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n196), .B(new_n197), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  OAI21_X1  g129(.A(G221), .B1(new_n315), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT11), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(G137), .ZN(new_n319));
  AND2_X1   g133(.A1(KEYINPUT64), .A2(G134), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT64), .A2(G134), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G137), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT11), .A3(G134), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(G137), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G131), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  OR2_X1    g141(.A1(KEYINPUT64), .A2(G134), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(KEYINPUT11), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT64), .A2(G134), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G131), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n324), .A4(new_n325), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n242), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n254), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT10), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n282), .A2(G128), .B1(new_n266), .B2(new_n268), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n223), .B(new_n226), .C1(new_n340), .C2(new_n276), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT65), .B(G128), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(G143), .B2(new_n265), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n277), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n271), .A2(new_n275), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n339), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n339), .A2(new_n341), .B1(new_n347), .B2(new_n227), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n335), .B1(new_n338), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n338), .A2(new_n335), .A3(new_n348), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n187), .A2(G227), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT78), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G140), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n345), .A2(new_n346), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n341), .B1(new_n357), .B2(new_n227), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n358), .A2(KEYINPUT12), .A3(new_n334), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT12), .B1(new_n358), .B2(new_n334), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n351), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n355), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n350), .A2(new_n356), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G469), .B1(new_n363), .B2(G902), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n338), .A2(new_n335), .A3(new_n348), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n362), .B1(new_n365), .B2(new_n349), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n351), .B(new_n355), .C1(new_n359), .C2(new_n360), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G469), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(new_n191), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n317), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G478), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(KEYINPUT15), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G217), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n315), .A2(new_n375), .A3(G953), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n267), .A2(G128), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT13), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT95), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n278), .A2(new_n280), .A3(G143), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n379), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT95), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n383), .A2(new_n267), .A3(KEYINPUT13), .A4(G128), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n380), .A2(new_n381), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G134), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n320), .A2(new_n321), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n381), .A2(KEYINPUT96), .A3(new_n387), .A4(new_n378), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n381), .A2(new_n387), .A3(new_n378), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT96), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n386), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n198), .A2(G122), .ZN(new_n393));
  INV_X1    g207(.A(G122), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G116), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT93), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n393), .B2(new_n395), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n219), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n393), .A2(new_n395), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT93), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(G107), .A3(new_n397), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT94), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n400), .A2(new_n403), .A3(KEYINPUT94), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n392), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n198), .A2(KEYINPUT14), .A3(G122), .ZN(new_n409));
  OAI211_X1 g223(.A(G107), .B(new_n409), .C1(new_n401), .C2(KEYINPUT14), .ZN(new_n410));
  INV_X1    g224(.A(new_n389), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n387), .B1(new_n381), .B2(new_n378), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n400), .B(new_n410), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n377), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n385), .A2(G134), .B1(new_n389), .B2(new_n390), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n400), .A2(new_n403), .A3(KEYINPUT94), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT94), .B1(new_n400), .B2(new_n403), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n388), .B(new_n416), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n413), .A3(new_n376), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n374), .B1(new_n421), .B2(new_n191), .ZN(new_n422));
  INV_X1    g236(.A(new_n191), .ZN(new_n423));
  AOI211_X1 g237(.A(new_n423), .B(new_n373), .C1(new_n415), .C2(new_n420), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(G237), .A2(G953), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G214), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n267), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(G143), .A3(G214), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n332), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n429), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G131), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT17), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n428), .A2(KEYINPUT87), .A3(new_n332), .A4(new_n429), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n432), .A2(new_n434), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT77), .ZN(new_n438));
  INV_X1    g252(.A(G125), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n439), .A2(KEYINPUT16), .A3(G140), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G140), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G125), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(G140), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT16), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n438), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n440), .A2(KEYINPUT77), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n265), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n447), .ZN(new_n449));
  XNOR2_X1  g263(.A(G125), .B(G140), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n440), .B1(new_n450), .B2(KEYINPUT16), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n449), .B(G146), .C1(new_n451), .C2(new_n438), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n433), .A2(KEYINPUT17), .A3(G131), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n437), .A2(new_n448), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(KEYINPUT18), .A2(G131), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n433), .B(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n443), .A2(new_n444), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT86), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT86), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n443), .A2(new_n444), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(G146), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n450), .A2(new_n265), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n454), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G113), .B(G122), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(new_n216), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n467), .B(KEYINPUT90), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n454), .A2(new_n464), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(G902), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT92), .B(G475), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT20), .ZN(new_n475));
  NOR2_X1   g289(.A1(G475), .A2(G902), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT19), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n443), .A2(new_n444), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT88), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n450), .A2(KEYINPUT88), .A3(new_n477), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n458), .A2(KEYINPUT19), .A3(new_n460), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n265), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n452), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT89), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n432), .A2(new_n436), .A3(new_n434), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(new_n489), .A3(new_n452), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n467), .B1(new_n491), .B2(new_n464), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n454), .A2(new_n464), .A3(new_n470), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n475), .B(new_n476), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT91), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n487), .B1(new_n485), .B2(KEYINPUT89), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n497), .A2(new_n490), .B1(new_n463), .B2(new_n456), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n471), .B1(new_n498), .B2(new_n467), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n499), .A2(KEYINPUT91), .A3(new_n475), .A4(new_n476), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n491), .A2(new_n464), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n493), .B1(new_n501), .B2(new_n468), .ZN(new_n502));
  INV_X1    g316(.A(new_n476), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT20), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n496), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n371), .A2(new_n425), .A3(new_n474), .A4(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n314), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n248), .A2(new_n215), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n332), .B1(G134), .B2(G137), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n328), .A2(new_n330), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(G137), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n333), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(new_n284), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n336), .B1(new_n327), .B2(new_n333), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT30), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n516));
  INV_X1    g330(.A(new_n336), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n322), .A2(G131), .A3(new_n326), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n324), .A2(new_n325), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n332), .B1(new_n519), .B2(new_n331), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n357), .A2(new_n333), .A3(new_n511), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n508), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n237), .A2(new_n238), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n426), .A2(G210), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT27), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT26), .B(G101), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT68), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT68), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n526), .A2(new_n533), .A3(new_n530), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n524), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT31), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT31), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n524), .A2(new_n532), .A3(new_n537), .A4(new_n534), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n513), .A2(new_n514), .A3(new_n508), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n525), .B1(new_n521), .B2(new_n522), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT28), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT28), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n526), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n530), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n536), .A2(new_n538), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(G472), .A2(G902), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT69), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT32), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n547), .A2(KEYINPUT69), .A3(new_n548), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n547), .A2(KEYINPUT32), .A3(new_n548), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n542), .B1(new_n556), .B2(new_n526), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n526), .A2(new_n542), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT29), .B1(new_n559), .B2(new_n530), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT70), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT30), .B1(new_n513), .B2(new_n514), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n521), .A2(new_n516), .A3(new_n522), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n539), .B1(new_n564), .B2(new_n508), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n561), .B1(new_n565), .B2(new_n530), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n525), .B1(new_n562), .B2(new_n563), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT70), .B(new_n545), .C1(new_n567), .C2(new_n539), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n560), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT71), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n559), .A2(new_n570), .A3(KEYINPUT29), .A4(new_n530), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n541), .A2(KEYINPUT29), .A3(new_n530), .A4(new_n543), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT71), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n574), .A3(new_n191), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT73), .B1(new_n575), .B2(G472), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT73), .ZN(new_n577));
  INV_X1    g391(.A(G472), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n423), .B1(new_n571), .B2(new_n573), .ZN(new_n579));
  AOI211_X1 g393(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n569), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n554), .B(new_n555), .C1(new_n576), .C2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n375), .B1(new_n191), .B2(G234), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n448), .A2(new_n452), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n278), .A2(new_n280), .A3(G119), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n200), .A2(G128), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT74), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n589), .A3(new_n586), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT24), .B(G110), .Z(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n342), .A2(KEYINPUT23), .A3(G119), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT75), .B1(new_n586), .B2(KEYINPUT23), .ZN(new_n594));
  OAI211_X1 g408(.A(KEYINPUT75), .B(KEYINPUT23), .C1(new_n274), .C2(G119), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n274), .A2(G119), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n593), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n598), .A2(KEYINPUT76), .A3(G110), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT76), .B1(new_n598), .B2(G110), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n584), .B(new_n592), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n591), .B1(new_n588), .B2(new_n590), .ZN(new_n602));
  INV_X1    g416(.A(G110), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n593), .B(new_n603), .C1(new_n594), .C2(new_n597), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n452), .B(new_n462), .C1(new_n602), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT22), .B(G137), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n609));
  XOR2_X1   g423(.A(new_n608), .B(new_n609), .Z(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n601), .A2(new_n606), .A3(new_n610), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n191), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT25), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n612), .A2(KEYINPUT25), .A3(new_n191), .A4(new_n613), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n583), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n612), .A2(new_n613), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n582), .A2(G902), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n507), .A2(new_n581), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  NAND2_X1  g439(.A1(new_n505), .A2(new_n474), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n421), .A2(new_n372), .A3(new_n191), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n408), .A2(new_n414), .A3(new_n377), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n376), .B1(new_n419), .B2(new_n413), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT33), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n415), .A2(new_n420), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n423), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n627), .B1(new_n633), .B2(new_n372), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT98), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n636), .B(new_n627), .C1(new_n633), .C2(new_n372), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n626), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n314), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n547), .A2(new_n191), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G472), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n551), .A2(new_n641), .A3(new_n553), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n623), .A2(new_n371), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT97), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n361), .A2(new_n362), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n350), .A2(new_n351), .A3(new_n355), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n646), .A3(G469), .ZN(new_n647));
  NAND2_X1  g461(.A1(G469), .A2(G902), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI211_X1 g463(.A(G469), .B(new_n423), .C1(new_n366), .C2(new_n367), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n316), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n651), .A2(new_n622), .A3(new_n618), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n547), .A2(KEYINPUT69), .A3(new_n548), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT69), .B1(new_n547), .B2(new_n548), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n652), .A2(new_n653), .A3(new_n656), .A4(new_n641), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n639), .A2(new_n644), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n504), .A2(new_n661), .A3(new_n494), .ZN(new_n662));
  INV_X1    g476(.A(new_n425), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n499), .A2(KEYINPUT99), .A3(new_n475), .A4(new_n476), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n662), .A2(new_n663), .A3(new_n474), .A4(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n314), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n644), .A3(new_n657), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  INV_X1    g483(.A(new_n642), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n616), .A2(new_n617), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n582), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n607), .A2(KEYINPUT100), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n611), .A2(KEYINPUT36), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n601), .A2(new_n675), .A3(new_n606), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n674), .B1(new_n673), .B2(new_n676), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n620), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n672), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n507), .A2(new_n670), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  OAI21_X1  g498(.A(new_n197), .B1(new_n312), .B2(new_n313), .ZN(new_n685));
  INV_X1    g499(.A(new_n680), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n371), .B1(new_n618), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n189), .B1(new_n192), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n472), .B2(new_n473), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n581), .A2(new_n688), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  NAND2_X1  g510(.A1(new_n556), .A2(new_n526), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n578), .B1(new_n697), .B2(new_n545), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n535), .A2(new_n698), .B1(G472), .B2(G902), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT102), .Z(new_n700));
  NAND3_X1  g514(.A1(new_n554), .A2(new_n555), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT103), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n554), .A2(new_n703), .A3(new_n700), .A4(new_n555), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n312), .A2(new_n313), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n691), .B(KEYINPUT39), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n371), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n711), .A2(new_n712), .A3(new_n681), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n197), .B1(new_n422), .B2(new_n424), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n505), .B2(new_n474), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n705), .A2(new_n708), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  AND4_X1   g531(.A1(new_n626), .A2(new_n635), .A3(new_n637), .A4(new_n692), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n581), .A2(new_n688), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  AOI21_X1  g534(.A(new_n369), .B1(new_n368), .B2(new_n191), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n721), .A2(new_n650), .A3(new_n317), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n639), .A2(new_n581), .A3(new_n623), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n623), .ZN(new_n726));
  INV_X1    g540(.A(new_n555), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n656), .B2(new_n552), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n575), .A2(G472), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n577), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n575), .A2(KEYINPUT73), .A3(G472), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n726), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(KEYINPUT104), .A3(new_n639), .A4(new_n722), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n725), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NAND4_X1  g551(.A1(new_n666), .A2(new_n581), .A3(new_n623), .A4(new_n722), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  AND3_X1   g553(.A1(new_n505), .A2(new_n425), .A3(new_n474), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n722), .B(new_n197), .C1(new_n312), .C2(new_n313), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n681), .A2(new_n196), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n581), .A2(new_n740), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT105), .B(G119), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G21));
  NAND2_X1  g560(.A1(new_n291), .A2(new_n310), .ZN(new_n747));
  INV_X1    g561(.A(new_n311), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n291), .A2(new_n310), .A3(new_n311), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(new_n715), .ZN(new_n752));
  AOI22_X1  g566(.A1(new_n535), .A2(KEYINPUT31), .B1(new_n544), .B2(new_n545), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n538), .B1(new_n753), .B2(KEYINPUT106), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n548), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n756), .A2(new_n623), .A3(new_n641), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n752), .A2(new_n757), .A3(new_n196), .A4(new_n722), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  AND3_X1   g573(.A1(new_n756), .A2(new_n641), .A3(new_n681), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n718), .A2(new_n742), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n749), .A2(new_n197), .A3(new_n750), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n651), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n733), .A2(new_n763), .A3(new_n718), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n576), .A2(new_n580), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT32), .B1(new_n547), .B2(new_n548), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(KEYINPUT107), .B2(new_n555), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n555), .A2(KEYINPUT107), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n623), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n765), .A2(new_n718), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT42), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n766), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT108), .B(G131), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G33));
  NAND3_X1  g591(.A1(new_n733), .A2(new_n694), .A3(new_n765), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n626), .B(KEYINPUT110), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n635), .A2(KEYINPUT43), .A3(new_n637), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n626), .B(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n782), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(KEYINPUT111), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT43), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n635), .A2(new_n637), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n505), .A2(new_n474), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n635), .A2(KEYINPUT109), .A3(new_n637), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n783), .A2(new_n787), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n681), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n795), .A2(new_n670), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(KEYINPUT44), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n798), .A2(KEYINPUT112), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(KEYINPUT112), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n363), .A2(KEYINPUT45), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n363), .A2(KEYINPUT45), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(G469), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n648), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT46), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n370), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n804), .A2(new_n805), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n316), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n709), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n764), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n797), .B2(KEYINPUT44), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n799), .A2(new_n800), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  XNOR2_X1  g630(.A(new_n809), .B(KEYINPUT47), .ZN(new_n817));
  INV_X1    g631(.A(new_n581), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(new_n726), .A3(new_n718), .A4(new_n812), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n794), .A2(new_n788), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n781), .A2(new_n780), .A3(new_n782), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT111), .B1(new_n785), .B2(new_n786), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n826), .A2(new_n189), .A3(new_n757), .ZN(new_n827));
  INV_X1    g641(.A(new_n722), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n708), .A2(new_n197), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(KEYINPUT50), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n826), .A2(new_n189), .A3(new_n757), .A4(new_n829), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT50), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n795), .A2(new_n190), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n764), .A2(new_n828), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n760), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n826), .A2(new_n189), .A3(new_n760), .A4(new_n837), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n705), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n764), .A2(new_n726), .A3(new_n828), .A4(new_n190), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n792), .A2(new_n842), .A3(new_n789), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n721), .A2(new_n650), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n317), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n764), .B1(new_n817), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n844), .B1(new_n847), .B2(new_n827), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n834), .A2(KEYINPUT51), .A3(new_n841), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT48), .ZN(new_n850));
  INV_X1    g664(.A(new_n772), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n835), .A2(new_n850), .A3(new_n851), .A4(new_n837), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n826), .A2(new_n189), .A3(new_n851), .A4(new_n837), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT48), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n188), .B(KEYINPUT118), .Z(new_n857));
  NAND2_X1  g671(.A1(new_n842), .A2(new_n843), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(new_n638), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n827), .B2(new_n742), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n855), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n856), .B1(new_n855), .B2(new_n860), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n849), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n834), .A2(KEYINPUT116), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n830), .A2(new_n833), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n865), .A2(new_n867), .A3(new_n841), .A4(new_n848), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n863), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n740), .B1(new_n626), .B2(new_n789), .ZN(new_n871));
  INV_X1    g685(.A(new_n314), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n644), .A3(new_n657), .A4(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n873), .A2(new_n682), .A3(new_n744), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n738), .A2(new_n624), .A3(new_n758), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n735), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n764), .A2(new_n687), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n693), .A2(new_n424), .A3(new_n422), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n664), .A3(new_n662), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT113), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT113), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n878), .A2(new_n662), .A3(new_n881), .A4(new_n664), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n877), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n718), .A2(new_n760), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n883), .A2(new_n581), .B1(new_n884), .B2(new_n765), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n774), .A3(new_n766), .A4(new_n778), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n876), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n651), .A2(new_n691), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n796), .A2(new_n751), .A3(new_n715), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n705), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n719), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n695), .A2(new_n761), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n888), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n719), .A2(KEYINPUT52), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n890), .B1(new_n702), .B2(new_n704), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT114), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n695), .A2(new_n761), .A3(KEYINPUT114), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n898), .A2(new_n900), .A3(KEYINPUT115), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n695), .A2(KEYINPUT114), .A3(new_n761), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT114), .B1(new_n695), .B2(new_n761), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT115), .B1(new_n906), .B2(new_n898), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n887), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n719), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n897), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n695), .A2(new_n761), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT52), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR4_X1   g728(.A1(new_n894), .A2(new_n897), .A3(new_n911), .A4(new_n888), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n887), .B(KEYINPUT53), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n870), .B1(new_n910), .B2(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n887), .B(KEYINPUT53), .C1(new_n903), .C2(new_n907), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n915), .A2(new_n914), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n873), .A2(new_n744), .A3(new_n682), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n738), .A2(new_n624), .A3(new_n758), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n884), .A2(new_n765), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n581), .A2(new_n877), .A3(new_n880), .A4(new_n882), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n778), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n922), .A2(new_n925), .A3(new_n775), .A4(new_n735), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n909), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n918), .A2(new_n927), .A3(new_n870), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n917), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(G952), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n869), .A2(new_n929), .B1(new_n930), .B2(new_n187), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n845), .B(KEYINPUT49), .Z(new_n932));
  NAND2_X1  g746(.A1(new_n316), .A2(new_n197), .ZN(new_n933));
  OR4_X1    g747(.A1(new_n726), .A2(new_n932), .A3(new_n789), .A4(new_n933), .ZN(new_n934));
  NOR4_X1   g748(.A1(new_n934), .A2(new_n705), .A3(new_n708), .A4(new_n781), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n822), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n868), .A2(new_n864), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n861), .A2(new_n862), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n929), .A2(new_n937), .A3(new_n938), .A4(new_n849), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n930), .A2(new_n187), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n935), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n941), .A2(KEYINPUT120), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n936), .A2(new_n943), .ZN(G75));
  NOR2_X1   g758(.A1(new_n187), .A2(G952), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n191), .B1(new_n918), .B2(new_n927), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT56), .B1(new_n947), .B2(new_n748), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n264), .A2(new_n290), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n288), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n946), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n947), .B(KEYINPUT121), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n748), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT56), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n952), .B1(new_n954), .B2(new_n956), .ZN(G51));
  INV_X1    g771(.A(new_n953), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n958), .A2(new_n803), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n918), .A2(new_n927), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT54), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n918), .A2(new_n927), .A3(new_n870), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n648), .B(KEYINPUT57), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n368), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n945), .B1(new_n959), .B2(new_n966), .ZN(G54));
  NAND2_X1  g781(.A1(KEYINPUT58), .A2(G475), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n958), .A2(new_n502), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n968), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n499), .B1(new_n953), .B2(new_n970), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n969), .A2(new_n971), .A3(new_n945), .ZN(G60));
  INV_X1    g786(.A(KEYINPUT122), .ZN(new_n973));
  NAND2_X1  g787(.A1(G478), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT59), .Z(new_n975));
  NAND3_X1  g789(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT115), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n902), .A3(new_n895), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT53), .B1(new_n979), .B2(new_n887), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n919), .A2(new_n926), .A3(new_n909), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT54), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n975), .B1(new_n982), .B2(new_n962), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n630), .A2(new_n632), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n973), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n975), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n917), .B2(new_n928), .ZN(new_n987));
  INV_X1    g801(.A(new_n984), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(KEYINPUT122), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n975), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n945), .B1(new_n963), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n985), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(KEYINPUT123), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT123), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n985), .A2(new_n989), .A3(new_n994), .A4(new_n991), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(G63));
  XOR2_X1   g810(.A(KEYINPUT124), .B(KEYINPUT60), .Z(new_n997));
  NAND2_X1  g811(.A1(G217), .A2(G902), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n960), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n945), .B1(new_n1000), .B2(new_n619), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n678), .A2(new_n679), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(new_n1000), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT61), .Z(G66));
  XNOR2_X1  g818(.A(new_n876), .B(KEYINPUT125), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n187), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT126), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n187), .B1(new_n195), .B2(G224), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n949), .B1(G898), .B2(new_n187), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1009), .B(new_n1010), .Z(G69));
  NOR2_X1   g825(.A1(new_n764), .A2(new_n710), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n733), .A2(new_n871), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n820), .A2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n904), .A2(new_n905), .A3(new_n911), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n716), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1014), .B1(new_n1016), .B2(KEYINPUT62), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n815), .B(new_n1017), .C1(KEYINPUT62), .C2(new_n1016), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n187), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n482), .A2(new_n483), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n564), .B(new_n1020), .Z(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(G900), .B2(G953), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n811), .A2(new_n851), .A3(new_n752), .ZN(new_n1025));
  AND4_X1   g839(.A1(new_n775), .A2(new_n820), .A3(new_n778), .A4(new_n1025), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n815), .A2(new_n1015), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1024), .B1(new_n1027), .B2(G953), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1030), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1023), .A2(new_n1032), .A3(new_n1028), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1031), .A2(new_n1033), .ZN(G72));
  NAND2_X1  g848(.A1(G472), .A2(G902), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT63), .Z(new_n1036));
  OAI21_X1  g850(.A(new_n1036), .B1(new_n1027), .B2(new_n1005), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1037), .A2(new_n545), .A3(new_n565), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n566), .A2(new_n568), .A3(new_n535), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(new_n1036), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1040), .B(KEYINPUT127), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1041), .B1(new_n980), .B2(new_n981), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1038), .A2(new_n946), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1036), .B1(new_n1018), .B2(new_n1005), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n565), .A2(new_n545), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(G57));
endmodule


