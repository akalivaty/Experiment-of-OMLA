

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(n565), .A2(G2104), .ZN(n895) );
  XNOR2_X1 U554 ( .A(n553), .B(KEYINPUT65), .ZN(n552) );
  AND2_X1 U555 ( .A1(n803), .A2(n804), .ZN(n753) );
  XNOR2_X1 U556 ( .A(KEYINPUT103), .B(KEYINPUT31), .ZN(n738) );
  INV_X1 U557 ( .A(n798), .ZN(n541) );
  NOR2_X1 U558 ( .A1(n539), .A2(KEYINPUT106), .ZN(n538) );
  INV_X1 U559 ( .A(n986), .ZN(n539) );
  INV_X1 U560 ( .A(G2105), .ZN(n565) );
  AND2_X1 U561 ( .A1(n753), .A2(G1996), .ZN(n741) );
  AND2_X1 U562 ( .A1(n551), .A2(n516), .ZN(n751) );
  AND2_X1 U563 ( .A1(n760), .A2(n535), .ZN(n534) );
  NAND2_X1 U564 ( .A1(n532), .A2(KEYINPUT29), .ZN(n531) );
  NAND2_X1 U565 ( .A1(n526), .A2(n524), .ZN(n523) );
  AND2_X1 U566 ( .A1(n525), .A2(n763), .ZN(n524) );
  NAND2_X1 U567 ( .A1(n530), .A2(KEYINPUT100), .ZN(n528) );
  AND2_X1 U568 ( .A1(n773), .A2(n767), .ZN(n768) );
  AND2_X1 U569 ( .A1(n781), .A2(n780), .ZN(n783) );
  NOR2_X1 U570 ( .A1(n540), .A2(n536), .ZN(n787) );
  NAND2_X1 U571 ( .A1(G8), .A2(n774), .ZN(n798) );
  XNOR2_X1 U572 ( .A(KEYINPUT91), .B(n727), .ZN(n803) );
  NOR2_X1 U573 ( .A1(n675), .A2(n582), .ZN(n558) );
  NAND2_X1 U574 ( .A1(n557), .A2(n555), .ZN(n554) );
  OR2_X1 U575 ( .A1(n802), .A2(n801), .ZN(n557) );
  INV_X1 U576 ( .A(n844), .ZN(n556) );
  XNOR2_X1 U577 ( .A(n633), .B(KEYINPUT15), .ZN(n987) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n583), .Z(n688) );
  XNOR2_X1 U579 ( .A(n579), .B(KEYINPUT66), .ZN(n689) );
  XNOR2_X1 U580 ( .A(n566), .B(n549), .ZN(n548) );
  XNOR2_X1 U581 ( .A(KEYINPUT67), .B(KEYINPUT23), .ZN(n549) );
  NOR2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n568) );
  AND2_X1 U583 ( .A1(n573), .A2(G113), .ZN(n550) );
  AND2_X1 U584 ( .A1(n545), .A2(n544), .ZN(G160) );
  AND2_X1 U585 ( .A1(n547), .A2(n546), .ZN(n545) );
  NAND2_X1 U586 ( .A1(n651), .A2(G137), .ZN(n544) );
  AND2_X1 U587 ( .A1(n548), .A2(n570), .ZN(n546) );
  OR2_X1 U588 ( .A1(G301), .A2(n762), .ZN(n515) );
  OR2_X1 U589 ( .A1(n749), .A2(n748), .ZN(n516) );
  AND2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n517) );
  NAND2_X1 U591 ( .A1(n748), .A2(n749), .ZN(n518) );
  AND2_X1 U592 ( .A1(n531), .A2(n515), .ZN(n519) );
  XNOR2_X2 U593 ( .A(n569), .B(KEYINPUT17), .ZN(n651) );
  OR2_X1 U594 ( .A1(n986), .A2(n542), .ZN(n520) );
  AND2_X1 U595 ( .A1(n541), .A2(n520), .ZN(n521) );
  INV_X1 U596 ( .A(KEYINPUT106), .ZN(n542) );
  AND2_X1 U597 ( .A1(KEYINPUT100), .A2(KEYINPUT29), .ZN(n522) );
  NAND2_X1 U598 ( .A1(n517), .A2(n523), .ZN(n764) );
  NAND2_X1 U599 ( .A1(n529), .A2(KEYINPUT29), .ZN(n525) );
  INV_X1 U600 ( .A(n530), .ZN(n526) );
  NAND2_X1 U601 ( .A1(n529), .A2(n522), .ZN(n527) );
  INV_X1 U602 ( .A(n761), .ZN(n529) );
  NAND2_X1 U603 ( .A1(n533), .A2(n519), .ZN(n530) );
  INV_X1 U604 ( .A(n760), .ZN(n532) );
  NAND2_X1 U605 ( .A1(n761), .A2(n534), .ZN(n533) );
  INV_X1 U606 ( .A(KEYINPUT29), .ZN(n535) );
  NAND2_X1 U607 ( .A1(n537), .A2(n521), .ZN(n536) );
  NAND2_X1 U608 ( .A1(n543), .A2(n538), .ZN(n537) );
  NOR2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n540) );
  NAND2_X1 U610 ( .A1(n792), .A2(n988), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n550), .B(KEYINPUT69), .ZN(n547) );
  NAND2_X1 U612 ( .A1(n552), .A2(n518), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n745), .A2(n744), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n850), .ZN(n852) );
  NOR2_X1 U615 ( .A1(n827), .A2(n556), .ZN(n555) );
  XOR2_X1 U616 ( .A(KEYINPUT76), .B(n629), .Z(n559) );
  AND2_X1 U617 ( .A1(n696), .A2(G43), .ZN(n560) );
  XNOR2_X1 U618 ( .A(KEYINPUT14), .B(n617), .ZN(n561) );
  OR2_X1 U619 ( .A1(n789), .A2(n798), .ZN(n562) );
  XOR2_X1 U620 ( .A(KEYINPUT101), .B(n728), .Z(n563) );
  INV_X1 U621 ( .A(KEYINPUT99), .ZN(n750) );
  INV_X1 U622 ( .A(KEYINPUT100), .ZN(n763) );
  XNOR2_X1 U623 ( .A(n739), .B(n738), .ZN(n765) );
  NAND2_X1 U624 ( .A1(n804), .A2(n803), .ZN(n774) );
  NAND2_X1 U625 ( .A1(G40), .A2(G160), .ZN(n727) );
  NAND2_X1 U626 ( .A1(n562), .A2(n1000), .ZN(n790) );
  NOR2_X1 U627 ( .A1(G164), .A2(G1384), .ZN(n804) );
  INV_X1 U628 ( .A(KEYINPUT0), .ZN(n578) );
  INV_X1 U629 ( .A(G2104), .ZN(n567) );
  XNOR2_X1 U630 ( .A(n578), .B(G543), .ZN(n675) );
  AND2_X1 U631 ( .A1(n567), .A2(G2105), .ZN(n898) );
  NOR2_X1 U632 ( .A1(n675), .A2(G651), .ZN(n696) );
  NAND2_X1 U633 ( .A1(n618), .A2(n561), .ZN(n994) );
  NAND2_X1 U634 ( .A1(G2104), .A2(G2105), .ZN(n564) );
  XOR2_X1 U635 ( .A(KEYINPUT68), .B(n564), .Z(n573) );
  NAND2_X1 U636 ( .A1(G101), .A2(n895), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n898), .A2(G125), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT70), .B(n568), .Z(n569) );
  NAND2_X1 U639 ( .A1(n895), .A2(G102), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G138), .A2(n651), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G126), .A2(n898), .ZN(n575) );
  BUF_X1 U643 ( .A(n573), .Z(n899) );
  NAND2_X1 U644 ( .A1(G114), .A2(n899), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U646 ( .A1(n577), .A2(n576), .ZN(G164) );
  INV_X1 U647 ( .A(G651), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n558), .A2(G72), .ZN(n581) );
  NOR2_X1 U649 ( .A1(G651), .A2(G543), .ZN(n579) );
  NAND2_X1 U650 ( .A1(G85), .A2(n689), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n587) );
  NOR2_X1 U652 ( .A1(G543), .A2(n582), .ZN(n583) );
  NAND2_X1 U653 ( .A1(G60), .A2(n688), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G47), .A2(n696), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  OR2_X1 U656 ( .A1(n587), .A2(n586), .ZN(G290) );
  XOR2_X1 U657 ( .A(G2438), .B(G2454), .Z(n589) );
  XNOR2_X1 U658 ( .A(G2435), .B(G2430), .ZN(n588) );
  XNOR2_X1 U659 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U660 ( .A(n590), .B(G2427), .Z(n592) );
  XNOR2_X1 U661 ( .A(G1348), .B(G1341), .ZN(n591) );
  XNOR2_X1 U662 ( .A(n592), .B(n591), .ZN(n596) );
  XOR2_X1 U663 ( .A(G2443), .B(G2446), .Z(n594) );
  XNOR2_X1 U664 ( .A(KEYINPUT108), .B(G2451), .ZN(n593) );
  XNOR2_X1 U665 ( .A(n594), .B(n593), .ZN(n595) );
  XOR2_X1 U666 ( .A(n596), .B(n595), .Z(n597) );
  AND2_X1 U667 ( .A1(G14), .A2(n597), .ZN(G401) );
  AND2_X1 U668 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U669 ( .A(G57), .ZN(G237) );
  INV_X1 U670 ( .A(G132), .ZN(G219) );
  NAND2_X1 U671 ( .A1(G63), .A2(n688), .ZN(n599) );
  NAND2_X1 U672 ( .A1(G51), .A2(n696), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U674 ( .A(KEYINPUT6), .B(n600), .ZN(n607) );
  NAND2_X1 U675 ( .A1(G89), .A2(n689), .ZN(n601) );
  XNOR2_X1 U676 ( .A(n601), .B(KEYINPUT4), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G76), .A2(n558), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U679 ( .A(KEYINPUT78), .B(n604), .Z(n605) );
  XNOR2_X1 U680 ( .A(KEYINPUT5), .B(n605), .ZN(n606) );
  NOR2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U682 ( .A(KEYINPUT7), .B(n608), .Z(G168) );
  XOR2_X1 U683 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U684 ( .A1(G7), .A2(G661), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U686 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n611) );
  INV_X1 U687 ( .A(G223), .ZN(n853) );
  NAND2_X1 U688 ( .A1(G567), .A2(n853), .ZN(n610) );
  XNOR2_X1 U689 ( .A(n611), .B(n610), .ZN(G234) );
  NAND2_X1 U690 ( .A1(G81), .A2(n689), .ZN(n612) );
  XNOR2_X1 U691 ( .A(n612), .B(KEYINPUT12), .ZN(n614) );
  NAND2_X1 U692 ( .A1(G68), .A2(n558), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U694 ( .A(KEYINPUT13), .B(n615), .Z(n616) );
  NOR2_X1 U695 ( .A1(n616), .A2(n560), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G56), .A2(n688), .ZN(n617) );
  INV_X1 U697 ( .A(G860), .ZN(n665) );
  OR2_X1 U698 ( .A1(n994), .A2(n665), .ZN(G153) );
  NAND2_X1 U699 ( .A1(n558), .A2(G77), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G90), .A2(n689), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U702 ( .A(KEYINPUT9), .B(n621), .ZN(n625) );
  NAND2_X1 U703 ( .A1(G64), .A2(n688), .ZN(n623) );
  NAND2_X1 U704 ( .A1(G52), .A2(n696), .ZN(n622) );
  AND2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(G301) );
  INV_X1 U707 ( .A(G301), .ZN(G171) );
  INV_X1 U708 ( .A(G868), .ZN(n708) );
  NOR2_X1 U709 ( .A1(n708), .A2(G171), .ZN(n626) );
  XNOR2_X1 U710 ( .A(n626), .B(KEYINPUT75), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G54), .A2(n696), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G66), .A2(n688), .ZN(n628) );
  NAND2_X1 U713 ( .A1(G79), .A2(n558), .ZN(n627) );
  NAND2_X1 U714 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n689), .A2(G92), .ZN(n629) );
  NOR2_X1 U716 ( .A1(n630), .A2(n559), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(n633) );
  INV_X1 U718 ( .A(n987), .ZN(n748) );
  NAND2_X1 U719 ( .A1(n708), .A2(n748), .ZN(n634) );
  NAND2_X1 U720 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U721 ( .A(KEYINPUT77), .B(n636), .Z(G284) );
  NAND2_X1 U722 ( .A1(G65), .A2(n688), .ZN(n638) );
  NAND2_X1 U723 ( .A1(G53), .A2(n696), .ZN(n637) );
  NAND2_X1 U724 ( .A1(n638), .A2(n637), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n558), .A2(G78), .ZN(n640) );
  NAND2_X1 U726 ( .A1(G91), .A2(n689), .ZN(n639) );
  NAND2_X1 U727 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U728 ( .A(KEYINPUT71), .B(n641), .Z(n642) );
  NOR2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n997) );
  XOR2_X1 U730 ( .A(n997), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U731 ( .A1(G299), .A2(G868), .ZN(n645) );
  NOR2_X1 U732 ( .A1(G286), .A2(n708), .ZN(n644) );
  NOR2_X1 U733 ( .A1(n645), .A2(n644), .ZN(G297) );
  NAND2_X1 U734 ( .A1(n665), .A2(G559), .ZN(n646) );
  NAND2_X1 U735 ( .A1(n646), .A2(n987), .ZN(n647) );
  XNOR2_X1 U736 ( .A(n647), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U737 ( .A1(G868), .A2(n994), .ZN(n650) );
  NAND2_X1 U738 ( .A1(G868), .A2(n987), .ZN(n648) );
  NOR2_X1 U739 ( .A1(G559), .A2(n648), .ZN(n649) );
  NOR2_X1 U740 ( .A1(n650), .A2(n649), .ZN(G282) );
  NAND2_X1 U741 ( .A1(n651), .A2(G135), .ZN(n652) );
  XNOR2_X1 U742 ( .A(n652), .B(KEYINPUT80), .ZN(n656) );
  XOR2_X1 U743 ( .A(KEYINPUT18), .B(KEYINPUT79), .Z(n654) );
  NAND2_X1 U744 ( .A1(G123), .A2(n898), .ZN(n653) );
  XNOR2_X1 U745 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U746 ( .A1(n656), .A2(n655), .ZN(n661) );
  NAND2_X1 U747 ( .A1(G99), .A2(n895), .ZN(n658) );
  NAND2_X1 U748 ( .A1(G111), .A2(n899), .ZN(n657) );
  NAND2_X1 U749 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U750 ( .A(KEYINPUT81), .B(n659), .Z(n660) );
  NOR2_X1 U751 ( .A1(n661), .A2(n660), .ZN(n936) );
  XNOR2_X1 U752 ( .A(n936), .B(G2096), .ZN(n663) );
  INV_X1 U753 ( .A(G2100), .ZN(n662) );
  NAND2_X1 U754 ( .A1(n663), .A2(n662), .ZN(G156) );
  NAND2_X1 U755 ( .A1(G559), .A2(n987), .ZN(n664) );
  XOR2_X1 U756 ( .A(n994), .B(n664), .Z(n706) );
  NAND2_X1 U757 ( .A1(n665), .A2(n706), .ZN(n674) );
  NAND2_X1 U758 ( .A1(n689), .A2(G93), .ZN(n666) );
  XNOR2_X1 U759 ( .A(n666), .B(KEYINPUT82), .ZN(n673) );
  NAND2_X1 U760 ( .A1(G67), .A2(n688), .ZN(n668) );
  NAND2_X1 U761 ( .A1(G55), .A2(n696), .ZN(n667) );
  NAND2_X1 U762 ( .A1(n668), .A2(n667), .ZN(n671) );
  NAND2_X1 U763 ( .A1(G80), .A2(n558), .ZN(n669) );
  XNOR2_X1 U764 ( .A(KEYINPUT83), .B(n669), .ZN(n670) );
  NOR2_X1 U765 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U766 ( .A1(n673), .A2(n672), .ZN(n709) );
  XNOR2_X1 U767 ( .A(n674), .B(n709), .ZN(G145) );
  NAND2_X1 U768 ( .A1(G87), .A2(n675), .ZN(n676) );
  XNOR2_X1 U769 ( .A(n676), .B(KEYINPUT84), .ZN(n681) );
  NAND2_X1 U770 ( .A1(G49), .A2(n696), .ZN(n678) );
  NAND2_X1 U771 ( .A1(G74), .A2(G651), .ZN(n677) );
  NAND2_X1 U772 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U773 ( .A1(n688), .A2(n679), .ZN(n680) );
  NAND2_X1 U774 ( .A1(n681), .A2(n680), .ZN(G288) );
  NAND2_X1 U775 ( .A1(n558), .A2(G75), .ZN(n683) );
  NAND2_X1 U776 ( .A1(G88), .A2(n689), .ZN(n682) );
  NAND2_X1 U777 ( .A1(n683), .A2(n682), .ZN(n687) );
  NAND2_X1 U778 ( .A1(G62), .A2(n688), .ZN(n685) );
  NAND2_X1 U779 ( .A1(G50), .A2(n696), .ZN(n684) );
  NAND2_X1 U780 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U781 ( .A1(n687), .A2(n686), .ZN(G166) );
  NAND2_X1 U782 ( .A1(G61), .A2(n688), .ZN(n691) );
  NAND2_X1 U783 ( .A1(G86), .A2(n689), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U785 ( .A1(G73), .A2(n558), .ZN(n692) );
  XNOR2_X1 U786 ( .A(n692), .B(KEYINPUT2), .ZN(n693) );
  XNOR2_X1 U787 ( .A(n693), .B(KEYINPUT85), .ZN(n694) );
  NOR2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n696), .A2(G48), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(G305) );
  XNOR2_X1 U791 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n700) );
  XNOR2_X1 U792 ( .A(G288), .B(KEYINPUT19), .ZN(n699) );
  XNOR2_X1 U793 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U794 ( .A(G299), .B(n701), .ZN(n703) );
  XNOR2_X1 U795 ( .A(G290), .B(G166), .ZN(n702) );
  XNOR2_X1 U796 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U797 ( .A(n704), .B(G305), .ZN(n705) );
  XNOR2_X1 U798 ( .A(n705), .B(n709), .ZN(n921) );
  XNOR2_X1 U799 ( .A(n706), .B(n921), .ZN(n707) );
  NOR2_X1 U800 ( .A1(n708), .A2(n707), .ZN(n711) );
  NOR2_X1 U801 ( .A1(G868), .A2(n709), .ZN(n710) );
  NOR2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U803 ( .A(KEYINPUT88), .B(n712), .ZN(G295) );
  NAND2_X1 U804 ( .A1(G2084), .A2(G2078), .ZN(n713) );
  XNOR2_X1 U805 ( .A(n713), .B(KEYINPUT89), .ZN(n714) );
  XNOR2_X1 U806 ( .A(n714), .B(KEYINPUT20), .ZN(n715) );
  NAND2_X1 U807 ( .A1(n715), .A2(G2090), .ZN(n716) );
  XNOR2_X1 U808 ( .A(KEYINPUT21), .B(n716), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n717), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U810 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U811 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  NOR2_X1 U812 ( .A1(G219), .A2(G220), .ZN(n718) );
  XOR2_X1 U813 ( .A(KEYINPUT22), .B(n718), .Z(n719) );
  NOR2_X1 U814 ( .A1(G218), .A2(n719), .ZN(n720) );
  XNOR2_X1 U815 ( .A(KEYINPUT90), .B(n720), .ZN(n721) );
  NAND2_X1 U816 ( .A1(n721), .A2(G96), .ZN(n932) );
  NAND2_X1 U817 ( .A1(G2106), .A2(n932), .ZN(n725) );
  NAND2_X1 U818 ( .A1(G69), .A2(G120), .ZN(n722) );
  NOR2_X1 U819 ( .A1(G237), .A2(n722), .ZN(n723) );
  NAND2_X1 U820 ( .A1(G108), .A2(n723), .ZN(n933) );
  NAND2_X1 U821 ( .A1(G567), .A2(n933), .ZN(n724) );
  NAND2_X1 U822 ( .A1(n725), .A2(n724), .ZN(n859) );
  NAND2_X1 U823 ( .A1(G483), .A2(G661), .ZN(n726) );
  NOR2_X1 U824 ( .A1(n859), .A2(n726), .ZN(n858) );
  NAND2_X1 U825 ( .A1(n858), .A2(G36), .ZN(G176) );
  INV_X1 U826 ( .A(G166), .ZN(G303) );
  NOR2_X1 U827 ( .A1(G2084), .A2(n774), .ZN(n769) );
  NOR2_X1 U828 ( .A1(G1966), .A2(n798), .ZN(n766) );
  NOR2_X1 U829 ( .A1(n769), .A2(n766), .ZN(n728) );
  NAND2_X1 U830 ( .A1(G8), .A2(n563), .ZN(n729) );
  XNOR2_X1 U831 ( .A(KEYINPUT30), .B(n729), .ZN(n730) );
  NOR2_X1 U832 ( .A1(G168), .A2(n730), .ZN(n737) );
  XNOR2_X1 U833 ( .A(G2078), .B(KEYINPUT25), .ZN(n731) );
  XNOR2_X1 U834 ( .A(n731), .B(KEYINPUT97), .ZN(n965) );
  NOR2_X1 U835 ( .A1(n965), .A2(n774), .ZN(n732) );
  XNOR2_X1 U836 ( .A(n732), .B(KEYINPUT98), .ZN(n734) );
  NOR2_X1 U837 ( .A1(n753), .A2(G1961), .ZN(n733) );
  NOR2_X1 U838 ( .A1(n734), .A2(n733), .ZN(n762) );
  NAND2_X1 U839 ( .A1(n762), .A2(G301), .ZN(n735) );
  XOR2_X1 U840 ( .A(KEYINPUT102), .B(n735), .Z(n736) );
  NOR2_X1 U841 ( .A1(n737), .A2(n736), .ZN(n739) );
  XOR2_X1 U842 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n740) );
  XNOR2_X1 U843 ( .A(n741), .B(n740), .ZN(n745) );
  NAND2_X1 U844 ( .A1(n774), .A2(G1341), .ZN(n743) );
  INV_X1 U845 ( .A(n994), .ZN(n742) );
  AND2_X1 U846 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U847 ( .A1(G1348), .A2(n774), .ZN(n747) );
  NAND2_X1 U848 ( .A1(n753), .A2(G2067), .ZN(n746) );
  NAND2_X1 U849 ( .A1(n747), .A2(n746), .ZN(n749) );
  XNOR2_X1 U850 ( .A(n751), .B(n750), .ZN(n757) );
  NAND2_X1 U851 ( .A1(n753), .A2(G2072), .ZN(n752) );
  XNOR2_X1 U852 ( .A(n752), .B(KEYINPUT27), .ZN(n755) );
  INV_X1 U853 ( .A(G1956), .ZN(n1016) );
  NOR2_X1 U854 ( .A1(n1016), .A2(n753), .ZN(n754) );
  NOR2_X1 U855 ( .A1(n755), .A2(n754), .ZN(n758) );
  NAND2_X1 U856 ( .A1(n758), .A2(n997), .ZN(n756) );
  NAND2_X1 U857 ( .A1(n757), .A2(n756), .ZN(n761) );
  NOR2_X1 U858 ( .A1(n758), .A2(n997), .ZN(n759) );
  XOR2_X1 U859 ( .A(n759), .B(KEYINPUT28), .Z(n760) );
  NAND2_X1 U860 ( .A1(n765), .A2(n764), .ZN(n773) );
  INV_X1 U861 ( .A(n766), .ZN(n767) );
  XNOR2_X1 U862 ( .A(n768), .B(KEYINPUT104), .ZN(n771) );
  NAND2_X1 U863 ( .A1(n769), .A2(G8), .ZN(n770) );
  NAND2_X1 U864 ( .A1(n771), .A2(n770), .ZN(n785) );
  AND2_X1 U865 ( .A1(G286), .A2(G8), .ZN(n772) );
  NAND2_X1 U866 ( .A1(n773), .A2(n772), .ZN(n781) );
  INV_X1 U867 ( .A(G8), .ZN(n779) );
  NOR2_X1 U868 ( .A1(G1971), .A2(n798), .ZN(n776) );
  NOR2_X1 U869 ( .A1(G2090), .A2(n774), .ZN(n775) );
  NOR2_X1 U870 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U871 ( .A1(n777), .A2(G303), .ZN(n778) );
  OR2_X1 U872 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U873 ( .A(KEYINPUT105), .B(KEYINPUT32), .Z(n782) );
  XNOR2_X1 U874 ( .A(n783), .B(n782), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n792) );
  NOR2_X1 U876 ( .A1(G1976), .A2(G288), .ZN(n788) );
  NOR2_X1 U877 ( .A1(G1971), .A2(G303), .ZN(n786) );
  NOR2_X1 U878 ( .A1(n788), .A2(n786), .ZN(n988) );
  NAND2_X1 U879 ( .A1(G1976), .A2(G288), .ZN(n986) );
  NOR2_X1 U880 ( .A1(KEYINPUT33), .A2(n787), .ZN(n791) );
  NAND2_X1 U881 ( .A1(n788), .A2(KEYINPUT33), .ZN(n789) );
  XOR2_X1 U882 ( .A(G1981), .B(G305), .Z(n1000) );
  NOR2_X1 U883 ( .A1(n791), .A2(n790), .ZN(n802) );
  NOR2_X1 U884 ( .A1(G2090), .A2(G303), .ZN(n793) );
  NAND2_X1 U885 ( .A1(G8), .A2(n793), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n792), .A2(n794), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n795), .A2(n798), .ZN(n800) );
  NOR2_X1 U888 ( .A1(G1981), .A2(G305), .ZN(n796) );
  XOR2_X1 U889 ( .A(n796), .B(KEYINPUT24), .Z(n797) );
  OR2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n801) );
  INV_X1 U892 ( .A(n803), .ZN(n805) );
  NOR2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U894 ( .A(n806), .B(KEYINPUT92), .ZN(n848) );
  INV_X1 U895 ( .A(n848), .ZN(n823) );
  NAND2_X1 U896 ( .A1(n651), .A2(G141), .ZN(n807) );
  XNOR2_X1 U897 ( .A(n807), .B(KEYINPUT96), .ZN(n814) );
  NAND2_X1 U898 ( .A1(G129), .A2(n898), .ZN(n809) );
  NAND2_X1 U899 ( .A1(G117), .A2(n899), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n895), .A2(G105), .ZN(n810) );
  XOR2_X1 U902 ( .A(KEYINPUT38), .B(n810), .Z(n811) );
  NOR2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n910) );
  AND2_X1 U905 ( .A1(n910), .A2(G1996), .ZN(n822) );
  NAND2_X1 U906 ( .A1(n895), .A2(G95), .ZN(n816) );
  NAND2_X1 U907 ( .A1(G131), .A2(n651), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n820) );
  NAND2_X1 U909 ( .A1(G119), .A2(n898), .ZN(n818) );
  NAND2_X1 U910 ( .A1(G107), .A2(n899), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n911) );
  INV_X1 U913 ( .A(G1991), .ZN(n963) );
  NOR2_X1 U914 ( .A1(n911), .A2(n963), .ZN(n821) );
  NOR2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n942) );
  NOR2_X1 U916 ( .A1(n823), .A2(n942), .ZN(n841) );
  INV_X1 U917 ( .A(n841), .ZN(n826) );
  XOR2_X1 U918 ( .A(G1986), .B(G290), .Z(n993) );
  NOR2_X1 U919 ( .A1(n823), .A2(n993), .ZN(n824) );
  XNOR2_X1 U920 ( .A(n824), .B(KEYINPUT93), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n895), .A2(G104), .ZN(n829) );
  NAND2_X1 U923 ( .A1(G140), .A2(n651), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U925 ( .A(KEYINPUT34), .B(n830), .ZN(n836) );
  NAND2_X1 U926 ( .A1(G128), .A2(n898), .ZN(n832) );
  NAND2_X1 U927 ( .A1(G116), .A2(n899), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n832), .A2(n831), .ZN(n833) );
  XOR2_X1 U929 ( .A(KEYINPUT35), .B(n833), .Z(n834) );
  XNOR2_X1 U930 ( .A(KEYINPUT94), .B(n834), .ZN(n835) );
  NOR2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  XOR2_X1 U932 ( .A(n837), .B(KEYINPUT36), .Z(n838) );
  XNOR2_X1 U933 ( .A(KEYINPUT95), .B(n838), .ZN(n918) );
  XNOR2_X1 U934 ( .A(G2067), .B(KEYINPUT37), .ZN(n846) );
  NOR2_X1 U935 ( .A1(n918), .A2(n846), .ZN(n937) );
  NAND2_X1 U936 ( .A1(n937), .A2(n848), .ZN(n844) );
  NOR2_X1 U937 ( .A1(G1996), .A2(n910), .ZN(n951) );
  NOR2_X1 U938 ( .A1(G1986), .A2(G290), .ZN(n839) );
  AND2_X1 U939 ( .A1(n963), .A2(n911), .ZN(n935) );
  NOR2_X1 U940 ( .A1(n839), .A2(n935), .ZN(n840) );
  NOR2_X1 U941 ( .A1(n841), .A2(n840), .ZN(n842) );
  NOR2_X1 U942 ( .A1(n951), .A2(n842), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n843), .B(KEYINPUT39), .ZN(n845) );
  NAND2_X1 U944 ( .A1(n845), .A2(n844), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n918), .A2(n846), .ZN(n941) );
  NAND2_X1 U946 ( .A1(n847), .A2(n941), .ZN(n849) );
  NAND2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n850) );
  XOR2_X1 U948 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(G329) );
  NAND2_X1 U950 ( .A1(G2106), .A2(n853), .ZN(G217) );
  NAND2_X1 U951 ( .A1(G15), .A2(G2), .ZN(n855) );
  INV_X1 U952 ( .A(G661), .ZN(n854) );
  NOR2_X1 U953 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n856), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U955 ( .A1(G3), .A2(G1), .ZN(n857) );
  NAND2_X1 U956 ( .A1(n858), .A2(n857), .ZN(G188) );
  XOR2_X1 U957 ( .A(G96), .B(KEYINPUT110), .Z(G221) );
  XNOR2_X1 U958 ( .A(KEYINPUT111), .B(n859), .ZN(G319) );
  XOR2_X1 U959 ( .A(G2100), .B(G2096), .Z(n861) );
  XNOR2_X1 U960 ( .A(KEYINPUT42), .B(G2678), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U962 ( .A(KEYINPUT43), .B(G2090), .Z(n863) );
  XNOR2_X1 U963 ( .A(G2067), .B(G2072), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U965 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U966 ( .A(G2084), .B(G2078), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(G227) );
  XNOR2_X1 U968 ( .A(G1961), .B(KEYINPUT112), .ZN(n877) );
  XOR2_X1 U969 ( .A(G1976), .B(G1971), .Z(n869) );
  XNOR2_X1 U970 ( .A(G1986), .B(G1956), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U972 ( .A(G1981), .B(G1966), .Z(n871) );
  XNOR2_X1 U973 ( .A(G1991), .B(G1996), .ZN(n870) );
  XNOR2_X1 U974 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U975 ( .A(n873), .B(n872), .Z(n875) );
  XNOR2_X1 U976 ( .A(G2474), .B(KEYINPUT41), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(G229) );
  NAND2_X1 U979 ( .A1(G100), .A2(n895), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G112), .A2(n899), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U982 ( .A(KEYINPUT114), .B(n880), .ZN(n886) );
  NAND2_X1 U983 ( .A1(G124), .A2(n898), .ZN(n881) );
  XOR2_X1 U984 ( .A(KEYINPUT113), .B(n881), .Z(n882) );
  XNOR2_X1 U985 ( .A(n882), .B(KEYINPUT44), .ZN(n884) );
  NAND2_X1 U986 ( .A1(G136), .A2(n651), .ZN(n883) );
  NAND2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U988 ( .A1(n886), .A2(n885), .ZN(G162) );
  NAND2_X1 U989 ( .A1(G130), .A2(n898), .ZN(n888) );
  NAND2_X1 U990 ( .A1(G118), .A2(n899), .ZN(n887) );
  NAND2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n895), .A2(G106), .ZN(n890) );
  NAND2_X1 U993 ( .A1(G142), .A2(n651), .ZN(n889) );
  NAND2_X1 U994 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U995 ( .A(KEYINPUT45), .B(n891), .Z(n892) );
  NOR2_X1 U996 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U997 ( .A(n894), .B(n936), .Z(n906) );
  NAND2_X1 U998 ( .A1(n895), .A2(G103), .ZN(n897) );
  NAND2_X1 U999 ( .A1(G139), .A2(n651), .ZN(n896) );
  NAND2_X1 U1000 ( .A1(n897), .A2(n896), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(G127), .A2(n898), .ZN(n901) );
  NAND2_X1 U1002 ( .A1(G115), .A2(n899), .ZN(n900) );
  NAND2_X1 U1003 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1004 ( .A(KEYINPUT47), .B(n902), .Z(n903) );
  NOR2_X1 U1005 ( .A1(n904), .A2(n903), .ZN(n943) );
  XNOR2_X1 U1006 ( .A(n943), .B(G162), .ZN(n905) );
  XNOR2_X1 U1007 ( .A(n906), .B(n905), .ZN(n915) );
  XOR2_X1 U1008 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n908) );
  XNOR2_X1 U1009 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n907) );
  XNOR2_X1 U1010 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1011 ( .A(n909), .B(KEYINPUT115), .Z(n913) );
  XOR2_X1 U1012 ( .A(n911), .B(n910), .Z(n912) );
  XNOR2_X1 U1013 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1014 ( .A(n915), .B(n914), .Z(n917) );
  XNOR2_X1 U1015 ( .A(G164), .B(G160), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n917), .B(n916), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n920), .ZN(G395) );
  XOR2_X1 U1019 ( .A(KEYINPUT118), .B(n921), .Z(n923) );
  XNOR2_X1 U1020 ( .A(G171), .B(n987), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n923), .B(n922), .ZN(n924) );
  XOR2_X1 U1022 ( .A(G286), .B(n924), .Z(n925) );
  XNOR2_X1 U1023 ( .A(n994), .B(n925), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(G37), .A2(n926), .ZN(G397) );
  NOR2_X1 U1025 ( .A1(G227), .A2(G229), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(G401), .A2(n928), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(G395), .A2(G397), .ZN(n929) );
  AND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(G319), .A2(n931), .ZN(G225) );
  XNOR2_X1 U1031 ( .A(KEYINPUT119), .B(G225), .ZN(G308) );
  INV_X1 U1033 ( .A(G120), .ZN(G236) );
  INV_X1 U1034 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(G325) );
  INV_X1 U1036 ( .A(G325), .ZN(G261) );
  INV_X1 U1037 ( .A(G108), .ZN(G238) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n981) );
  XOR2_X1 U1039 ( .A(G2084), .B(G160), .Z(n934) );
  NOR2_X1 U1040 ( .A1(n935), .A2(n934), .ZN(n939) );
  NOR2_X1 U1041 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1042 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1043 ( .A(KEYINPUT120), .B(n940), .ZN(n956) );
  NAND2_X1 U1044 ( .A1(n942), .A2(n941), .ZN(n948) );
  XOR2_X1 U1045 ( .A(G2072), .B(n943), .Z(n945) );
  XOR2_X1 U1046 ( .A(G164), .B(G2078), .Z(n944) );
  NOR2_X1 U1047 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1048 ( .A(KEYINPUT50), .B(n946), .Z(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G2090), .B(G162), .ZN(n949) );
  XNOR2_X1 U1051 ( .A(n949), .B(KEYINPUT121), .ZN(n950) );
  NOR2_X1 U1052 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1053 ( .A(KEYINPUT51), .B(n952), .Z(n953) );
  NAND2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(KEYINPUT122), .B(KEYINPUT52), .ZN(n957) );
  XNOR2_X1 U1057 ( .A(n958), .B(n957), .ZN(n959) );
  NAND2_X1 U1058 ( .A1(n981), .A2(n959), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(n960), .A2(G29), .ZN(n1040) );
  XNOR2_X1 U1060 ( .A(G2090), .B(G35), .ZN(n975) );
  XNOR2_X1 U1061 ( .A(G1996), .B(G32), .ZN(n962) );
  XNOR2_X1 U1062 ( .A(G33), .B(G2072), .ZN(n961) );
  NOR2_X1 U1063 ( .A1(n962), .A2(n961), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(G25), .B(n963), .ZN(n964) );
  NAND2_X1 U1065 ( .A1(n964), .A2(G28), .ZN(n968) );
  XOR2_X1 U1066 ( .A(G27), .B(n965), .Z(n966) );
  XNOR2_X1 U1067 ( .A(KEYINPUT123), .B(n966), .ZN(n967) );
  NOR2_X1 U1068 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1069 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1070 ( .A(G26), .B(G2067), .ZN(n971) );
  NOR2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1072 ( .A(KEYINPUT53), .B(n973), .ZN(n974) );
  NOR2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(n976), .B(KEYINPUT124), .ZN(n979) );
  XOR2_X1 U1075 ( .A(G2084), .B(G34), .Z(n977) );
  XNOR2_X1 U1076 ( .A(KEYINPUT54), .B(n977), .ZN(n978) );
  NAND2_X1 U1077 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1078 ( .A(n981), .B(n980), .ZN(n983) );
  INV_X1 U1079 ( .A(G29), .ZN(n982) );
  NAND2_X1 U1080 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n984), .ZN(n1038) );
  XNOR2_X1 U1082 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  NAND2_X1 U1083 ( .A1(G1971), .A2(G303), .ZN(n985) );
  NAND2_X1 U1084 ( .A1(n986), .A2(n985), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(n987), .B(G1348), .ZN(n989) );
  NAND2_X1 U1086 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(G1341), .B(n994), .ZN(n995) );
  NOR2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(n997), .B(G1956), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(G171), .B(G1961), .ZN(n998) );
  NAND2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G168), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1096 ( .A(KEYINPUT57), .B(n1002), .Z(n1003) );
  NOR2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1036) );
  INV_X1 U1100 ( .A(G16), .ZN(n1034) );
  XOR2_X1 U1101 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n1015) );
  XNOR2_X1 U1102 ( .A(G1986), .B(G24), .ZN(n1010) );
  XNOR2_X1 U1103 ( .A(G1971), .B(G22), .ZN(n1009) );
  NOR2_X1 U1104 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XOR2_X1 U1105 ( .A(G1976), .B(KEYINPUT126), .Z(n1011) );
  XNOR2_X1 U1106 ( .A(G23), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1107 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1108 ( .A(n1015), .B(n1014), .ZN(n1027) );
  XNOR2_X1 U1109 ( .A(G20), .B(n1016), .ZN(n1020) );
  XNOR2_X1 U1110 ( .A(G1341), .B(G19), .ZN(n1018) );
  XNOR2_X1 U1111 ( .A(G1981), .B(G6), .ZN(n1017) );
  NOR2_X1 U1112 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1113 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XOR2_X1 U1114 ( .A(KEYINPUT59), .B(G1348), .Z(n1021) );
  XNOR2_X1 U1115 ( .A(G4), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1116 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1117 ( .A(KEYINPUT125), .B(n1024), .ZN(n1025) );
  XNOR2_X1 U1118 ( .A(KEYINPUT60), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1119 ( .A1(n1027), .A2(n1026), .ZN(n1031) );
  XNOR2_X1 U1120 ( .A(G1966), .B(G21), .ZN(n1029) );
  XNOR2_X1 U1121 ( .A(G1961), .B(G5), .ZN(n1028) );
  NOR2_X1 U1122 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1123 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1124 ( .A(KEYINPUT61), .B(n1032), .Z(n1033) );
  NAND2_X1 U1125 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1126 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1127 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1128 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1129 ( .A(KEYINPUT62), .B(n1041), .Z(G311) );
  INV_X1 U1130 ( .A(G311), .ZN(G150) );
endmodule

