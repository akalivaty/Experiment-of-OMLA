//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n852, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G169gat), .B2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT23), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n209), .B1(G169gat), .B2(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n205), .B(new_n208), .C1(new_n210), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n217));
  OR2_X1    g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n203), .B1(new_n213), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n218), .A3(new_n217), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n209), .A2(G169gat), .A3(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n222), .A2(new_n225), .A3(new_n205), .A4(new_n208), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(new_n203), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n225), .A2(KEYINPUT25), .A3(new_n205), .A4(new_n208), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n231));
  INV_X1    g030(.A(G183gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n214), .A2(KEYINPUT66), .A3(new_n215), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n234), .A2(new_n236), .A3(new_n217), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n230), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n228), .A3(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(G127gat), .B(G134gat), .Z(new_n241));
  INV_X1    g040(.A(G113gat), .ZN(new_n242));
  INV_X1    g041(.A(G120gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G113gat), .A2(G120gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n241), .A2(new_n246), .A3(KEYINPUT1), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(G113gat), .A2(G120gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(G113gat), .A2(G120gat), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT69), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n244), .A2(new_n252), .A3(new_n245), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n256));
  NOR2_X1   g055(.A1(G127gat), .A2(G134gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT68), .B(G127gat), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(G134gat), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n255), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n256), .B1(new_n255), .B2(new_n259), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n248), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n231), .A2(new_n233), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT28), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT27), .B(G183gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(KEYINPUT27), .B(G183gat), .Z(new_n268));
  OAI21_X1  g067(.A(KEYINPUT28), .B1(new_n268), .B2(new_n263), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n270));
  OR3_X1    g069(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n225), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND4_X1   g071(.A1(new_n267), .A2(new_n269), .A3(new_n214), .A4(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n240), .A2(new_n262), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n262), .B1(new_n240), .B2(new_n274), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G227gat), .ZN(new_n278));
  INV_X1    g077(.A(G233gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n202), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n280), .ZN(new_n282));
  OAI211_X1 g081(.A(KEYINPUT34), .B(new_n282), .C1(new_n275), .C2(new_n276), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n275), .A2(new_n276), .A3(new_n282), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT71), .B1(new_n285), .B2(KEYINPUT33), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n240), .A2(new_n274), .ZN(new_n287));
  INV_X1    g086(.A(new_n262), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n240), .A2(new_n262), .A3(new_n274), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n280), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT33), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G15gat), .B(G43gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G71gat), .B(G99gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(new_n291), .B2(KEYINPUT32), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n286), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n286), .A2(new_n298), .A3(new_n301), .A4(new_n294), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n291), .A2(KEYINPUT32), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n297), .A2(new_n293), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n284), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G22gat), .B(G50gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G228gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G141gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT77), .B1(new_n312), .B2(G148gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(G141gat), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n313), .B(new_n316), .C1(G141gat), .C2(new_n315), .ZN(new_n317));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  INV_X1    g117(.A(G155gat), .ZN(new_n319));
  INV_X1    g118(.A(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n318), .B1(new_n321), .B2(KEYINPUT2), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G141gat), .B(G148gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n318), .B(new_n321), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G197gat), .B(G204gat), .ZN(new_n328));
  INV_X1    g127(.A(G218gat), .ZN(new_n329));
  INV_X1    g128(.A(G211gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT74), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G211gat), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT73), .B(KEYINPUT22), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n328), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G211gat), .B(G218gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n337), .B(new_n328), .C1(new_n334), .C2(new_n335), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n327), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n339), .A2(new_n340), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n323), .A2(new_n326), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n342), .B1(new_n347), .B2(KEYINPUT3), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n311), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT31), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n339), .A2(KEYINPUT82), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n336), .B2(new_n338), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n340), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n342), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n327), .B1(new_n359), .B2(new_n344), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n349), .A2(KEYINPUT83), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n348), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n310), .A3(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n351), .B(new_n354), .C1(new_n360), .C2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n311), .B1(new_n349), .B2(KEYINPUT83), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT3), .B1(new_n358), .B2(new_n342), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n363), .B(new_n367), .C1(new_n368), .C2(new_n327), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n354), .B1(new_n369), .B2(new_n351), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n309), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n351), .B1(new_n360), .B2(new_n364), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n353), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(new_n308), .A3(new_n365), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n306), .A2(new_n284), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(new_n300), .B2(new_n302), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n307), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n220), .A2(KEYINPUT65), .B1(new_n230), .B2(new_n238), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n273), .B1(new_n380), .B2(new_n228), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n381), .B2(KEYINPUT29), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n382), .B(new_n341), .C1(new_n379), .C2(new_n381), .ZN(new_n383));
  XNOR2_X1  g182(.A(G8gat), .B(G36gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(G64gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n385), .B(G92gat), .Z(new_n386));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n381), .B2(new_n379), .ZN(new_n388));
  INV_X1    g187(.A(new_n379), .ZN(new_n389));
  INV_X1    g188(.A(new_n228), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n234), .A2(new_n217), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n236), .A2(new_n237), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n229), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n227), .B1(new_n226), .B2(new_n203), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n390), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(KEYINPUT75), .B(new_n389), .C1(new_n395), .C2(new_n273), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n342), .B1(new_n395), .B2(new_n273), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n388), .A2(new_n396), .B1(new_n397), .B2(new_n379), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n383), .B(new_n386), .C1(new_n398), .C2(new_n341), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT75), .B1(new_n287), .B2(new_n389), .ZN(new_n402));
  AOI211_X1 g201(.A(new_n387), .B(new_n379), .C1(new_n240), .C2(new_n274), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n382), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n346), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n405), .A2(KEYINPUT30), .A3(new_n383), .A4(new_n386), .ZN(new_n406));
  INV_X1    g205(.A(new_n386), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n396), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n341), .B1(new_n408), .B2(new_n382), .ZN(new_n409));
  INV_X1    g208(.A(new_n383), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n401), .A2(new_n406), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G225gat), .A2(G233gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n323), .A2(new_n326), .A3(new_n344), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n344), .B1(new_n323), .B2(new_n326), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI211_X1 g218(.A(new_n414), .B(new_n416), .C1(new_n419), .C2(new_n262), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n327), .B(new_n248), .C1(new_n260), .C2(new_n261), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT4), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n255), .A2(new_n259), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT70), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n255), .A2(new_n256), .A3(new_n259), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n327), .A4(new_n248), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT80), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n422), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n288), .A2(KEYINPUT80), .A3(new_n427), .A4(new_n327), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n420), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n420), .A2(new_n430), .A3(KEYINPUT81), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n262), .A2(new_n347), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n438), .A2(new_n421), .ZN(new_n439));
  OAI211_X1 g238(.A(KEYINPUT79), .B(new_n414), .C1(new_n439), .C2(new_n415), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n428), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n419), .A2(new_n262), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n415), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT79), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n415), .B1(new_n438), .B2(new_n421), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n413), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n440), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G1gat), .B(G29gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(KEYINPUT0), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(G57gat), .ZN(new_n450));
  INV_X1    g249(.A(G85gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n447), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n447), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(KEYINPUT6), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n437), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n412), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n378), .A2(KEYINPUT86), .A3(KEYINPUT35), .A4(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n376), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n375), .B1(new_n303), .B2(new_n461), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n300), .A2(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n462), .B(new_n459), .C1(new_n284), .C2(new_n463), .ZN(new_n464));
  OR2_X1    g263(.A1(KEYINPUT86), .A2(KEYINPUT35), .ZN(new_n465));
  NAND2_X1  g264(.A1(KEYINPUT86), .A2(KEYINPUT35), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n455), .A2(new_n453), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n412), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n430), .A2(new_n431), .A3(new_n442), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n416), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT39), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n439), .B2(new_n415), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n470), .A2(new_n472), .A3(new_n416), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n475), .A2(KEYINPUT84), .A3(new_n452), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT84), .B1(new_n475), .B2(new_n452), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT40), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT40), .B(new_n474), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n469), .A2(KEYINPUT85), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT85), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n412), .A3(new_n468), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n475), .A2(new_n452), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n475), .A2(KEYINPUT84), .A3(new_n452), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT40), .B1(new_n489), .B2(new_n474), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n483), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n458), .A2(new_n454), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n409), .A2(new_n410), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT37), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n407), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n494), .A2(new_n495), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT38), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n386), .B1(new_n494), .B2(new_n495), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n389), .B1(new_n287), .B2(new_n342), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n381), .A2(new_n379), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n495), .B1(new_n503), .B2(new_n346), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n404), .A2(new_n341), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT38), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n500), .A2(new_n506), .B1(new_n494), .B2(new_n386), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n493), .A2(new_n499), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n375), .ZN(new_n509));
  AND4_X1   g308(.A1(new_n482), .A2(new_n491), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT36), .B1(new_n307), .B2(new_n377), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n375), .B1(new_n493), .B2(new_n412), .ZN(new_n512));
  INV_X1    g311(.A(new_n377), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n513), .B(new_n514), .C1(new_n284), .C2(new_n463), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n460), .B(new_n467), .C1(new_n510), .C2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G8gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT16), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(G1gat), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n521), .A2(KEYINPUT91), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(KEYINPUT91), .ZN(new_n523));
  OAI221_X1 g322(.A(new_n518), .B1(G1gat), .B2(new_n519), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  OR3_X1    g323(.A1(new_n519), .A2(KEYINPUT90), .A3(G1gat), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT90), .B1(new_n519), .B2(G1gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(G8gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G29gat), .ZN(new_n530));
  INV_X1    g329(.A(G36gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT14), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(G29gat), .B2(G36gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(G29gat), .A2(G36gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(KEYINPUT15), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT88), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n537), .B(KEYINPUT15), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n541), .A2(new_n536), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n529), .B1(new_n543), .B2(KEYINPUT17), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n542), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(KEYINPUT89), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT89), .B1(new_n545), .B2(new_n546), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n529), .A2(new_n545), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT18), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n551), .A4(new_n552), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT92), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(new_n529), .B2(new_n545), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n543), .A2(KEYINPUT92), .A3(new_n528), .A4(new_n524), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n559), .A3(new_n552), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n551), .B(KEYINPUT13), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n564));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G169gat), .B(G197gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT12), .Z(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n569), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n555), .A2(new_n571), .A3(new_n556), .A4(new_n562), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n517), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT41), .ZN(new_n576));
  NAND3_X1  g375(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT7), .ZN(new_n578));
  INV_X1    g377(.A(G99gat), .ZN(new_n579));
  INV_X1    g378(.A(G106gat), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT8), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT100), .B(G92gat), .Z(new_n582));
  OAI211_X1 g381(.A(new_n578), .B(new_n581), .C1(G85gat), .C2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G99gat), .B(G106gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(new_n545), .B2(new_n546), .ZN(new_n587));
  INV_X1    g386(.A(new_n549), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(new_n547), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n545), .A2(new_n585), .B1(KEYINPUT41), .B2(new_n575), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT101), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n548), .A2(new_n549), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n593), .B(new_n590), .C1(new_n594), .C2(new_n587), .ZN(new_n595));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT98), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n596), .B1(new_n592), .B2(new_n595), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n576), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT97), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n592), .A2(new_n595), .ZN(new_n603));
  INV_X1    g402(.A(new_n596), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n576), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n605), .A2(KEYINPUT98), .A3(new_n606), .A4(new_n597), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n600), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n602), .B1(new_n600), .B2(new_n607), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G71gat), .B(G78gat), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT93), .Z(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT94), .B(G57gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(G64gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT95), .Z(new_n617));
  INV_X1    g416(.A(G64gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(G57gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT96), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n612), .B(new_n614), .C1(new_n617), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G57gat), .B(G64gat), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n614), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n611), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n529), .B1(new_n625), .B2(KEYINPUT21), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n232), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n627), .B(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n625), .A2(KEYINPUT21), .ZN(new_n632));
  XNOR2_X1  g431(.A(G127gat), .B(G155gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n330), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n631), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n610), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n584), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT102), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n621), .A2(new_n624), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n586), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n621), .A2(new_n624), .A3(new_n585), .A4(new_n640), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n625), .A2(KEYINPUT10), .A3(new_n585), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT103), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n642), .B2(new_n644), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT104), .B(G120gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  NAND3_X1  g456(.A1(new_n651), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n649), .B1(new_n645), .B2(new_n646), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n660), .B2(new_n652), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(KEYINPUT105), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n663), .B(new_n659), .C1(new_n660), .C2(new_n652), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n638), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n574), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n492), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(G1gat), .Z(G1324gat));
  INV_X1    g468(.A(new_n412), .ZN(new_n670));
  OAI21_X1  g469(.A(G8gat), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n667), .A2(new_n670), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT16), .B(G8gat), .Z(new_n677));
  AND3_X1   g476(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n676), .B1(new_n675), .B2(new_n677), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n673), .B(new_n674), .C1(new_n678), .C2(new_n679), .ZN(G1325gat));
  AND2_X1   g479(.A1(new_n511), .A2(new_n515), .ZN(new_n681));
  OAI21_X1  g480(.A(G15gat), .B1(new_n667), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n307), .A2(new_n377), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n684), .A2(G15gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n682), .B1(new_n667), .B2(new_n685), .ZN(G1326gat));
  NOR2_X1   g485(.A1(new_n667), .A2(new_n509), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT43), .B(G22gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT107), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n687), .B(new_n689), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n637), .A2(new_n665), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n600), .A2(new_n607), .ZN(new_n692));
  INV_X1    g491(.A(new_n602), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n600), .A2(new_n602), .A3(new_n607), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n574), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(new_n530), .A3(new_n493), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT45), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n696), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT108), .B1(new_n510), .B2(new_n516), .ZN(new_n705));
  INV_X1    g504(.A(new_n516), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n491), .A2(new_n508), .A3(new_n482), .A4(new_n509), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n466), .B1(new_n464), .B2(new_n465), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT109), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n460), .A2(new_n714), .A3(new_n467), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n704), .B1(new_n710), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n517), .B2(new_n696), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n691), .A2(new_n573), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n493), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n702), .B1(new_n530), .B2(new_n724), .ZN(G1328gat));
  NOR3_X1   g524(.A1(new_n699), .A2(G36gat), .A3(new_n670), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT46), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n722), .A2(new_n412), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n729), .B2(new_n531), .ZN(G1329gat));
  INV_X1    g529(.A(new_n681), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n722), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n699), .A2(G43gat), .A3(new_n684), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  INV_X1    g536(.A(G43gat), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(new_n722), .B2(new_n731), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n739), .B2(new_n734), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n736), .A2(new_n740), .ZN(G1330gat));
  XNOR2_X1  g540(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n717), .A2(new_n719), .ZN(new_n743));
  INV_X1    g542(.A(new_n721), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(new_n375), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n509), .A2(G50gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n699), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n742), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n742), .ZN(new_n751));
  AOI211_X1 g550(.A(new_n751), .B(new_n748), .C1(new_n745), .C2(G50gat), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n750), .A2(new_n752), .ZN(G1331gat));
  NOR3_X1   g552(.A1(new_n510), .A2(KEYINPUT108), .A3(new_n516), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n707), .B1(new_n706), .B2(new_n708), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n460), .A2(new_n714), .A3(new_n467), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n714), .B1(new_n460), .B2(new_n467), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n754), .A2(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n665), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n638), .A2(new_n573), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n492), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n615), .ZN(G1332gat));
  NOR2_X1   g562(.A1(new_n761), .A2(new_n670), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  AND2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n764), .B2(new_n765), .ZN(G1333gat));
  NOR3_X1   g567(.A1(new_n761), .A2(G71gat), .A3(new_n684), .ZN(new_n769));
  INV_X1    g568(.A(new_n761), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n731), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(G71gat), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n375), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g574(.A1(new_n665), .A2(new_n451), .A3(new_n493), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT114), .Z(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n705), .A2(new_n709), .B1(new_n713), .B2(new_n715), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n637), .A2(new_n573), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n696), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n781), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n758), .A2(KEYINPUT51), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(KEYINPUT113), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(KEYINPUT113), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n777), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n780), .A2(new_n665), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT112), .Z(new_n790));
  NAND2_X1  g589(.A1(new_n743), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791), .B2(new_n492), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n792), .ZN(G1336gat));
  NOR2_X1   g592(.A1(new_n670), .A2(G92gat), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n759), .B(new_n795), .C1(new_n782), .C2(new_n784), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n790), .B(new_n412), .C1(new_n717), .C2(new_n719), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n582), .ZN(new_n799));
  XNOR2_X1  g598(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n798), .A2(new_n802), .A3(new_n582), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n798), .B2(new_n582), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n803), .A2(new_n804), .A3(new_n796), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n801), .B1(new_n805), .B2(new_n806), .ZN(G1337gat));
  NOR3_X1   g606(.A1(new_n684), .A2(G99gat), .A3(new_n759), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n786), .B2(new_n787), .ZN(new_n809));
  OAI21_X1  g608(.A(G99gat), .B1(new_n791), .B2(new_n681), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1338gat));
  NAND4_X1  g610(.A1(new_n785), .A2(new_n580), .A3(new_n375), .A4(new_n665), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n790), .B(new_n375), .C1(new_n717), .C2(new_n719), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G106gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(KEYINPUT117), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT53), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n812), .A2(KEYINPUT117), .A3(new_n817), .A4(new_n814), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1339gat));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n657), .B1(new_n660), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n651), .A2(KEYINPUT54), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n647), .A2(new_n650), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT55), .B(new_n821), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n826), .A2(new_n573), .A3(new_n658), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n560), .A2(new_n561), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n568), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n662), .A2(new_n572), .A3(new_n664), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n572), .A2(new_n831), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n664), .A4(new_n662), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n828), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n610), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n826), .A2(new_n834), .A3(new_n658), .A4(new_n827), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n696), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n636), .ZN(new_n843));
  INV_X1    g642(.A(new_n573), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n610), .A2(new_n637), .A3(new_n844), .A4(new_n759), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n492), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n670), .A3(new_n378), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n844), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(new_n242), .ZN(G1340gat));
  NOR2_X1   g648(.A1(new_n847), .A2(new_n759), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(new_n243), .ZN(G1341gat));
  NOR2_X1   g650(.A1(new_n847), .A2(new_n636), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(new_n258), .Z(G1342gat));
  AOI211_X1 g652(.A(new_n610), .B(new_n847), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n854));
  NOR2_X1   g653(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1343gat));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(KEYINPUT58), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n857), .A2(KEYINPUT58), .ZN(new_n859));
  INV_X1    g658(.A(new_n845), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n828), .A2(new_n832), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n610), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n841), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n860), .B1(new_n863), .B2(new_n636), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT57), .B1(new_n864), .B2(new_n509), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n839), .B1(new_n694), .B2(new_n695), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n610), .B2(new_n837), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n845), .B1(new_n867), .B2(new_n637), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n509), .A2(KEYINPUT57), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n731), .A2(new_n492), .A3(new_n412), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n865), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(G141gat), .B1(new_n872), .B2(new_n844), .ZN(new_n873));
  AND4_X1   g672(.A1(new_n670), .A2(new_n846), .A3(new_n375), .A4(new_n681), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n312), .A3(new_n573), .ZN(new_n875));
  AOI211_X1 g674(.A(new_n858), .B(new_n859), .C1(new_n873), .C2(new_n875), .ZN(new_n876));
  AND4_X1   g675(.A1(new_n857), .A2(new_n873), .A3(new_n875), .A4(KEYINPUT58), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(G1344gat));
  NAND3_X1  g677(.A1(new_n874), .A2(new_n315), .A3(new_n665), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n863), .A2(KEYINPUT120), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n636), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n863), .A2(KEYINPUT120), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n845), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n375), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n884), .A2(new_n869), .B1(KEYINPUT57), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n665), .A3(new_n871), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n880), .B1(new_n887), .B2(G148gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n759), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(KEYINPUT59), .A3(new_n315), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n879), .B1(new_n888), .B2(new_n890), .ZN(G1345gat));
  OAI21_X1  g690(.A(G155gat), .B1(new_n872), .B2(new_n636), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n319), .A3(new_n637), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT121), .ZN(G1346gat));
  OAI21_X1  g694(.A(G162gat), .B1(new_n872), .B2(new_n610), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n874), .A2(new_n320), .A3(new_n696), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1347gat));
  AND2_X1   g697(.A1(new_n378), .A2(new_n412), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n637), .B1(new_n838), .B2(new_n841), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n492), .B(new_n899), .C1(new_n900), .C2(new_n860), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(new_n206), .A3(new_n844), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT122), .B1(new_n868), .B2(new_n492), .ZN(new_n903));
  OAI211_X1 g702(.A(KEYINPUT122), .B(new_n492), .C1(new_n900), .C2(new_n860), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(new_n899), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n573), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n902), .B1(new_n908), .B2(new_n206), .ZN(G1348gat));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n207), .A3(new_n665), .ZN(new_n910));
  OAI21_X1  g709(.A(G176gat), .B1(new_n901), .B2(new_n759), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1349gat));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n493), .B1(new_n843), .B2(new_n845), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n914), .A2(new_n915), .A3(new_n637), .A4(new_n899), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT123), .B1(new_n901), .B2(new_n636), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(G183gat), .A3(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n636), .A2(new_n268), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n899), .B(new_n920), .C1(new_n903), .C2(new_n905), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n919), .B1(new_n918), .B2(new_n921), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n913), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n918), .A2(new_n921), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT124), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(KEYINPUT60), .A3(new_n922), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n928), .ZN(G1350gat));
  NAND3_X1  g728(.A1(new_n907), .A2(new_n264), .A3(new_n696), .ZN(new_n930));
  OAI21_X1  g729(.A(G190gat), .B1(new_n901), .B2(new_n610), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT61), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1351gat));
  NOR3_X1   g732(.A1(new_n731), .A2(new_n670), .A3(new_n509), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n934), .B1(new_n903), .B2(new_n905), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n935), .B(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(G197gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(new_n938), .A3(new_n573), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n731), .A2(new_n493), .A3(new_n670), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n886), .A2(new_n573), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G197gat), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n939), .A2(new_n942), .ZN(G1352gat));
  NAND3_X1  g742(.A1(new_n886), .A2(new_n665), .A3(new_n940), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n886), .A2(KEYINPUT126), .A3(new_n665), .A4(new_n940), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(G204gat), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n935), .A2(G204gat), .A3(new_n759), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n948), .A2(new_n951), .A3(new_n952), .ZN(G1353gat));
  AND3_X1   g752(.A1(new_n637), .A2(new_n331), .A3(new_n333), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n884), .A2(new_n869), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n885), .A2(KEYINPUT57), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n956), .A2(new_n637), .A3(new_n957), .A4(new_n940), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n886), .A2(new_n962), .A3(new_n940), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n696), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n962), .B1(new_n886), .B2(new_n940), .ZN(new_n965));
  OAI21_X1  g764(.A(G218gat), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n937), .A2(new_n329), .A3(new_n696), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1355gat));
endmodule


