//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  AND2_X1   g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G211gat), .A2(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G197gat), .B(G204gat), .Z(new_n207));
  NOR2_X1   g006(.A1(new_n204), .A2(KEYINPUT22), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(G197gat), .B(G204gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n210), .B(new_n211), .C1(KEYINPUT22), .C2(new_n204), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT29), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT3), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT78), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G141gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n220), .A3(G148gat), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G141gat), .ZN(new_n223));
  AND2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n221), .A2(new_n223), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G155gat), .B(G162gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n217), .A2(G148gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n230), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n216), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n224), .A2(new_n226), .ZN(new_n235));
  XNOR2_X1  g034(.A(G141gat), .B(G148gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(KEYINPUT2), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n217), .A2(G148gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT78), .B(G141gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(G148gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n224), .B1(new_n227), .B2(new_n226), .ZN(new_n241));
  OAI211_X1 g040(.A(KEYINPUT79), .B(new_n237), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n234), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n215), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n245), .B(new_n237), .C1(new_n240), .C2(new_n241), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n213), .B1(new_n246), .B2(new_n214), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n203), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n221), .A2(new_n223), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n228), .A2(new_n225), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n222), .A2(G141gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n227), .B1(new_n238), .B2(new_n251), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n249), .A2(new_n250), .B1(new_n252), .B2(new_n235), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT82), .B1(new_n215), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT29), .B1(new_n209), .B2(new_n212), .ZN(new_n256));
  OAI221_X1 g055(.A(new_n255), .B1(new_n229), .B2(new_n233), .C1(new_n256), .C2(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n246), .A2(new_n214), .ZN(new_n258));
  INV_X1    g057(.A(new_n213), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n203), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n254), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT31), .B(G50gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n248), .B2(new_n261), .ZN(new_n266));
  XNOR2_X1  g065(.A(G78gat), .B(G106gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(G22gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n265), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n248), .A2(new_n261), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n262), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n272), .B2(new_n264), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G226gat), .A2(G233gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n280), .A2(KEYINPUT67), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT67), .B1(new_n280), .B2(new_n281), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT27), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT27), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n286), .B1(new_n292), .B2(KEYINPUT28), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT27), .B(G183gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n295), .A3(new_n291), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n284), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G169gat), .ZN(new_n298));
  INV_X1    g097(.A(G176gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT23), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n302), .A3(new_n278), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n285), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n303), .B1(new_n307), .B2(KEYINPUT64), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT64), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n309), .A3(new_n306), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT25), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(KEYINPUT66), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n313), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n312), .A2(new_n314), .B1(new_n285), .B2(new_n304), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n302), .A2(KEYINPUT25), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT65), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n278), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n315), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n297), .B1(new_n311), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n276), .B1(new_n322), .B2(new_n214), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n300), .A2(new_n302), .A3(new_n278), .ZN(new_n325));
  AND2_X1   g124(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n285), .A2(new_n304), .B1(new_n326), .B2(G190gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n327), .B2(new_n309), .ZN(new_n328));
  INV_X1    g127(.A(new_n310), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n321), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n275), .B1(new_n332), .B2(new_n297), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n259), .B1(new_n323), .B2(new_n333), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n284), .A2(new_n293), .A3(new_n296), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n330), .B2(new_n331), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n275), .B1(new_n336), .B2(KEYINPUT29), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n276), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n213), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G8gat), .B(G36gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  NAND3_X1  g141(.A1(new_n334), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT30), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n234), .A2(KEYINPUT3), .A3(new_n242), .ZN(new_n347));
  INV_X1    g146(.A(G120gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G113gat), .ZN(new_n349));
  INV_X1    g148(.A(G113gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G120gat), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT1), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G127gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G134gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(KEYINPUT68), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G134gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G127gat), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n354), .A2(new_n358), .A3(KEYINPUT68), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n350), .A2(KEYINPUT69), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT69), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G113gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n364), .A3(G120gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT70), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n366), .A3(new_n349), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n354), .A2(new_n358), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n366), .B1(new_n365), .B2(new_n349), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n361), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n347), .A2(new_n373), .A3(new_n246), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n253), .B(new_n361), .C1(new_n372), .C2(new_n371), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n359), .A2(new_n352), .A3(new_n355), .ZN(new_n378));
  INV_X1    g177(.A(new_n349), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT69), .B(G113gat), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(G120gat), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n369), .B1(new_n381), .B2(new_n366), .ZN(new_n382));
  INV_X1    g181(.A(new_n372), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(KEYINPUT4), .A3(new_n253), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n374), .A2(new_n377), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT80), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n234), .A3(new_n242), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n375), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT5), .ZN(new_n392));
  OAI22_X1  g191(.A1(new_n386), .A2(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n375), .B(KEYINPUT4), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n394), .A2(KEYINPUT5), .A3(new_n389), .A4(new_n374), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT0), .ZN(new_n398));
  XNOR2_X1  g197(.A(G57gat), .B(G85gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n393), .A2(new_n395), .A3(new_n400), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n393), .A2(new_n395), .A3(new_n400), .ZN(new_n406));
  INV_X1    g205(.A(new_n404), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n346), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n334), .A2(new_n339), .ZN(new_n410));
  INV_X1    g209(.A(new_n342), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n334), .A2(new_n339), .A3(KEYINPUT30), .A4(new_n342), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT77), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n412), .B2(new_n413), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n274), .B1(new_n409), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n400), .B(KEYINPUT83), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n393), .A2(new_n395), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n404), .A3(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n421), .A2(new_n408), .A3(new_n343), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n323), .A2(new_n333), .A3(new_n259), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n213), .B1(new_n337), .B2(new_n338), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT37), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT37), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n334), .A2(new_n339), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n427), .A3(new_n411), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT38), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT38), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n425), .A2(new_n430), .A3(new_n427), .A4(new_n411), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT85), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n342), .B1(new_n410), .B2(KEYINPUT37), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n430), .A4(new_n427), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n422), .A2(new_n429), .A3(new_n432), .A4(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n274), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n386), .A2(new_n388), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n389), .B(new_n375), .C1(new_n243), .C2(new_n384), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n439), .A2(KEYINPUT39), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n419), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT39), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n386), .A2(new_n443), .A3(new_n388), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n441), .A2(KEYINPUT40), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n420), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT40), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n442), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n439), .A2(KEYINPUT39), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n388), .B2(new_n386), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n447), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT84), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n453), .B(new_n447), .C1(new_n448), .C2(new_n450), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n446), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n345), .A2(new_n412), .A3(new_n413), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n437), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n418), .B1(new_n436), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n307), .A2(KEYINPUT64), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(new_n310), .A3(new_n325), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n321), .B1(new_n460), .B2(new_n324), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n384), .B1(new_n461), .B2(new_n335), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n373), .B(new_n297), .C1(new_n311), .C2(new_n321), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G227gat), .ZN(new_n465));
  INV_X1    g264(.A(G233gat), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(KEYINPUT74), .A2(KEYINPUT34), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(KEYINPUT74), .A2(KEYINPUT34), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n467), .B2(new_n469), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n465), .A2(new_n466), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n462), .A2(new_n476), .A3(new_n463), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT71), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(KEYINPUT71), .A3(new_n478), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G43gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(G71gat), .B(G99gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n477), .B2(KEYINPUT32), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n485), .A2(new_n478), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n477), .A2(KEYINPUT32), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT72), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n477), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n487), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT36), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n487), .A2(new_n493), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT73), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT73), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n487), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n474), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT75), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n475), .B1(new_n496), .B2(KEYINPUT73), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(KEYINPUT75), .A3(new_n499), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n495), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n496), .A2(new_n474), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n494), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n458), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n413), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n342), .B1(new_n334), .B2(new_n339), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n274), .A2(new_n513), .A3(new_n345), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n403), .A2(new_n404), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n400), .B1(new_n393), .B2(new_n395), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(new_n407), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n517), .B2(new_n420), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT35), .B1(new_n519), .B2(new_n507), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n494), .A2(new_n274), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n502), .B2(new_n504), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n409), .A2(new_n417), .A3(KEYINPUT35), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n510), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G169gat), .B(G197gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G29gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT14), .B(G29gat), .Z(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(G36gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n538));
  NAND2_X1  g337(.A1(G43gat), .A2(G50gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT88), .B(G50gat), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n538), .B(new_n539), .C1(new_n540), .C2(G43gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(G43gat), .A2(G50gat), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n538), .B1(new_n543), .B2(new_n539), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n537), .A2(new_n544), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G15gat), .B(G22gat), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n549), .A2(G1gat), .ZN(new_n550));
  INV_X1    g349(.A(G8gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT16), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n549), .B1(new_n552), .B2(G1gat), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n551), .B1(new_n550), .B2(new_n553), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n548), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n558), .B(KEYINPUT13), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562));
  INV_X1    g361(.A(new_n547), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n544), .B1(new_n537), .B2(new_n541), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(KEYINPUT89), .A2(KEYINPUT17), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n562), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n546), .A2(new_n547), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n556), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT90), .B1(new_n548), .B2(new_n556), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(new_n556), .B2(new_n569), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n558), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT18), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n560), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n569), .A2(new_n556), .ZN(new_n578));
  INV_X1    g377(.A(new_n573), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n580), .A2(new_n571), .B1(G229gat), .B2(G233gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(KEYINPUT18), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n533), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n560), .B(new_n532), .C1(new_n575), .C2(new_n576), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT91), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(new_n581), .B2(KEYINPUT18), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n575), .A2(KEYINPUT91), .A3(new_n576), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n583), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n525), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT92), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n592));
  INV_X1    g391(.A(G57gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(G64gat), .ZN(new_n594));
  INV_X1    g393(.A(G64gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(G57gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n592), .B1(new_n597), .B2(KEYINPUT94), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(KEYINPUT94), .B2(new_n597), .ZN(new_n599));
  XOR2_X1   g398(.A(G71gat), .B(G78gat), .Z(new_n600));
  OR2_X1    g399(.A1(new_n600), .A2(KEYINPUT93), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(KEYINPUT93), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n600), .A2(new_n592), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n596), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n596), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n594), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n604), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n612));
  XNOR2_X1  g411(.A(G127gat), .B(G155gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  AOI211_X1 g413(.A(new_n555), .B(new_n554), .C1(new_n611), .C2(KEYINPUT21), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT96), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n616), .A2(new_n622), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT98), .B(G85gat), .Z(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT99), .B(G92gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G85gat), .A2(G92gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT7), .ZN(new_n630));
  INV_X1    g429(.A(G99gat), .ZN(new_n631));
  INV_X1    g430(.A(G106gat), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT8), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G99gat), .B(G106gat), .Z(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n569), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n636), .A2(new_n546), .A3(new_n547), .A4(new_n637), .ZN(new_n640));
  NAND2_X1  g439(.A1(G232gat), .A2(G233gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT97), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT41), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n640), .A2(KEYINPUT100), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT100), .B1(new_n640), .B2(new_n644), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n639), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n643), .A2(KEYINPUT41), .ZN(new_n651));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n639), .B(new_n648), .C1(new_n645), .C2(new_n646), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n655), .A2(KEYINPUT101), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(KEYINPUT101), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n653), .B1(new_n650), .B2(new_n654), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI211_X1 g459(.A(KEYINPUT102), .B(new_n653), .C1(new_n650), .C2(new_n654), .ZN(new_n661));
  OAI22_X1  g460(.A1(new_n656), .A2(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n638), .A2(new_n610), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n636), .A2(new_n637), .A3(new_n603), .A4(new_n609), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n667), .A2(new_n666), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n667), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(new_n671), .B2(new_n664), .ZN(new_n672));
  XOR2_X1   g471(.A(G120gat), .B(G148gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT103), .ZN(new_n674));
  XNOR2_X1  g473(.A(G176gat), .B(G204gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n668), .A2(new_n669), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n663), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n671), .A2(new_n664), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n676), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n625), .A2(new_n662), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n591), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n405), .A2(new_n408), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g488(.A(new_n551), .B1(new_n685), .B2(new_n456), .ZN(new_n690));
  INV_X1    g489(.A(new_n456), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT16), .B(G8gat), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n684), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT42), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(KEYINPUT42), .B2(new_n693), .ZN(G1325gat));
  INV_X1    g494(.A(new_n495), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n500), .A2(new_n501), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT75), .B1(new_n503), .B2(new_n499), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n509), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G15gat), .B1(new_n684), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n507), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n703), .A2(G15gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n684), .B2(new_n704), .ZN(G1326gat));
  NOR2_X1   g504(.A1(new_n684), .A2(new_n274), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT43), .B(G22gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  INV_X1    g507(.A(new_n682), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n625), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n662), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n591), .A2(new_n534), .A3(new_n687), .A4(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n406), .A2(new_n516), .A3(new_n407), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n345), .B1(new_n716), .B2(new_n515), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT77), .B1(new_n511), .B2(new_n512), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n412), .A2(new_n414), .A3(new_n413), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n437), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n429), .A2(new_n408), .A3(new_n343), .A4(new_n421), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n432), .A2(new_n435), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n445), .A2(new_n420), .ZN(new_n725));
  INV_X1    g524(.A(new_n454), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n453), .B1(new_n727), .B2(new_n447), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n456), .B(new_n725), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n274), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n721), .B1(new_n724), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n700), .B2(new_n699), .ZN(new_n732));
  INV_X1    g531(.A(new_n521), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n523), .B(new_n733), .C1(new_n697), .C2(new_n698), .ZN(new_n734));
  INV_X1    g533(.A(new_n520), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n662), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n711), .B1(new_n510), .B2(new_n524), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT44), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n589), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n710), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G29gat), .B1(new_n745), .B2(new_n686), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n713), .A2(new_n714), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n715), .A2(new_n746), .A3(new_n747), .ZN(G1328gat));
  NAND2_X1  g547(.A1(new_n591), .A2(new_n712), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n749), .A2(G36gat), .A3(new_n691), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n750), .A2(KEYINPUT46), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(KEYINPUT46), .ZN(new_n752));
  OAI21_X1  g551(.A(G36gat), .B1(new_n745), .B2(new_n691), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(G1329gat));
  INV_X1    g553(.A(new_n745), .ZN(new_n755));
  INV_X1    g554(.A(new_n701), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(G43gat), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(G43gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n749), .B2(new_n703), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1330gat));
  NAND4_X1  g561(.A1(new_n742), .A2(new_n540), .A3(new_n437), .A4(new_n744), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n749), .A2(new_n274), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n540), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g565(.A1(new_n623), .A2(new_n624), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n711), .A2(new_n743), .A3(new_n682), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT105), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n525), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n686), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(new_n593), .ZN(G1332gat));
  NOR2_X1   g571(.A1(new_n770), .A2(new_n691), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  AND2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n773), .B2(new_n774), .ZN(G1333gat));
  INV_X1    g576(.A(new_n770), .ZN(new_n778));
  INV_X1    g577(.A(G71gat), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n701), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT106), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n779), .B1(new_n770), .B2(new_n703), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g585(.A1(new_n778), .A2(new_n437), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g587(.A1(new_n767), .A2(new_n589), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n709), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n742), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n686), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT51), .B1(new_n740), .B2(new_n789), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n662), .B(new_n789), .C1(new_n732), .C2(new_n736), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT107), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT107), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n740), .A2(new_n798), .A3(KEYINPUT51), .A4(new_n789), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n794), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n687), .A2(new_n682), .A3(new_n626), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n793), .A2(new_n626), .B1(new_n800), .B2(new_n801), .ZN(G1336gat));
  OR3_X1    g601(.A1(new_n709), .A2(G92gat), .A3(new_n691), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT108), .Z(new_n804));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT51), .B1(new_n795), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n805), .B2(new_n795), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n797), .A2(new_n799), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(KEYINPUT110), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n739), .A2(new_n741), .A3(new_n456), .A4(new_n791), .ZN(new_n811));
  INV_X1    g610(.A(new_n627), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n809), .B2(KEYINPUT110), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT52), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n794), .ZN(new_n816));
  AOI211_X1 g615(.A(new_n711), .B(new_n790), .C1(new_n510), .C2(new_n524), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n798), .B1(new_n817), .B2(KEYINPUT51), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n795), .A2(KEYINPUT107), .A3(new_n796), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n804), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(KEYINPUT111), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n800), .B2(new_n804), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n811), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n627), .B1(new_n811), .B2(new_n827), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n825), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n826), .B1(new_n825), .B2(new_n830), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n815), .B1(new_n831), .B2(new_n832), .ZN(G1337gat));
  OAI21_X1  g632(.A(G99gat), .B1(new_n792), .B2(new_n701), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n507), .A2(new_n631), .A3(new_n682), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n834), .B1(new_n800), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT114), .ZN(G1338gat));
  NOR2_X1   g636(.A1(new_n792), .A2(new_n274), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n632), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n682), .A2(new_n632), .A3(new_n437), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n807), .B2(new_n808), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT53), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  OAI221_X1 g642(.A(new_n843), .B1(new_n800), .B2(new_n840), .C1(new_n838), .C2(new_n632), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(G1339gat));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n668), .A2(new_n669), .A3(new_n664), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n679), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n676), .B1(new_n670), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(KEYINPUT55), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n681), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT55), .B1(new_n848), .B2(new_n850), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n846), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n848), .A2(new_n850), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n857), .A2(KEYINPUT115), .A3(new_n681), .A4(new_n851), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n854), .A2(new_n589), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n580), .A2(G229gat), .A3(G233gat), .A4(new_n571), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n557), .A2(new_n559), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n530), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n586), .A2(new_n587), .ZN(new_n863));
  INV_X1    g662(.A(new_n584), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n682), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n662), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  AND4_X1   g666(.A1(new_n662), .A2(new_n854), .A3(new_n865), .A4(new_n858), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n625), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n711), .A2(new_n743), .A3(new_n709), .A4(new_n767), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n437), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n507), .B1(new_n871), .B2(KEYINPUT116), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n873), .B(new_n437), .C1(new_n869), .C2(new_n870), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n686), .A2(new_n456), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G113gat), .B1(new_n877), .B2(new_n743), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n686), .B1(new_n869), .B2(new_n870), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n879), .A2(new_n691), .A3(new_n522), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n380), .A3(new_n589), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n878), .A2(new_n881), .ZN(G1340gat));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n348), .A3(new_n682), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n884));
  INV_X1    g683(.A(new_n877), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n682), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n886), .B2(G120gat), .ZN(new_n887));
  AOI211_X1 g686(.A(KEYINPUT117), .B(new_n348), .C1(new_n885), .C2(new_n682), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n883), .B1(new_n887), .B2(new_n888), .ZN(G1341gat));
  OAI21_X1  g688(.A(G127gat), .B1(new_n877), .B2(new_n625), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n880), .A2(new_n353), .A3(new_n767), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1342gat));
  NAND3_X1  g691(.A1(new_n880), .A2(new_n357), .A3(new_n662), .ZN(new_n893));
  XOR2_X1   g692(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n894));
  XNOR2_X1  g693(.A(new_n893), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n877), .B2(new_n711), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1343gat));
  NOR2_X1   g696(.A1(new_n756), .A2(new_n274), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT120), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n879), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n691), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n743), .A2(G141gat), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OR3_X1    g704(.A1(new_n903), .A2(KEYINPUT121), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT121), .B1(new_n903), .B2(new_n905), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n701), .A2(new_n876), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n869), .A2(new_n870), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT57), .B1(new_n911), .B2(new_n437), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n852), .A2(new_n853), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n589), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n866), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n868), .B1(new_n711), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n870), .B1(new_n918), .B2(new_n767), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n274), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n912), .B2(new_n913), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n589), .B(new_n910), .C1(new_n914), .C2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n239), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n899), .A2(new_n456), .A3(new_n905), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n927), .B1(new_n924), .B2(new_n925), .ZN(new_n928));
  OAI22_X1  g727(.A1(new_n909), .A2(new_n926), .B1(new_n907), .B2(new_n928), .ZN(G1344gat));
  XNOR2_X1  g728(.A(new_n870), .B(KEYINPUT122), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n662), .B1(new_n866), .B2(new_n916), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n662), .A2(new_n865), .A3(new_n915), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n625), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n274), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(KEYINPUT123), .A3(new_n920), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n937), .B1(new_n934), .B2(KEYINPUT57), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n911), .A2(new_n921), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n682), .A3(new_n910), .ZN(new_n941));
  AND2_X1   g740(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n914), .A2(new_n923), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n910), .A2(new_n682), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(KEYINPUT59), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n941), .A2(new_n942), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT59), .B1(new_n903), .B2(new_n709), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n222), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1345gat));
  NAND2_X1  g748(.A1(new_n943), .A2(new_n910), .ZN(new_n950));
  OAI21_X1  g749(.A(G155gat), .B1(new_n950), .B2(new_n625), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n625), .A2(G155gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n903), .B2(new_n952), .ZN(G1346gat));
  OAI21_X1  g752(.A(G162gat), .B1(new_n950), .B2(new_n711), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n711), .A2(G162gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n903), .B2(new_n955), .ZN(G1347gat));
  NAND2_X1  g755(.A1(new_n911), .A2(new_n274), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n873), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n871), .A2(KEYINPUT116), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n687), .A2(new_n691), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT124), .Z(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n958), .A2(new_n507), .A3(new_n959), .A4(new_n962), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n963), .A2(new_n298), .A3(new_n743), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n911), .A2(new_n960), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n965), .A2(new_n522), .ZN(new_n966));
  AOI21_X1  g765(.A(G169gat), .B1(new_n966), .B2(new_n589), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n964), .A2(new_n967), .ZN(G1348gat));
  OAI21_X1  g767(.A(G176gat), .B1(new_n963), .B2(new_n709), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n299), .A3(new_n682), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1349gat));
  NAND3_X1  g770(.A1(new_n966), .A2(new_n294), .A3(new_n767), .ZN(new_n972));
  NOR4_X1   g771(.A1(new_n872), .A2(new_n874), .A3(new_n625), .A4(new_n961), .ZN(new_n973));
  OAI21_X1  g772(.A(G183gat), .B1(new_n973), .B2(KEYINPUT125), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n963), .A2(new_n975), .A3(new_n625), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n972), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT60), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT60), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n979), .B(new_n972), .C1(new_n974), .C2(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1350gat));
  NAND3_X1  g780(.A1(new_n966), .A2(new_n291), .A3(new_n662), .ZN(new_n982));
  OAI21_X1  g781(.A(G190gat), .B1(new_n963), .B2(new_n711), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n983), .A2(KEYINPUT61), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(KEYINPUT61), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  AND2_X1   g785(.A1(new_n965), .A2(new_n898), .ZN(new_n987));
  AOI21_X1  g786(.A(G197gat), .B1(new_n987), .B2(new_n589), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n756), .A2(new_n961), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n940), .A2(new_n989), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n589), .A2(G197gat), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(G1352gat));
  NAND2_X1  g791(.A1(new_n940), .A2(new_n989), .ZN(new_n993));
  OAI21_X1  g792(.A(G204gat), .B1(new_n993), .B2(new_n709), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n965), .A2(new_n898), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n995), .A2(G204gat), .A3(new_n709), .ZN(new_n996));
  XNOR2_X1  g795(.A(new_n996), .B(KEYINPUT62), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n994), .A2(new_n997), .ZN(G1353gat));
  OR3_X1    g797(.A1(new_n995), .A2(G211gat), .A3(new_n625), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n940), .A2(new_n767), .A3(new_n989), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n1000), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1001));
  AOI21_X1  g800(.A(KEYINPUT63), .B1(new_n1000), .B2(G211gat), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(G1354gat));
  INV_X1    g802(.A(G218gat), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1004), .B1(new_n995), .B2(new_n711), .ZN(new_n1005));
  XNOR2_X1  g804(.A(new_n1005), .B(KEYINPUT126), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n662), .A2(G218gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1007), .B1(new_n990), .B2(KEYINPUT127), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1006), .B1(new_n1008), .B2(new_n1010), .ZN(G1355gat));
endmodule


