//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n545, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  NAND2_X1  g030(.A1(G113), .A2(G2104), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT65), .B1(new_n457), .B2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n458), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n457), .A2(KEYINPUT65), .A3(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n466), .A2(G137), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n459), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n464), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND3_X1  g048(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n474));
  INV_X1    g049(.A(G136), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n467), .A2(G112), .ZN(new_n477));
  OAI22_X1  g052(.A1(new_n474), .A2(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n479), .B1(KEYINPUT3), .B2(new_n459), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n481));
  OAI211_X1 g056(.A(G2105), .B(new_n468), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n466), .A2(KEYINPUT66), .A3(G2105), .A4(new_n468), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n478), .B1(new_n486), .B2(G124), .ZN(G162));
  NAND4_X1  g062(.A1(new_n466), .A2(G138), .A3(new_n467), .A4(new_n468), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n467), .A2(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n461), .A2(KEYINPUT4), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n488), .A2(KEYINPUT4), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n482), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n491), .A2(new_n495), .ZN(G164));
  XNOR2_X1  g071(.A(KEYINPUT5), .B(G543), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  OR2_X1    g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT67), .B1(new_n501), .B2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(new_n499), .A3(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(G651), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n505), .A2(G88), .A3(new_n497), .A4(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n505), .A2(G50), .A3(G543), .A4(new_n506), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT68), .B1(new_n507), .B2(new_n508), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n500), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G166));
  AND3_X1   g089(.A1(new_n505), .A2(new_n497), .A3(new_n506), .ZN(new_n515));
  AND2_X1   g090(.A1(G63), .A2(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n515), .A2(G89), .B1(new_n497), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n503), .B1(KEYINPUT6), .B2(new_n499), .ZN(new_n518));
  NOR3_X1   g093(.A1(new_n501), .A2(KEYINPUT67), .A3(G651), .ZN(new_n519));
  OAI211_X1 g094(.A(G543), .B(new_n506), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT69), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n505), .A2(new_n522), .A3(G543), .A4(new_n506), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n521), .A2(G51), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT70), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n517), .A2(new_n524), .A3(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  XOR2_X1   g104(.A(KEYINPUT71), .B(G52), .Z(new_n530));
  NAND3_X1  g105(.A1(new_n521), .A2(new_n523), .A3(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n497), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(new_n499), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n515), .A2(G90), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  NAND3_X1  g111(.A1(new_n521), .A2(G43), .A3(new_n523), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n497), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n499), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT72), .B(G81), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n515), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n537), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G188));
  INV_X1    g124(.A(new_n520), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n550), .A2(KEYINPUT9), .A3(G53), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n497), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n499), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n515), .A2(G91), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n520), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n551), .A2(new_n553), .A3(new_n554), .A4(new_n557), .ZN(G299));
  XNOR2_X1  g133(.A(new_n509), .B(new_n510), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n559), .A2(KEYINPUT73), .A3(new_n500), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n513), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(G303));
  NAND2_X1  g138(.A1(new_n550), .A2(G49), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n515), .A2(G87), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT74), .ZN(G288));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  INV_X1    g144(.A(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT5), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT5), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n569), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n497), .A2(KEYINPUT75), .A3(G61), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT76), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n550), .A2(G48), .B1(new_n515), .B2(G86), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n579), .A2(new_n583), .A3(G651), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(G305));
  NAND3_X1  g160(.A1(new_n521), .A2(G47), .A3(new_n523), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n499), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n515), .A2(G85), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n515), .A2(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n515), .A2(KEYINPUT10), .A3(G92), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n521), .A2(G54), .A3(new_n523), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  XOR2_X1   g173(.A(KEYINPUT77), .B(G66), .Z(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n574), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n591), .B1(new_n602), .B2(G868), .ZN(G321));
  XOR2_X1   g178(.A(G321), .B(KEYINPUT78), .Z(G284));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT79), .ZN(G148));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n609), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g190(.A(new_n474), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G135), .ZN(new_n617));
  OR2_X1    g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n486), .B2(G123), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2096), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n623));
  NOR3_X1   g198(.A1(new_n457), .A2(new_n459), .A3(G2105), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n623), .B(new_n624), .Z(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT13), .B(G2100), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n622), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT15), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2435), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XOR2_X1   g208(.A(G2443), .B(G2446), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G1341), .B(G1348), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G14), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n644), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n646), .A2(new_n647), .ZN(new_n653));
  AOI21_X1  g228(.A(KEYINPUT18), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n651), .B(new_n654), .Z(G227));
  XNOR2_X1  g230(.A(G1961), .B(G1966), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT81), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  AND2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1971), .B(G1976), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n657), .A2(new_n658), .ZN(new_n664));
  AOI22_X1  g239(.A1(new_n662), .A2(new_n663), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  OR3_X1    g240(.A1(new_n659), .A2(new_n664), .A3(new_n661), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n666), .C1(new_n663), .C2(new_n662), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT82), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(new_n673), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G229));
  NAND2_X1  g250(.A1(G115), .A2(G2104), .ZN(new_n676));
  INV_X1    g251(.A(G127), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(new_n461), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT92), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G2105), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n616), .A2(G139), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n470), .A2(G103), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G29), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G29), .B2(G33), .ZN(new_n688));
  INV_X1    g263(.A(G2072), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(G171), .A2(G16), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G5), .B2(G16), .ZN(new_n693));
  INV_X1    g268(.A(G1961), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT85), .B(G16), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G19), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n543), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G1341), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n690), .A2(new_n691), .A3(new_n695), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n616), .A2(G141), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n470), .A2(G105), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT26), .Z(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT93), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n486), .B2(G129), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n486), .A2(new_n707), .A3(G129), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n706), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G29), .B2(G32), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT27), .B(G1996), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G35), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G162), .B2(new_n717), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G2090), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n701), .A2(new_n716), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n693), .A2(new_n694), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT96), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT96), .ZN(new_n726));
  NOR2_X1   g301(.A1(G27), .A2(G29), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G164), .B2(G29), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n725), .A2(new_n726), .B1(G2078), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n602), .A2(G16), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G4), .B2(G16), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT88), .B(G1348), .Z(new_n732));
  OAI22_X1  g307(.A1(new_n731), .A2(new_n732), .B1(G2078), .B2(new_n728), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n731), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G21), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G168), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT94), .B(G1966), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n729), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT89), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n486), .A2(G128), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n467), .A2(G116), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G140), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n474), .B2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n740), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G128), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n484), .B2(new_n485), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n751), .A2(KEYINPUT89), .A3(new_n747), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(new_n717), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n717), .A2(G26), .ZN(new_n755));
  OAI21_X1  g330(.A(KEYINPUT28), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(KEYINPUT28), .B2(new_n755), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT90), .B(G2067), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n697), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT98), .B(KEYINPUT23), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G299), .ZN(new_n763));
  INV_X1    g338(.A(G16), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT99), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1956), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n621), .A2(G29), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G28), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT95), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n771), .B(new_n717), .C1(new_n769), .C2(G28), .ZN(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  AND2_X1   g348(.A1(KEYINPUT24), .A2(G34), .ZN(new_n774));
  NOR2_X1   g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n774), .A2(new_n775), .A3(G29), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n472), .B2(G29), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n768), .B(new_n772), .C1(new_n773), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n713), .B2(new_n715), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n723), .A2(new_n739), .A3(new_n759), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n764), .A2(G6), .ZN(new_n782));
  INV_X1    g357(.A(G305), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n764), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT32), .B(G1981), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT86), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n784), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n697), .A2(G22), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G166), .B2(new_n697), .ZN(new_n789));
  INV_X1    g364(.A(G1971), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G16), .A2(G23), .ZN(new_n792));
  INV_X1    g367(.A(new_n567), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT33), .B(G1976), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n787), .A2(new_n791), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT34), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n697), .A2(G24), .ZN(new_n799));
  INV_X1    g374(.A(G290), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n697), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n797), .A2(KEYINPUT34), .B1(G1986), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(G1986), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G25), .ZN(new_n805));
  OAI21_X1  g380(.A(KEYINPUT83), .B1(new_n805), .B2(G29), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n805), .A2(KEYINPUT83), .A3(G29), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n486), .A2(G119), .ZN(new_n808));
  INV_X1    g383(.A(G131), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n467), .A2(G107), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n474), .A2(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n806), .B(new_n807), .C1(new_n813), .C2(new_n717), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT35), .B(G1991), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT84), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n814), .B(new_n816), .Z(new_n817));
  NAND4_X1  g392(.A1(new_n798), .A2(new_n802), .A3(new_n804), .A4(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT87), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(KEYINPUT36), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n781), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n818), .B1(new_n819), .B2(KEYINPUT36), .ZN(new_n822));
  INV_X1    g397(.A(new_n820), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n777), .A2(new_n773), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT31), .B(G11), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n821), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n699), .A2(G1341), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(G311));
  AND2_X1   g404(.A1(new_n821), .A2(new_n824), .ZN(new_n830));
  INV_X1    g405(.A(new_n828), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n830), .A2(new_n831), .A3(new_n825), .A4(new_n826), .ZN(G150));
  NAND3_X1  g407(.A1(new_n521), .A2(G55), .A3(new_n523), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n571), .A2(new_n573), .A3(G67), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n499), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n515), .B2(G93), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n833), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n833), .B2(new_n837), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  OAI21_X1  g418(.A(new_n542), .B1(new_n839), .B2(new_n840), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT101), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n833), .A2(new_n837), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n543), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(new_n542), .C1(new_n839), .C2(new_n840), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n609), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n850), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT39), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n853), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n843), .B1(new_n856), .B2(G860), .ZN(G145));
  XNOR2_X1  g432(.A(new_n621), .B(new_n472), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G162), .ZN(new_n859));
  INV_X1    g434(.A(G142), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n467), .A2(G118), .ZN(new_n862));
  OAI22_X1  g437(.A1(new_n474), .A2(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n486), .B2(G130), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n813), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n859), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n867));
  INV_X1    g442(.A(new_n706), .ZN(new_n868));
  INV_X1    g443(.A(new_n710), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n869), .B2(new_n708), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n741), .A2(new_n740), .A3(new_n748), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n491), .A2(new_n495), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT89), .B1(new_n751), .B2(new_n747), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n872), .B1(new_n871), .B2(new_n873), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n877));
  OAI21_X1  g452(.A(G164), .B1(new_n749), .B2(new_n752), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n711), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n877), .B1(new_n876), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n685), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n685), .B1(new_n876), .B2(new_n880), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n867), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n874), .A2(new_n875), .A3(new_n870), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n711), .B1(new_n878), .B2(new_n879), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT103), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT104), .B1(new_n891), .B2(new_n685), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n886), .A2(new_n625), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n625), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n686), .B1(new_n889), .B2(new_n890), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT104), .B1(new_n895), .B2(new_n884), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n883), .A2(new_n867), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n866), .B1(new_n893), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n625), .B1(new_n886), .B2(new_n892), .ZN(new_n901));
  INV_X1    g476(.A(new_n866), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n896), .A2(new_n894), .A3(new_n897), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g481(.A(new_n850), .B(new_n612), .Z(new_n907));
  NAND2_X1  g482(.A1(new_n602), .A2(new_n763), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n851), .A2(G299), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n851), .A2(G299), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n851), .A2(G299), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT41), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n908), .A2(new_n909), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(KEYINPUT105), .B2(KEYINPUT42), .ZN(new_n920));
  NAND2_X1  g495(.A1(G166), .A2(new_n793), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n513), .A2(new_n567), .ZN(new_n922));
  AOI21_X1  g497(.A(G290), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n922), .A3(G290), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n924), .A2(new_n783), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n783), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n930), .B(new_n931), .C1(new_n911), .C2(new_n918), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n920), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n920), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(G868), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n841), .A2(new_n605), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(G295));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n937), .ZN(G331));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n940));
  XNOR2_X1  g515(.A(G286), .B(G301), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n850), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n845), .A2(new_n941), .A3(new_n847), .A4(new_n849), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT106), .B1(new_n850), .B2(new_n942), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n945), .A2(new_n910), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n944), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n917), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n929), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(KEYINPUT106), .ZN(new_n952));
  INV_X1    g527(.A(new_n910), .ZN(new_n953));
  INV_X1    g528(.A(new_n946), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n928), .A3(new_n949), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n956), .A3(new_n900), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(new_n900), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n914), .A2(KEYINPUT108), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n910), .A2(new_n962), .A3(KEYINPUT41), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n916), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT107), .A4(new_n915), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n961), .A2(new_n963), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n945), .B2(new_n946), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n943), .A2(new_n953), .A3(new_n944), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n928), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n960), .A2(new_n958), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT44), .B1(new_n959), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  NOR4_X1   g548(.A1(new_n960), .A2(new_n973), .A3(KEYINPUT43), .A4(new_n970), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT109), .ZN(new_n976));
  INV_X1    g551(.A(new_n960), .ZN(new_n977));
  INV_X1    g552(.A(new_n970), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n958), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n974), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n972), .B1(new_n980), .B2(KEYINPUT44), .ZN(G397));
  NAND4_X1  g556(.A1(new_n464), .A2(G40), .A3(new_n469), .A4(new_n471), .ZN(new_n982));
  INV_X1    g557(.A(G1384), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n491), .B2(new_n495), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(KEYINPUT45), .B(new_n983), .C1(new_n491), .C2(new_n495), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT56), .B(G2072), .Z(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n990), .A2(KEYINPUT120), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(KEYINPUT120), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n872), .A2(KEYINPUT116), .A3(new_n993), .A4(new_n983), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n993), .B(new_n983), .C1(new_n491), .C2(new_n495), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n999));
  INV_X1    g574(.A(new_n982), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT115), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n982), .B1(new_n984), .B2(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n998), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n991), .B(new_n992), .C1(new_n1006), .C2(G1956), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1008));
  XNOR2_X1  g583(.A(G299), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n995), .B(KEYINPUT116), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1012));
  AOI211_X1 g587(.A(KEYINPUT115), .B(new_n982), .C1(new_n984), .C2(KEYINPUT50), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1956), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1009), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n991), .A4(new_n992), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1010), .A2(KEYINPUT61), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT61), .B1(new_n1010), .B2(new_n1018), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n872), .A2(new_n1000), .A3(KEYINPUT121), .A4(new_n983), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT121), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n984), .B2(new_n982), .ZN(new_n1023));
  INV_X1    g598(.A(G2067), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1348), .B1(new_n1003), .B2(new_n995), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n851), .A2(KEYINPUT123), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT123), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n602), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1027), .A2(KEYINPUT60), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT60), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n999), .A2(new_n1000), .A3(new_n995), .ZN(new_n1034));
  INV_X1    g609(.A(G1348), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n1030), .A3(new_n1037), .A4(KEYINPUT60), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(KEYINPUT123), .A3(new_n851), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1031), .A2(new_n1033), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n984), .A2(new_n985), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1041), .A2(new_n1000), .A3(new_n987), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G1996), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT58), .B(G1341), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n543), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT59), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(new_n543), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1040), .A2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1019), .A2(new_n1020), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1027), .A2(new_n851), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1018), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1014), .A2(new_n1015), .B1(KEYINPUT120), .B2(new_n990), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1017), .B1(new_n1058), .B2(new_n991), .ZN(new_n1059));
  OAI211_X1 g634(.A(KEYINPUT122), .B(new_n1018), .C1(new_n1059), .C2(new_n1054), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT124), .B1(new_n1052), .B2(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n986), .A2(KEYINPUT125), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n986), .B2(KEYINPUT125), .ZN(new_n1065));
  INV_X1    g640(.A(G2078), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .A4(new_n987), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n986), .A2(new_n1066), .A3(new_n987), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1068), .A2(new_n1064), .B1(new_n1034), .B2(new_n694), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(G301), .A3(new_n1069), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n1068), .A2(new_n1064), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1071), .A2(new_n1069), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1072), .B2(G301), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1042), .A2(new_n737), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT117), .B(G2084), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1003), .A2(new_n995), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1076), .B1(new_n1080), .B2(G286), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1077), .A2(new_n1079), .A3(G168), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G8), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1076), .B1(new_n1082), .B2(G8), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1075), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(G301), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1087), .A2(KEYINPUT126), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1074), .B1(new_n1072), .B2(G301), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(KEYINPUT126), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1034), .A2(G2090), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1971), .B1(new_n986), .B2(new_n987), .ZN(new_n1093));
  OAI21_X1  g668(.A(G8), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G303), .A2(G8), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1094), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G8), .ZN(new_n1101));
  INV_X1    g676(.A(new_n984), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n1000), .ZN(new_n1103));
  NAND2_X1  g678(.A1(G305), .A2(G1981), .ZN(new_n1104));
  INV_X1    g679(.A(G1981), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n581), .A2(new_n1105), .A3(new_n582), .A4(new_n584), .ZN(new_n1106));
  OR2_X1    g681(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n1110));
  OAI211_X1 g685(.A(new_n1103), .B(new_n1108), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n793), .A2(G1976), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1103), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT52), .ZN(new_n1114));
  INV_X1    g689(.A(G1976), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT52), .B1(G288), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(new_n1103), .A3(new_n1112), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1111), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1014), .A2(G2090), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1093), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1101), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1100), .B(new_n1119), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1086), .A2(new_n1091), .A3(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1040), .A2(new_n1050), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1010), .A2(KEYINPUT61), .A3(new_n1018), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1130), .A2(new_n1131), .A3(new_n1057), .A4(new_n1060), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1062), .A2(new_n1125), .A3(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1094), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT118), .B1(new_n1134), .B2(new_n1118), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1114), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1110), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1109), .B2(new_n1107), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1138), .B2(new_n1103), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1094), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1139), .A2(new_n1140), .A3(new_n1117), .A4(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1080), .A2(G8), .A3(G168), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1099), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1135), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT63), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1138), .A2(G1976), .A3(G288), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1106), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1103), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT62), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1072), .A2(G301), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1153), .B(new_n1154), .C1(new_n1083), .C2(new_n1081), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1143), .A2(KEYINPUT63), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1124), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1100), .A2(new_n1118), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1150), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1133), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n753), .A2(new_n1024), .ZN(new_n1162));
  OAI21_X1  g737(.A(G2067), .B1(new_n749), .B2(new_n752), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1041), .A2(new_n982), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT111), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n870), .B(G1996), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1165), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT112), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1167), .A2(KEYINPUT112), .A3(new_n1169), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n813), .B(new_n816), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n1165), .ZN(new_n1175));
  INV_X1    g750(.A(G1986), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n800), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT110), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1176), .B2(new_n800), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n1165), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1172), .A2(new_n1173), .A3(new_n1175), .A4(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT113), .Z(new_n1182));
  NAND2_X1  g757(.A1(new_n1161), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1165), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n808), .A2(new_n816), .A3(new_n812), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1172), .A2(new_n1173), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1184), .B1(new_n1186), .B2(new_n1162), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1178), .A2(new_n1184), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT48), .Z(new_n1189));
  AND4_X1   g764(.A1(new_n1172), .A2(new_n1189), .A3(new_n1173), .A4(new_n1175), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1164), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1192), .A2(KEYINPUT46), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1191), .B(new_n711), .C1(G1996), .C2(new_n1193), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n1184), .A2(G1996), .ZN(new_n1195));
  XOR2_X1   g770(.A(KEYINPUT127), .B(KEYINPUT46), .Z(new_n1196));
  AOI22_X1  g771(.A1(new_n1194), .A2(new_n1165), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT47), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1187), .A2(new_n1190), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1183), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g775(.A(G227), .ZN(new_n1202));
  NAND3_X1  g776(.A1(new_n905), .A2(new_n1202), .A3(new_n674), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n642), .A2(G319), .ZN(new_n1204));
  NOR3_X1   g778(.A1(new_n980), .A2(new_n1203), .A3(new_n1204), .ZN(G308));
  AND2_X1   g779(.A1(new_n905), .A2(new_n674), .ZN(new_n1206));
  INV_X1    g780(.A(new_n1204), .ZN(new_n1207));
  NAND4_X1  g781(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT109), .A4(new_n958), .ZN(new_n1208));
  AOI21_X1  g782(.A(new_n973), .B1(new_n957), .B2(KEYINPUT43), .ZN(new_n1209));
  NOR3_X1   g783(.A1(new_n960), .A2(KEYINPUT43), .A3(new_n970), .ZN(new_n1210));
  OAI21_X1  g784(.A(new_n1208), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND4_X1  g785(.A1(new_n1206), .A2(new_n1207), .A3(new_n1202), .A4(new_n1211), .ZN(G225));
endmodule


