

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779;

  BUF_X1 U377 ( .A(n567), .Z(n588) );
  AND2_X1 U378 ( .A1(n542), .A2(n476), .ZN(n708) );
  NOR2_X1 U379 ( .A1(n749), .A2(G902), .ZN(n472) );
  BUF_X1 U380 ( .A(G116), .Z(n356) );
  INV_X1 U381 ( .A(KEYINPUT64), .ZN(n458) );
  AND2_X2 U382 ( .A1(n726), .A2(n437), .ZN(n436) );
  AND2_X2 U383 ( .A1(n428), .A2(n427), .ZN(n426) );
  XNOR2_X1 U384 ( .A(n355), .B(n506), .ZN(n467) );
  NAND2_X1 U385 ( .A1(n511), .A2(G221), .ZN(n355) );
  XNOR2_X2 U386 ( .A(n522), .B(n521), .ZN(n761) );
  NAND2_X2 U387 ( .A1(n442), .A2(n440), .ZN(n552) );
  NAND2_X2 U388 ( .A1(n383), .A2(n648), .ZN(n655) );
  NAND2_X1 U389 ( .A1(n369), .A2(n368), .ZN(n374) );
  NOR2_X1 U390 ( .A1(n379), .A2(n414), .ZN(n413) );
  XNOR2_X1 U391 ( .A(n400), .B(n412), .ZN(n399) );
  XNOR2_X1 U392 ( .A(n642), .B(KEYINPUT46), .ZN(n387) );
  NOR2_X1 U393 ( .A1(n625), .A2(KEYINPUT85), .ZN(n626) );
  INV_X1 U394 ( .A(n588), .ZN(n357) );
  XNOR2_X1 U395 ( .A(n418), .B(n557), .ZN(n567) );
  NAND2_X1 U396 ( .A1(n614), .A2(n362), .ZN(n418) );
  AND2_X1 U397 ( .A1(n367), .A2(n443), .ZN(n442) );
  BUF_X1 U398 ( .A(n541), .Z(n607) );
  XNOR2_X1 U399 ( .A(n510), .B(n509), .ZN(n558) );
  XNOR2_X1 U400 ( .A(n467), .B(n466), .ZN(n749) );
  XNOR2_X1 U401 ( .A(n439), .B(n438), .ZN(n769) );
  XNOR2_X1 U402 ( .A(KEYINPUT10), .B(G125), .ZN(n439) );
  XNOR2_X1 U403 ( .A(G110), .B(G137), .ZN(n461) );
  XOR2_X1 U404 ( .A(G128), .B(G119), .Z(n464) );
  XOR2_X1 U405 ( .A(G131), .B(KEYINPUT68), .Z(n495) );
  NAND2_X1 U406 ( .A1(n697), .A2(KEYINPUT2), .ZN(n358) );
  AND2_X1 U407 ( .A1(n755), .A2(n770), .ZN(n697) );
  BUF_X1 U408 ( .A(n761), .Z(n359) );
  INV_X1 U409 ( .A(n748), .ZN(n360) );
  AND2_X2 U410 ( .A1(n655), .A2(n358), .ZN(n662) );
  XNOR2_X2 U411 ( .A(n472), .B(n471), .ZN(n542) );
  AND2_X1 U412 ( .A1(n629), .A2(n363), .ZN(n393) );
  XNOR2_X1 U413 ( .A(n492), .B(n491), .ZN(n548) );
  XNOR2_X1 U414 ( .A(n456), .B(n656), .ZN(n541) );
  XNOR2_X1 U415 ( .A(G110), .B(G107), .ZN(n485) );
  XNOR2_X1 U416 ( .A(n518), .B(n517), .ZN(n671) );
  XNOR2_X1 U417 ( .A(n531), .B(n455), .ZN(n768) );
  XNOR2_X1 U418 ( .A(KEYINPUT69), .B(G137), .ZN(n453) );
  INV_X1 U419 ( .A(n671), .ZN(n375) );
  NAND2_X1 U420 ( .A1(n393), .A2(n382), .ZN(n386) );
  AND2_X1 U421 ( .A1(n387), .A2(n392), .ZN(n382) );
  NAND2_X1 U422 ( .A1(n390), .A2(KEYINPUT48), .ZN(n389) );
  NAND2_X1 U423 ( .A1(n401), .A2(n602), .ZN(n400) );
  NAND2_X1 U424 ( .A1(n770), .A2(n415), .ZN(n414) );
  NAND2_X1 U425 ( .A1(n603), .A2(KEYINPUT86), .ZN(n415) );
  XNOR2_X1 U426 ( .A(KEYINPUT65), .B(KEYINPUT81), .ZN(n450) );
  XOR2_X1 U427 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n523) );
  XNOR2_X1 U428 ( .A(n508), .B(G475), .ZN(n509) );
  NAND2_X1 U429 ( .A1(n587), .A2(n420), .ZN(n566) );
  INV_X1 U430 ( .A(n595), .ZN(n420) );
  AND2_X1 U431 ( .A1(n431), .A2(n424), .ZN(n423) );
  AND2_X1 U432 ( .A1(n371), .A2(n364), .ZN(n369) );
  NAND2_X1 U433 ( .A1(n662), .A2(n372), .ZN(n371) );
  INV_X1 U434 ( .A(n741), .ZN(n748) );
  XNOR2_X1 U435 ( .A(n768), .B(n489), .ZN(n744) );
  INV_X1 U436 ( .A(G953), .ZN(n754) );
  NOR2_X1 U437 ( .A1(n779), .A2(n778), .ZN(n642) );
  XNOR2_X1 U438 ( .A(n409), .B(n408), .ZN(n717) );
  INV_X1 U439 ( .A(KEYINPUT104), .ZN(n408) );
  INV_X1 U440 ( .A(n444), .ZN(n435) );
  INV_X1 U441 ( .A(KEYINPUT88), .ZN(n412) );
  INV_X1 U442 ( .A(G140), .ZN(n438) );
  XNOR2_X1 U443 ( .A(n411), .B(n410), .ZN(n514) );
  XNOR2_X1 U444 ( .A(KEYINPUT7), .B(KEYINPUT101), .ZN(n410) );
  XNOR2_X1 U445 ( .A(n512), .B(KEYINPUT9), .ZN(n411) );
  XNOR2_X1 U446 ( .A(G107), .B(G134), .ZN(n512) );
  XNOR2_X1 U447 ( .A(G122), .B(G113), .ZN(n496) );
  XNOR2_X1 U448 ( .A(G143), .B(G104), .ZN(n497) );
  XOR2_X1 U449 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n498) );
  XNOR2_X1 U450 ( .A(KEYINPUT67), .B(G101), .ZN(n483) );
  XNOR2_X1 U451 ( .A(n548), .B(n547), .ZN(n565) );
  INV_X1 U452 ( .A(n607), .ZN(n705) );
  NOR2_X2 U453 ( .A1(n391), .A2(n388), .ZN(n770) );
  NAND2_X1 U454 ( .A1(n389), .A2(n646), .ZN(n388) );
  NOR2_X1 U455 ( .A1(n375), .A2(n670), .ZN(n372) );
  XNOR2_X1 U456 ( .A(n761), .B(n530), .ZN(n366) );
  INV_X1 U457 ( .A(KEYINPUT41), .ZN(n637) );
  XNOR2_X1 U458 ( .A(n690), .B(KEYINPUT103), .ZN(n643) );
  BUF_X1 U459 ( .A(n565), .Z(n707) );
  AND2_X1 U460 ( .A1(n394), .A2(n494), .ZN(n632) );
  XNOR2_X1 U461 ( .A(n395), .B(KEYINPUT30), .ZN(n394) );
  NOR2_X1 U462 ( .A1(n607), .A2(n396), .ZN(n395) );
  XNOR2_X1 U463 ( .A(n558), .B(n381), .ZN(n591) );
  INV_X1 U464 ( .A(KEYINPUT100), .ZN(n381) );
  NAND2_X1 U465 ( .A1(n567), .A2(n559), .ZN(n561) );
  INV_X1 U466 ( .A(n707), .ZN(n594) );
  XNOR2_X1 U467 ( .A(n541), .B(n540), .ZN(n595) );
  NAND2_X1 U468 ( .A1(n425), .A2(n423), .ZN(n422) );
  XOR2_X1 U469 ( .A(n749), .B(KEYINPUT125), .Z(n750) );
  XNOR2_X1 U470 ( .A(n374), .B(n373), .ZN(G63) );
  INV_X1 U471 ( .A(KEYINPUT124), .ZN(n373) );
  XNOR2_X1 U472 ( .A(n744), .B(n743), .ZN(n745) );
  NAND2_X1 U473 ( .A1(n445), .A2(n754), .ZN(n737) );
  AND2_X1 U474 ( .A1(n582), .A2(n581), .ZN(n361) );
  OR2_X1 U475 ( .A1(n556), .A2(n555), .ZN(n362) );
  XOR2_X1 U476 ( .A(n605), .B(KEYINPUT84), .Z(n363) );
  NAND2_X1 U477 ( .A1(n655), .A2(n699), .ZN(n741) );
  NAND2_X1 U478 ( .A1(n534), .A2(G214), .ZN(n719) );
  INV_X1 U479 ( .A(n719), .ZN(n396) );
  OR2_X1 U480 ( .A1(n525), .A2(G952), .ZN(n672) );
  XNOR2_X1 U481 ( .A(n366), .B(n533), .ZN(n663) );
  AND2_X1 U482 ( .A1(n370), .A2(n672), .ZN(n364) );
  AND2_X1 U483 ( .A1(n647), .A2(n417), .ZN(n365) );
  NAND2_X1 U484 ( .A1(n755), .A2(n365), .ZN(n416) );
  NOR2_X1 U485 ( .A1(n755), .A2(n417), .ZN(n379) );
  XNOR2_X2 U486 ( .A(n380), .B(KEYINPUT45), .ZN(n755) );
  NAND2_X1 U487 ( .A1(n663), .A2(n537), .ZN(n367) );
  NAND2_X1 U488 ( .A1(n360), .A2(n375), .ZN(n368) );
  NAND2_X1 U489 ( .A1(n375), .A2(n670), .ZN(n370) );
  XNOR2_X2 U490 ( .A(n376), .B(n446), .ZN(n522) );
  XNOR2_X2 U491 ( .A(n378), .B(n377), .ZN(n376) );
  XNOR2_X2 U492 ( .A(G113), .B(KEYINPUT72), .ZN(n377) );
  XNOR2_X2 U493 ( .A(G119), .B(G116), .ZN(n378) );
  NAND2_X1 U494 ( .A1(n402), .A2(n399), .ZN(n380) );
  XNOR2_X2 U495 ( .A(n592), .B(KEYINPUT102), .ZN(n690) );
  NAND2_X1 U496 ( .A1(n404), .A2(n361), .ZN(n403) );
  INV_X1 U497 ( .A(n579), .ZN(n404) );
  NOR2_X2 U498 ( .A1(n576), .A2(n578), .ZN(n577) );
  NAND2_X1 U499 ( .A1(n413), .A2(n416), .ZN(n383) );
  NOR2_X2 U500 ( .A1(n741), .A2(n656), .ZN(n659) );
  NAND2_X1 U501 ( .A1(n386), .A2(n384), .ZN(n391) );
  NAND2_X1 U502 ( .A1(n385), .A2(KEYINPUT48), .ZN(n384) );
  INV_X1 U503 ( .A(n387), .ZN(n385) );
  INV_X1 U504 ( .A(n393), .ZN(n390) );
  INV_X1 U505 ( .A(KEYINPUT48), .ZN(n392) );
  XNOR2_X1 U506 ( .A(n768), .B(n397), .ZN(n657) );
  XNOR2_X1 U507 ( .A(n398), .B(n449), .ZN(n397) );
  XNOR2_X1 U508 ( .A(n522), .B(n447), .ZN(n398) );
  NAND2_X1 U509 ( .A1(n601), .A2(KEYINPUT44), .ZN(n401) );
  NAND2_X1 U510 ( .A1(n405), .A2(n403), .ZN(n402) );
  NAND2_X1 U511 ( .A1(n406), .A2(n580), .ZN(n405) );
  XNOR2_X1 U512 ( .A(n577), .B(KEYINPUT75), .ZN(n406) );
  NAND2_X1 U513 ( .A1(n407), .A2(n604), .ZN(n605) );
  NAND2_X1 U514 ( .A1(n717), .A2(KEYINPUT47), .ZN(n407) );
  NAND2_X1 U515 ( .A1(n643), .A2(n635), .ZN(n409) );
  INV_X1 U516 ( .A(KEYINPUT86), .ZN(n417) );
  XNOR2_X2 U517 ( .A(n419), .B(KEYINPUT19), .ZN(n614) );
  NAND2_X1 U518 ( .A1(n552), .A2(n719), .ZN(n419) );
  XNOR2_X2 U519 ( .A(n421), .B(KEYINPUT77), .ZN(n587) );
  NAND2_X1 U520 ( .A1(n565), .A2(n708), .ZN(n421) );
  NAND2_X1 U521 ( .A1(n357), .A2(n435), .ZN(n434) );
  NAND2_X2 U522 ( .A1(n426), .A2(n422), .ZN(n600) );
  INV_X1 U523 ( .A(n570), .ZN(n424) );
  NOR2_X1 U524 ( .A1(n436), .A2(n433), .ZN(n425) );
  NAND2_X1 U525 ( .A1(n436), .A2(n570), .ZN(n427) );
  NAND2_X1 U526 ( .A1(n429), .A2(n570), .ZN(n428) );
  NAND2_X1 U527 ( .A1(n430), .A2(n431), .ZN(n429) );
  INV_X1 U528 ( .A(n433), .ZN(n430) );
  NAND2_X1 U529 ( .A1(n432), .A2(n435), .ZN(n431) );
  INV_X1 U530 ( .A(n726), .ZN(n432) );
  NAND2_X1 U531 ( .A1(n434), .A2(n569), .ZN(n433) );
  AND2_X1 U532 ( .A1(n588), .A2(n444), .ZN(n437) );
  OR2_X1 U533 ( .A1(n663), .A2(n441), .ZN(n440) );
  OR2_X1 U534 ( .A1(n537), .A2(n647), .ZN(n441) );
  NAND2_X1 U535 ( .A1(n537), .A2(n647), .ZN(n443) );
  XOR2_X1 U536 ( .A(KEYINPUT76), .B(KEYINPUT34), .Z(n444) );
  NOR2_X1 U537 ( .A1(n736), .A2(n735), .ZN(n445) );
  INV_X1 U538 ( .A(KEYINPUT1), .ZN(n547) );
  NOR2_X1 U539 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U540 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n446) );
  NOR2_X1 U541 ( .A1(G953), .A2(G237), .ZN(n501) );
  NAND2_X1 U542 ( .A1(n501), .A2(G210), .ZN(n447) );
  XOR2_X1 U543 ( .A(n483), .B(KEYINPUT5), .Z(n448) );
  XNOR2_X1 U544 ( .A(n448), .B(KEYINPUT78), .ZN(n449) );
  XNOR2_X1 U545 ( .A(G143), .B(G128), .ZN(n451) );
  XNOR2_X1 U546 ( .A(n451), .B(n450), .ZN(n515) );
  XNOR2_X1 U547 ( .A(KEYINPUT4), .B(G146), .ZN(n452) );
  XNOR2_X1 U548 ( .A(n515), .B(n452), .ZN(n531) );
  XNOR2_X1 U549 ( .A(n453), .B(G134), .ZN(n454) );
  XNOR2_X1 U550 ( .A(n495), .B(n454), .ZN(n455) );
  INV_X1 U551 ( .A(G902), .ZN(n519) );
  NAND2_X1 U552 ( .A1(n657), .A2(n519), .ZN(n456) );
  INV_X1 U553 ( .A(G472), .ZN(n656) );
  INV_X1 U554 ( .A(G237), .ZN(n457) );
  NAND2_X1 U555 ( .A1(n519), .A2(n457), .ZN(n534) );
  XNOR2_X2 U556 ( .A(n458), .B(G953), .ZN(n525) );
  NAND2_X1 U557 ( .A1(n525), .A2(G234), .ZN(n459) );
  XOR2_X1 U558 ( .A(KEYINPUT8), .B(n459), .Z(n511) );
  XNOR2_X1 U559 ( .A(n769), .B(G146), .ZN(n506) );
  XNOR2_X1 U560 ( .A(n461), .B(KEYINPUT94), .ZN(n463) );
  XOR2_X1 U561 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n462) );
  XNOR2_X1 U562 ( .A(n463), .B(n462), .ZN(n465) );
  XOR2_X1 U563 ( .A(n465), .B(n464), .Z(n466) );
  XOR2_X1 U564 ( .A(KEYINPUT25), .B(KEYINPUT79), .Z(n470) );
  XNOR2_X1 U565 ( .A(G902), .B(KEYINPUT15), .ZN(n603) );
  NAND2_X1 U566 ( .A1(n603), .A2(G234), .ZN(n468) );
  XNOR2_X1 U567 ( .A(n468), .B(KEYINPUT20), .ZN(n473) );
  NAND2_X1 U568 ( .A1(n473), .A2(G217), .ZN(n469) );
  XNOR2_X1 U569 ( .A(n470), .B(n469), .ZN(n471) );
  AND2_X1 U570 ( .A1(n473), .A2(G221), .ZN(n475) );
  XNOR2_X1 U571 ( .A(KEYINPUT95), .B(KEYINPUT21), .ZN(n474) );
  XNOR2_X1 U572 ( .A(n475), .B(n474), .ZN(n702) );
  INV_X1 U573 ( .A(n702), .ZN(n476) );
  NAND2_X1 U574 ( .A1(G237), .A2(G234), .ZN(n477) );
  XNOR2_X1 U575 ( .A(n477), .B(KEYINPUT14), .ZN(n479) );
  NAND2_X1 U576 ( .A1(n479), .A2(G952), .ZN(n478) );
  XNOR2_X1 U577 ( .A(n478), .B(KEYINPUT92), .ZN(n733) );
  NOR2_X1 U578 ( .A1(n733), .A2(G953), .ZN(n556) );
  NAND2_X1 U579 ( .A1(G902), .A2(n479), .ZN(n554) );
  NOR2_X1 U580 ( .A1(n525), .A2(n554), .ZN(n480) );
  XOR2_X1 U581 ( .A(KEYINPUT106), .B(n480), .Z(n481) );
  NOR2_X1 U582 ( .A1(G900), .A2(n481), .ZN(n482) );
  OR2_X1 U583 ( .A1(n556), .A2(n482), .ZN(n543) );
  NAND2_X1 U584 ( .A1(n708), .A2(n543), .ZN(n493) );
  XNOR2_X1 U585 ( .A(n483), .B(KEYINPUT74), .ZN(n486) );
  INV_X1 U586 ( .A(G104), .ZN(n484) );
  XNOR2_X1 U587 ( .A(n485), .B(n484), .ZN(n762) );
  XNOR2_X1 U588 ( .A(n486), .B(n762), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n525), .A2(G227), .ZN(n487) );
  XNOR2_X1 U590 ( .A(n487), .B(G140), .ZN(n488) );
  XNOR2_X1 U591 ( .A(n532), .B(n488), .ZN(n489) );
  NAND2_X1 U592 ( .A1(n744), .A2(n519), .ZN(n492) );
  XNOR2_X1 U593 ( .A(KEYINPUT71), .B(G469), .ZN(n490) );
  XNOR2_X1 U594 ( .A(n490), .B(KEYINPUT70), .ZN(n491) );
  BUF_X1 U595 ( .A(n548), .Z(n612) );
  NOR2_X1 U596 ( .A1(n493), .A2(n612), .ZN(n494) );
  XNOR2_X1 U597 ( .A(n496), .B(n495), .ZN(n500) );
  XNOR2_X1 U598 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U599 ( .A(n500), .B(n499), .ZN(n505) );
  XOR2_X1 U600 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n503) );
  NAND2_X1 U601 ( .A1(n501), .A2(G214), .ZN(n502) );
  XNOR2_X1 U602 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U603 ( .A(n505), .B(n504), .ZN(n507) );
  XNOR2_X1 U604 ( .A(n507), .B(n506), .ZN(n649) );
  NOR2_X1 U605 ( .A1(G902), .A2(n649), .ZN(n510) );
  XNOR2_X1 U606 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n508) );
  NAND2_X1 U607 ( .A1(n511), .A2(G217), .ZN(n518) );
  XNOR2_X1 U608 ( .A(n356), .B(G122), .ZN(n513) );
  XNOR2_X1 U609 ( .A(n514), .B(n513), .ZN(n516) );
  XNOR2_X1 U610 ( .A(n516), .B(n515), .ZN(n517) );
  NAND2_X1 U611 ( .A1(n671), .A2(n519), .ZN(n520) );
  INV_X1 U612 ( .A(G478), .ZN(n670) );
  XNOR2_X1 U613 ( .A(n520), .B(n670), .ZN(n590) );
  OR2_X1 U614 ( .A1(n558), .A2(n590), .ZN(n568) );
  XNOR2_X1 U615 ( .A(KEYINPUT16), .B(G122), .ZN(n521) );
  XOR2_X1 U616 ( .A(G125), .B(KEYINPUT90), .Z(n524) );
  XNOR2_X1 U617 ( .A(n524), .B(n523), .ZN(n529) );
  NAND2_X1 U618 ( .A1(n525), .A2(G224), .ZN(n527) );
  XNOR2_X1 U619 ( .A(KEYINPUT91), .B(KEYINPUT80), .ZN(n526) );
  XNOR2_X1 U620 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U621 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U622 ( .A(n532), .B(n531), .ZN(n533) );
  INV_X1 U623 ( .A(n603), .ZN(n647) );
  NAND2_X1 U624 ( .A1(n534), .A2(G210), .ZN(n536) );
  INV_X1 U625 ( .A(KEYINPUT82), .ZN(n535) );
  XNOR2_X1 U626 ( .A(n536), .B(n535), .ZN(n537) );
  BUF_X1 U627 ( .A(n552), .Z(n631) );
  INV_X1 U628 ( .A(n631), .ZN(n620) );
  NOR2_X1 U629 ( .A1(n568), .A2(n620), .ZN(n538) );
  NAND2_X1 U630 ( .A1(n632), .A2(n538), .ZN(n604) );
  XOR2_X1 U631 ( .A(G143), .B(KEYINPUT113), .Z(n539) );
  XNOR2_X1 U632 ( .A(n604), .B(n539), .ZN(G45) );
  AND2_X1 U633 ( .A1(n591), .A2(n590), .ZN(n687) );
  INV_X1 U634 ( .A(KEYINPUT6), .ZN(n540) );
  NOR2_X1 U635 ( .A1(n702), .A2(n542), .ZN(n609) );
  INV_X1 U636 ( .A(n543), .ZN(n606) );
  NOR2_X1 U637 ( .A1(n606), .A2(n396), .ZN(n544) );
  NAND2_X1 U638 ( .A1(n609), .A2(n544), .ZN(n545) );
  NOR2_X1 U639 ( .A1(n595), .A2(n545), .ZN(n546) );
  NAND2_X1 U640 ( .A1(n687), .A2(n546), .ZN(n621) );
  NOR2_X1 U641 ( .A1(n621), .A2(n707), .ZN(n550) );
  XNOR2_X1 U642 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n549) );
  XNOR2_X1 U643 ( .A(n550), .B(n549), .ZN(n551) );
  AND2_X1 U644 ( .A1(n551), .A2(n620), .ZN(n645) );
  XOR2_X1 U645 ( .A(G140), .B(n645), .Z(G42) );
  NOR2_X1 U646 ( .A1(n754), .A2(G898), .ZN(n553) );
  XNOR2_X1 U647 ( .A(n553), .B(KEYINPUT93), .ZN(n764) );
  NOR2_X1 U648 ( .A1(n764), .A2(n554), .ZN(n555) );
  XNOR2_X1 U649 ( .A(KEYINPUT89), .B(KEYINPUT0), .ZN(n557) );
  NAND2_X1 U650 ( .A1(n590), .A2(n558), .ZN(n722) );
  NOR2_X1 U651 ( .A1(n722), .A2(n702), .ZN(n559) );
  INV_X1 U652 ( .A(KEYINPUT22), .ZN(n560) );
  XNOR2_X2 U653 ( .A(n561), .B(n560), .ZN(n598) );
  NOR2_X1 U654 ( .A1(n542), .A2(n594), .ZN(n562) );
  AND2_X1 U655 ( .A1(n562), .A2(n595), .ZN(n563) );
  NAND2_X1 U656 ( .A1(n598), .A2(n563), .ZN(n564) );
  XNOR2_X1 U657 ( .A(n564), .B(KEYINPUT32), .ZN(n582) );
  XNOR2_X1 U658 ( .A(n582), .B(G119), .ZN(G21) );
  XNOR2_X2 U659 ( .A(n566), .B(KEYINPUT33), .ZN(n726) );
  INV_X1 U660 ( .A(n568), .ZN(n569) );
  XNOR2_X1 U661 ( .A(KEYINPUT87), .B(KEYINPUT35), .ZN(n570) );
  NAND2_X1 U662 ( .A1(n600), .A2(n582), .ZN(n576) );
  NOR2_X1 U663 ( .A1(n707), .A2(n705), .ZN(n571) );
  NAND2_X1 U664 ( .A1(n598), .A2(n571), .ZN(n573) );
  INV_X1 U665 ( .A(KEYINPUT66), .ZN(n572) );
  XNOR2_X1 U666 ( .A(n573), .B(n572), .ZN(n574) );
  INV_X1 U667 ( .A(n542), .ZN(n701) );
  NAND2_X1 U668 ( .A1(n574), .A2(n701), .ZN(n575) );
  XNOR2_X1 U669 ( .A(n575), .B(KEYINPUT105), .ZN(n578) );
  BUF_X1 U670 ( .A(n578), .Z(n579) );
  INV_X1 U671 ( .A(KEYINPUT44), .ZN(n580) );
  NOR2_X1 U672 ( .A1(n580), .A2(KEYINPUT75), .ZN(n581) );
  INV_X1 U673 ( .A(n708), .ZN(n583) );
  NOR2_X1 U674 ( .A1(n583), .A2(n612), .ZN(n584) );
  NAND2_X1 U675 ( .A1(n584), .A2(n607), .ZN(n585) );
  NOR2_X1 U676 ( .A1(n357), .A2(n585), .ZN(n586) );
  XNOR2_X1 U677 ( .A(n586), .B(KEYINPUT96), .ZN(n677) );
  AND2_X1 U678 ( .A1(n587), .A2(n705), .ZN(n712) );
  NAND2_X1 U679 ( .A1(n712), .A2(n588), .ZN(n589) );
  XNOR2_X1 U680 ( .A(n589), .B(KEYINPUT31), .ZN(n689) );
  NOR2_X1 U681 ( .A1(n677), .A2(n689), .ZN(n593) );
  INV_X1 U682 ( .A(n687), .ZN(n635) );
  NOR2_X1 U683 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U684 ( .A1(n593), .A2(n717), .ZN(n599) );
  AND2_X1 U685 ( .A1(n542), .A2(n594), .ZN(n596) );
  AND2_X1 U686 ( .A1(n596), .A2(n595), .ZN(n597) );
  AND2_X1 U687 ( .A1(n598), .A2(n597), .ZN(n674) );
  NOR2_X1 U688 ( .A1(n599), .A2(n674), .ZN(n602) );
  INV_X1 U689 ( .A(n600), .ZN(n601) );
  NOR2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U692 ( .A(KEYINPUT28), .B(n610), .ZN(n611) );
  XNOR2_X1 U693 ( .A(n611), .B(KEYINPUT108), .ZN(n613) );
  NOR2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n639) );
  BUF_X1 U695 ( .A(n614), .Z(n615) );
  NAND2_X1 U696 ( .A1(n639), .A2(n615), .ZN(n681) );
  NAND2_X1 U697 ( .A1(n681), .A2(KEYINPUT85), .ZN(n619) );
  INV_X1 U698 ( .A(KEYINPUT85), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n681), .A2(KEYINPUT47), .ZN(n616) );
  NAND2_X1 U700 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n624) );
  NOR2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U703 ( .A(n622), .B(KEYINPUT36), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n623), .A2(n707), .ZN(n694) );
  NAND2_X1 U705 ( .A1(n624), .A2(n694), .ZN(n628) );
  NOR2_X1 U706 ( .A1(n717), .A2(n681), .ZN(n625) );
  NOR2_X1 U707 ( .A1(n626), .A2(KEYINPUT47), .ZN(n627) );
  NOR2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  INV_X1 U709 ( .A(KEYINPUT38), .ZN(n630) );
  XNOR2_X1 U710 ( .A(n631), .B(n630), .ZN(n720) );
  NAND2_X1 U711 ( .A1(n632), .A2(n720), .ZN(n634) );
  INV_X1 U712 ( .A(KEYINPUT39), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n634), .B(n633), .ZN(n644) );
  NOR2_X1 U714 ( .A1(n635), .A2(n644), .ZN(n636) );
  XNOR2_X1 U715 ( .A(n636), .B(KEYINPUT40), .ZN(n779) );
  XNOR2_X1 U716 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n720), .A2(n719), .ZN(n718) );
  NOR2_X1 U718 ( .A1(n718), .A2(n722), .ZN(n638) );
  XNOR2_X1 U719 ( .A(n638), .B(n637), .ZN(n734) );
  NAND2_X1 U720 ( .A1(n639), .A2(n734), .ZN(n640) );
  XNOR2_X1 U721 ( .A(n641), .B(n640), .ZN(n778) );
  NOR2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n696) );
  NOR2_X1 U723 ( .A1(n696), .A2(n645), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n647), .A2(KEYINPUT2), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n697), .A2(KEYINPUT2), .ZN(n699) );
  NAND2_X1 U726 ( .A1(n662), .A2(G475), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n649), .B(KEYINPUT59), .ZN(n650) );
  XNOR2_X1 U728 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n652), .A2(n672), .ZN(n654) );
  XNOR2_X1 U730 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n654), .B(n653), .ZN(G60) );
  XOR2_X1 U732 ( .A(KEYINPUT62), .B(n657), .Z(n658) );
  XNOR2_X1 U733 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U734 ( .A1(n660), .A2(n672), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n661), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U736 ( .A1(n662), .A2(G210), .ZN(n666) );
  XNOR2_X1 U737 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n663), .B(n664), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U740 ( .A1(n667), .A2(n672), .ZN(n669) );
  XNOR2_X1 U741 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n669), .B(n668), .ZN(G51) );
  INV_X1 U743 ( .A(n672), .ZN(n753) );
  XNOR2_X1 U744 ( .A(G110), .B(KEYINPUT111), .ZN(n673) );
  XNOR2_X1 U745 ( .A(n579), .B(n673), .ZN(G12) );
  XNOR2_X1 U746 ( .A(n600), .B(G122), .ZN(G24) );
  XOR2_X1 U747 ( .A(G101), .B(n674), .Z(G3) );
  NAND2_X1 U748 ( .A1(n677), .A2(n687), .ZN(n675) );
  XNOR2_X1 U749 ( .A(n675), .B(KEYINPUT110), .ZN(n676) );
  XNOR2_X1 U750 ( .A(G104), .B(n676), .ZN(G6) );
  XOR2_X1 U751 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n679) );
  NAND2_X1 U752 ( .A1(n677), .A2(n690), .ZN(n678) );
  XNOR2_X1 U753 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U754 ( .A(G107), .B(n680), .ZN(G9) );
  XOR2_X1 U755 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n683) );
  INV_X1 U756 ( .A(n681), .ZN(n685) );
  NAND2_X1 U757 ( .A1(n685), .A2(n690), .ZN(n682) );
  XNOR2_X1 U758 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U759 ( .A(G128), .B(n684), .ZN(G30) );
  NAND2_X1 U760 ( .A1(n685), .A2(n687), .ZN(n686) );
  XNOR2_X1 U761 ( .A(n686), .B(G146), .ZN(G48) );
  NAND2_X1 U762 ( .A1(n689), .A2(n687), .ZN(n688) );
  XNOR2_X1 U763 ( .A(n688), .B(G113), .ZN(G15) );
  NAND2_X1 U764 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U765 ( .A(n691), .B(KEYINPUT114), .ZN(n692) );
  XNOR2_X1 U766 ( .A(n356), .B(n692), .ZN(G18) );
  XNOR2_X1 U767 ( .A(KEYINPUT115), .B(KEYINPUT37), .ZN(n693) );
  XNOR2_X1 U768 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U769 ( .A(G125), .B(n695), .ZN(G27) );
  XOR2_X1 U770 ( .A(G134), .B(n696), .Z(G36) );
  NOR2_X1 U771 ( .A1(n697), .A2(KEYINPUT2), .ZN(n698) );
  XNOR2_X1 U772 ( .A(n698), .B(KEYINPUT83), .ZN(n700) );
  AND2_X1 U773 ( .A1(n700), .A2(n699), .ZN(n738) );
  XNOR2_X1 U774 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n715) );
  NAND2_X1 U775 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U776 ( .A(KEYINPUT49), .B(n703), .ZN(n704) );
  NOR2_X1 U777 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U778 ( .A(KEYINPUT116), .B(n706), .Z(n711) );
  NOR2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U780 ( .A(n709), .B(KEYINPUT50), .ZN(n710) );
  NOR2_X1 U781 ( .A1(n711), .A2(n710), .ZN(n713) );
  NOR2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U783 ( .A(n715), .B(n714), .Z(n716) );
  NAND2_X1 U784 ( .A1(n734), .A2(n716), .ZN(n729) );
  OR2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n725) );
  NOR2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U787 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U788 ( .A(KEYINPUT118), .B(n723), .Z(n724) );
  NAND2_X1 U789 ( .A1(n725), .A2(n724), .ZN(n727) );
  NAND2_X1 U790 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U791 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U792 ( .A(n730), .B(KEYINPUT119), .ZN(n731) );
  XNOR2_X1 U793 ( .A(KEYINPUT52), .B(n731), .ZN(n732) );
  NOR2_X1 U794 ( .A1(n733), .A2(n732), .ZN(n736) );
  AND2_X1 U795 ( .A1(n726), .A2(n734), .ZN(n735) );
  XNOR2_X1 U796 ( .A(KEYINPUT53), .B(KEYINPUT120), .ZN(n739) );
  XNOR2_X1 U797 ( .A(n740), .B(n739), .ZN(G75) );
  NAND2_X1 U798 ( .A1(n748), .A2(G469), .ZN(n746) );
  XOR2_X1 U799 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n742) );
  XOR2_X1 U800 ( .A(n742), .B(KEYINPUT122), .Z(n743) );
  XNOR2_X1 U801 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U802 ( .A1(n753), .A2(n747), .ZN(G54) );
  NAND2_X1 U803 ( .A1(n748), .A2(G217), .ZN(n751) );
  XNOR2_X1 U804 ( .A(n751), .B(n750), .ZN(n752) );
  NOR2_X1 U805 ( .A1(n753), .A2(n752), .ZN(G66) );
  NAND2_X1 U806 ( .A1(n755), .A2(n754), .ZN(n759) );
  NAND2_X1 U807 ( .A1(G953), .A2(G224), .ZN(n756) );
  XNOR2_X1 U808 ( .A(KEYINPUT61), .B(n756), .ZN(n757) );
  NAND2_X1 U809 ( .A1(n757), .A2(G898), .ZN(n758) );
  NAND2_X1 U810 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U811 ( .A(n760), .B(KEYINPUT126), .ZN(n767) );
  XOR2_X1 U812 ( .A(G101), .B(n762), .Z(n763) );
  XNOR2_X1 U813 ( .A(n359), .B(n763), .ZN(n765) );
  NAND2_X1 U814 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U815 ( .A(n767), .B(n766), .Z(G69) );
  XOR2_X1 U816 ( .A(n769), .B(n768), .Z(n772) );
  XNOR2_X1 U817 ( .A(n770), .B(n772), .ZN(n771) );
  NAND2_X1 U818 ( .A1(n771), .A2(n525), .ZN(n777) );
  XOR2_X1 U819 ( .A(n772), .B(G227), .Z(n773) );
  NAND2_X1 U820 ( .A1(n773), .A2(G900), .ZN(n774) );
  XOR2_X1 U821 ( .A(KEYINPUT127), .B(n774), .Z(n775) );
  NAND2_X1 U822 ( .A1(n775), .A2(G953), .ZN(n776) );
  NAND2_X1 U823 ( .A1(n777), .A2(n776), .ZN(G72) );
  XOR2_X1 U824 ( .A(n778), .B(G137), .Z(G39) );
  XOR2_X1 U825 ( .A(G131), .B(n779), .Z(G33) );
endmodule

