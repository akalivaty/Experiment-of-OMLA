//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT15), .ZN(new_n206));
  INV_X1    g005(.A(G43gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G50gat), .ZN(new_n208));
  INV_X1    g007(.A(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G43gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n205), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NOR3_X1   g011(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(KEYINPUT78), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(new_n203), .A3(new_n204), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT78), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n211), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(KEYINPUT76), .A2(G43gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT76), .A2(G43gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n209), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT77), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n207), .A2(G50gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n225), .B(new_n209), .C1(new_n220), .C2(new_n221), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n219), .B1(new_n206), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n210), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT75), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n216), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n213), .A2(KEYINPUT75), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(new_n212), .ZN(new_n233));
  INV_X1    g032(.A(new_n205), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n229), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n202), .B1(new_n228), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n234), .ZN(new_n237));
  INV_X1    g036(.A(new_n229), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n222), .A2(KEYINPUT77), .B1(new_n207), .B2(G50gat), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT15), .B1(new_n240), .B2(new_n226), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n239), .B(KEYINPUT79), .C1(new_n241), .C2(new_n219), .ZN(new_n242));
  XNOR2_X1  g041(.A(G15gat), .B(G22gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT16), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(G1gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(G1gat), .B2(new_n243), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(G8gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n236), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n236), .A2(KEYINPUT81), .A3(new_n242), .A4(new_n247), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G229gat), .A2(G233gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n242), .A3(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n246), .B(G8gat), .Z(new_n257));
  OAI211_X1 g056(.A(new_n239), .B(KEYINPUT17), .C1(new_n241), .C2(new_n219), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n252), .A2(new_n253), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT18), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n252), .A2(KEYINPUT18), .A3(new_n253), .A4(new_n259), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G113gat), .B(G141gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT74), .B(KEYINPUT11), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G169gat), .B(G197gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT12), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n236), .A2(new_n242), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n257), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n253), .B(KEYINPUT13), .Z(new_n275));
  AOI21_X1  g074(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n275), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n262), .A2(new_n277), .A3(new_n263), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n264), .A2(new_n276), .B1(new_n278), .B2(new_n271), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n280));
  NOR2_X1   g079(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT64), .B(G183gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(new_n282), .B2(KEYINPUT27), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n280), .B1(new_n283), .B2(G190gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT27), .B(G183gat), .ZN(new_n285));
  INV_X1    g084(.A(G190gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT28), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT26), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT26), .ZN(new_n292));
  INV_X1    g091(.A(G169gat), .ZN(new_n293));
  INV_X1    g092(.A(G176gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n289), .B(new_n291), .C1(new_n295), .C2(new_n290), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n290), .A2(KEYINPUT23), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n298), .B(new_n300), .C1(new_n293), .C2(new_n294), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n289), .A2(KEYINPUT24), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n282), .B2(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(new_n304), .B2(new_n306), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n302), .B1(new_n301), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n297), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G113gat), .B(G120gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(KEYINPUT1), .ZN(new_n317));
  XNOR2_X1  g116(.A(G127gat), .B(G134gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n317), .B(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n288), .A2(new_n296), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n320), .A3(new_n313), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(KEYINPUT65), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT34), .ZN(new_n325));
  NAND2_X1  g124(.A1(G227gat), .A2(G233gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT65), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n315), .A2(new_n327), .A3(new_n320), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n324), .A2(new_n325), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(KEYINPUT65), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(new_n313), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n317), .B(new_n318), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n326), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT34), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G15gat), .B(G43gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G71gat), .B(G99gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n334), .A2(new_n335), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT33), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(KEYINPUT32), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT33), .B1(new_n334), .B2(new_n335), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n329), .B(new_n336), .C1(new_n347), .C2(new_n340), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n344), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(G141gat), .B(G148gat), .Z(new_n350));
  INV_X1    g149(.A(G155gat), .ZN(new_n351));
  INV_X1    g150(.A(G162gat), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT2), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(G155gat), .B(G162gat), .Z(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n354), .B(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G211gat), .B(G218gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT66), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n360));
  INV_X1    g159(.A(G197gat), .ZN(new_n361));
  INV_X1    g160(.A(G204gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n360), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n359), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n357), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G228gat), .A2(G233gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n357), .A2(new_n369), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n366), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  OR3_X1    g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G22gat), .ZN(new_n375));
  INV_X1    g174(.A(G228gat), .ZN(new_n376));
  INV_X1    g175(.A(G233gat), .ZN(new_n377));
  OAI22_X1  g176(.A1(new_n370), .A2(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT70), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(G78gat), .B(G106gat), .Z(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT31), .B(G50gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n374), .A2(new_n378), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G22gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n379), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n387), .A2(KEYINPUT70), .A3(new_n379), .A4(new_n384), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n346), .B1(new_n344), .B2(new_n348), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n349), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n394), .B(new_n395), .Z(new_n396));
  AOI22_X1  g195(.A1(new_n331), .A2(new_n367), .B1(G226gat), .B2(G233gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n315), .A2(new_n398), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n397), .A2(new_n366), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n366), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n331), .A2(G226gat), .A3(G233gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n398), .B1(new_n315), .B2(KEYINPUT29), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(KEYINPUT30), .B(new_n396), .C1(new_n400), .C2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n366), .B1(new_n397), .B2(new_n399), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n403), .A3(new_n401), .ZN(new_n407));
  INV_X1    g206(.A(new_n396), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT67), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n396), .B1(new_n400), .B2(new_n404), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n408), .B1(new_n406), .B2(new_n407), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n415), .A2(KEYINPUT67), .A3(KEYINPUT30), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n410), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n357), .A2(new_n320), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT4), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n354), .B(new_n355), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT3), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n372), .A2(new_n421), .A3(new_n332), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n423), .B(KEYINPUT68), .Z(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n419), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n332), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n418), .A2(new_n427), .A3(KEYINPUT69), .ZN(new_n428));
  OR3_X1    g227(.A1(new_n357), .A2(new_n320), .A3(KEYINPUT69), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n424), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT5), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n419), .A2(new_n422), .A3(KEYINPUT5), .A4(new_n425), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT71), .ZN(new_n435));
  XNOR2_X1  g234(.A(G1gat), .B(G29gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT0), .ZN(new_n437));
  XNOR2_X1  g236(.A(G57gat), .B(G85gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT71), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n432), .A2(new_n441), .A3(new_n433), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n435), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT6), .B1(new_n434), .B2(new_n439), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n434), .A2(new_n439), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n443), .A2(new_n444), .B1(KEYINPUT6), .B2(new_n445), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n417), .A2(new_n446), .A3(KEYINPUT35), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n393), .A2(new_n447), .A3(KEYINPUT73), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT73), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n344), .A2(new_n348), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n345), .ZN(new_n451));
  INV_X1    g250(.A(new_n390), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n381), .A2(new_n384), .B1(new_n387), .B2(new_n379), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n344), .A2(new_n346), .A3(new_n348), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n443), .A2(new_n444), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n445), .A2(KEYINPUT6), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n405), .A2(new_n409), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT67), .B1(new_n415), .B2(KEYINPUT30), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n412), .A2(new_n411), .A3(new_n413), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT35), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n459), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n449), .B1(new_n456), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n444), .B1(new_n439), .B2(new_n434), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n458), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT35), .B1(new_n456), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n448), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT72), .B1(new_n400), .B2(new_n404), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT37), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT72), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n406), .B2(new_n407), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n477), .A3(new_n408), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT38), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n473), .A2(new_n477), .A3(new_n480), .A4(new_n408), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n479), .A2(new_n446), .A3(new_n481), .A4(new_n412), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n419), .A2(new_n422), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n424), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n428), .A2(new_n429), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n484), .B(KEYINPUT39), .C1(new_n424), .C2(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(new_n439), .C1(KEYINPUT39), .C2(new_n484), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT40), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(new_n443), .A3(new_n417), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n482), .A2(new_n489), .A3(new_n454), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(new_n349), .B2(new_n392), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n451), .A2(KEYINPUT36), .A3(new_n455), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n469), .A2(new_n391), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n490), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n279), .B1(new_n471), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT21), .ZN(new_n498));
  NAND2_X1  g297(.A1(G71gat), .A2(G78gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT9), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT83), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(KEYINPUT83), .A3(new_n500), .ZN(new_n504));
  INV_X1    g303(.A(G57gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(G64gat), .ZN(new_n506));
  INV_X1    g305(.A(G64gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(G57gat), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n503), .B(new_n504), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(G71gat), .A2(G78gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT82), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n499), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n512), .B1(new_n511), .B2(new_n510), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(new_n505), .B2(G64gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n507), .A2(KEYINPUT84), .A3(G57gat), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n516), .B(new_n517), .C1(G57gat), .C2(new_n507), .ZN(new_n518));
  INV_X1    g317(.A(new_n499), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(new_n510), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n518), .A2(new_n521), .A3(new_n504), .A4(new_n503), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n257), .B1(new_n498), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT85), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(new_n351), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n525), .B(new_n527), .Z(new_n528));
  NAND2_X1  g327(.A1(new_n523), .A2(new_n498), .ZN(new_n529));
  NAND2_X1  g328(.A1(G231gat), .A2(G233gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G127gat), .ZN(new_n532));
  XOR2_X1   g331(.A(G183gat), .B(G211gat), .Z(new_n533));
  OR2_X1    g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n528), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n525), .B(new_n527), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT88), .ZN(new_n541));
  XNOR2_X1  g340(.A(G190gat), .B(G218gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT41), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT87), .ZN(new_n546));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g347(.A1(G85gat), .A2(G92gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  INV_X1    g351(.A(G92gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n548), .A2(new_n551), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G99gat), .B(G106gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n546), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n551), .A2(new_n555), .ZN(new_n560));
  AOI22_X1  g359(.A1(KEYINPUT8), .A2(new_n547), .B1(new_n552), .B2(new_n553), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n560), .A2(KEYINPUT87), .A3(new_n557), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n556), .A2(new_n558), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n545), .B1(new_n272), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n256), .A2(new_n258), .A3(new_n565), .ZN(new_n568));
  AOI211_X1 g367(.A(new_n541), .B(new_n543), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n568), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n542), .B1(new_n571), .B2(new_n566), .ZN(new_n572));
  INV_X1    g371(.A(new_n272), .ZN(new_n573));
  INV_X1    g372(.A(new_n565), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n575), .A2(new_n568), .A3(new_n545), .A4(new_n543), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(new_n541), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT86), .B(G134gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(new_n352), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n544), .A2(KEYINPUT41), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n582), .B1(new_n576), .B2(KEYINPUT89), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n570), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n570), .B2(new_n577), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n540), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n558), .A2(KEYINPUT90), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT90), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n557), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n556), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n563), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n503), .A2(new_n504), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(new_n520), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n594), .A2(new_n518), .B1(new_n509), .B2(new_n513), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n523), .A2(new_n563), .A3(new_n564), .ZN(new_n597));
  AND4_X1   g396(.A1(G230gat), .A2(new_n596), .A3(G233gat), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT10), .B1(new_n596), .B2(new_n597), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT10), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n565), .A2(new_n523), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n604), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n605), .A2(new_n607), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n604), .B(KEYINPUT92), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n598), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n601), .B(KEYINPUT91), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n609), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n497), .A2(new_n587), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n468), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT93), .B(G1gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(G1324gat));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n417), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(G8gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT42), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT16), .B(G8gat), .Z(new_n626));
  NAND3_X1  g425(.A1(new_n618), .A2(new_n417), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n627), .A2(KEYINPUT94), .A3(new_n625), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT94), .B1(new_n627), .B2(new_n625), .ZN(new_n629));
  OAI221_X1 g428(.A(new_n624), .B1(new_n625), .B2(new_n627), .C1(new_n628), .C2(new_n629), .ZN(G1325gat));
  INV_X1    g429(.A(G15gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n451), .A2(new_n455), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n494), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n618), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n636), .B2(new_n631), .ZN(G1326gat));
  NAND2_X1  g436(.A1(new_n618), .A2(new_n391), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT95), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT95), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n618), .A2(new_n640), .A3(new_n391), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT43), .B(G22gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n642), .B(new_n644), .ZN(G1327gat));
  NAND2_X1  g444(.A1(new_n471), .A2(new_n496), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n586), .ZN(new_n647));
  INV_X1    g446(.A(new_n540), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(new_n616), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n278), .A2(new_n271), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n276), .A2(new_n262), .A3(new_n263), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(new_n203), .A3(new_n619), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT45), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n653), .ZN(new_n659));
  INV_X1    g458(.A(new_n586), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(new_n471), .B2(new_n496), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT44), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n658), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(G29gat), .B1(new_n663), .B2(new_n468), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n656), .A2(new_n664), .ZN(G1328gat));
  NAND3_X1  g464(.A1(new_n654), .A2(new_n204), .A3(new_n417), .ZN(new_n666));
  AND2_X1   g465(.A1(KEYINPUT96), .A2(KEYINPUT46), .ZN(new_n667));
  NOR2_X1   g466(.A1(KEYINPUT96), .A2(KEYINPUT46), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(G36gat), .B1(new_n663), .B2(new_n463), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n669), .B(new_n670), .C1(new_n667), .C2(new_n666), .ZN(G1329gat));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n633), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n220), .A2(new_n221), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n494), .A2(new_n673), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n663), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT47), .ZN(G1330gat));
  AND4_X1   g476(.A1(new_n209), .A2(new_n649), .A3(new_n391), .A4(new_n586), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n497), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT98), .Z(new_n680));
  NAND4_X1  g479(.A1(new_n658), .A2(new_n391), .A3(new_n659), .A4(new_n662), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G50gat), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT48), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT97), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n680), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(KEYINPUT97), .A3(G50gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n682), .A2(new_n679), .A3(new_n684), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n685), .A2(new_n686), .B1(KEYINPUT48), .B2(new_n687), .ZN(G1331gat));
  NAND2_X1  g487(.A1(new_n651), .A2(new_n616), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n587), .A2(new_n650), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n471), .B2(new_n496), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n619), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT100), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT99), .B(G57gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1332gat));
  AOI21_X1  g495(.A(new_n463), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT101), .Z(new_n698));
  NAND2_X1  g497(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT102), .Z(new_n700));
  NOR2_X1   g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1333gat));
  NAND3_X1  g501(.A1(new_n692), .A2(G71gat), .A3(new_n635), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n633), .A2(KEYINPUT103), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n632), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n692), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n703), .B1(new_n708), .B2(G71gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g509(.A1(new_n692), .A2(new_n391), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g511(.A1(new_n468), .A2(G85gat), .A3(new_n617), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n648), .A2(new_n652), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  AOI211_X1 g515(.A(new_n660), .B(new_n716), .C1(new_n471), .C2(new_n496), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT51), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n646), .A2(new_n586), .A3(new_n715), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT105), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT104), .B1(new_n720), .B2(new_n721), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n717), .A2(new_n725), .A3(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n714), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n716), .A2(new_n617), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n658), .A2(new_n619), .A3(new_n662), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G85gat), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT106), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n724), .A2(new_n726), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n718), .B1(new_n717), .B2(KEYINPUT51), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n720), .A2(KEYINPUT105), .A3(new_n721), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n713), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n739), .A3(new_n731), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n733), .A2(new_n740), .ZN(G1336gat));
  NAND3_X1  g540(.A1(new_n417), .A2(new_n553), .A3(new_n616), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT51), .B1(new_n720), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n743), .B2(new_n720), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n742), .B1(new_n745), .B2(new_n727), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n658), .A2(new_n417), .A3(new_n662), .A4(new_n729), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(G92gat), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT52), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT52), .B1(new_n747), .B2(G92gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n737), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n742), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(G1337gat));
  XOR2_X1   g552(.A(KEYINPUT108), .B(G99gat), .Z(new_n754));
  NAND3_X1  g553(.A1(new_n658), .A2(new_n662), .A3(new_n729), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(new_n494), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n632), .A2(new_n617), .A3(new_n754), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n751), .B2(new_n757), .ZN(G1338gat));
  OR3_X1    g557(.A1(new_n454), .A2(G106gat), .A3(new_n617), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n745), .B2(new_n727), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n658), .A2(new_n391), .A3(new_n662), .A4(new_n729), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(G106gat), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT53), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT53), .B1(new_n761), .B2(G106gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n751), .B2(new_n759), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1339gat));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767));
  INV_X1    g566(.A(new_n269), .ZN(new_n768));
  INV_X1    g567(.A(new_n275), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n252), .A2(new_n273), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n252), .A2(new_n259), .ZN(new_n771));
  INV_X1    g570(.A(new_n253), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n770), .A2(KEYINPUT110), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n252), .A2(new_n774), .A3(new_n273), .A4(new_n769), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n768), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n767), .B1(new_n689), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n770), .A2(KEYINPUT110), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n771), .A2(new_n772), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n269), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n781), .A2(KEYINPUT111), .A3(new_n651), .A4(new_n616), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT54), .B(new_n608), .C1(new_n610), .C2(new_n612), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n784), .B(new_n612), .C1(new_n605), .C2(new_n607), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n785), .A2(KEYINPUT109), .A3(new_n602), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT109), .B1(new_n785), .B2(new_n602), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(KEYINPUT55), .B(new_n783), .C1(new_n786), .C2(new_n787), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n609), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n777), .B(new_n782), .C1(new_n279), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n660), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n790), .A2(new_n609), .A3(new_n791), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n586), .A2(new_n795), .A3(new_n651), .A4(new_n781), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n540), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n587), .A2(new_n279), .A3(new_n617), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n391), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n632), .A2(new_n468), .A3(new_n417), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(G113gat), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n803), .A2(new_n804), .A3(new_n279), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n468), .B1(new_n798), .B2(new_n799), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n393), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(KEYINPUT112), .A3(new_n393), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n417), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n652), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n805), .B1(new_n812), .B2(new_n804), .ZN(G1340gat));
  NOR2_X1   g612(.A1(new_n617), .A2(G120gat), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT113), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G120gat), .B1(new_n803), .B2(new_n617), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1341gat));
  INV_X1    g617(.A(G127gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n648), .A2(new_n819), .ZN(new_n820));
  AOI211_X1 g619(.A(new_n417), .B(new_n820), .C1(new_n809), .C2(new_n810), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n819), .B1(new_n802), .B2(new_n648), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n821), .B2(new_n824), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1342gat));
  NAND2_X1  g627(.A1(new_n586), .A2(new_n463), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT115), .ZN(new_n830));
  AOI211_X1 g629(.A(G134gat), .B(new_n830), .C1(new_n809), .C2(new_n810), .ZN(new_n831));
  XOR2_X1   g630(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n832));
  NAND2_X1  g631(.A1(new_n802), .A2(new_n586), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n831), .A2(new_n832), .B1(G134gat), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n831), .B2(new_n832), .ZN(G1343gat));
  AOI211_X1 g634(.A(new_n468), .B(new_n417), .C1(new_n492), .C2(new_n493), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n454), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n583), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n576), .A2(new_n541), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n543), .B1(new_n567), .B2(new_n568), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n840), .B1(new_n843), .B2(new_n569), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n570), .A2(new_n577), .A3(new_n583), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n844), .A2(new_n781), .A3(new_n845), .A4(new_n651), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n792), .ZN(new_n847));
  OAI22_X1  g646(.A1(new_n279), .A2(new_n792), .B1(new_n689), .B2(new_n776), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n660), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n540), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n839), .B1(new_n853), .B2(new_n799), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n847), .B1(new_n793), .B2(new_n660), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n799), .B1(new_n855), .B2(new_n648), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n856), .B2(new_n391), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n836), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G141gat), .B1(new_n858), .B2(new_n279), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT119), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n635), .A2(new_n454), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT118), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(KEYINPUT118), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n806), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n417), .ZN(new_n865));
  INV_X1    g664(.A(G141gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n866), .A3(new_n652), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n859), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n860), .A2(new_n868), .A3(KEYINPUT58), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n859), .B(new_n867), .C1(KEYINPUT119), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1344gat));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n873), .B(G148gat), .C1(new_n858), .C2(new_n617), .ZN(new_n874));
  INV_X1    g673(.A(G148gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n836), .A2(new_n616), .ZN(new_n876));
  NOR4_X1   g675(.A1(new_n540), .A2(new_n586), .A3(new_n652), .A4(new_n616), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n795), .A2(new_n652), .B1(new_n690), .B2(new_n781), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n796), .B1(new_n878), .B2(new_n586), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n879), .B2(new_n540), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n837), .B1(new_n880), .B2(new_n454), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n856), .A2(new_n838), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n876), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n875), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n648), .B1(new_n849), .B2(new_n796), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n391), .B1(new_n886), .B2(new_n877), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n837), .A2(new_n887), .B1(new_n856), .B2(new_n838), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT120), .B1(new_n888), .B2(new_n876), .ZN(new_n889));
  AOI211_X1 g688(.A(KEYINPUT121), .B(new_n873), .C1(new_n885), .C2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  INV_X1    g690(.A(new_n876), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n839), .B1(new_n798), .B2(new_n799), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n847), .B1(new_n660), .B2(new_n848), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n799), .B1(new_n894), .B2(new_n648), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n895), .B2(new_n391), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n884), .B(new_n892), .C1(new_n893), .C2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n889), .A2(G148gat), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n891), .B1(new_n898), .B2(KEYINPUT59), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n874), .B1(new_n890), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n865), .A2(new_n875), .A3(new_n616), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1345gat));
  OAI21_X1  g701(.A(G155gat), .B1(new_n858), .B2(new_n540), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n865), .A2(new_n351), .A3(new_n648), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1346gat));
  OAI21_X1  g704(.A(G162gat), .B1(new_n858), .B2(new_n660), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n830), .A2(G162gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n864), .B2(new_n907), .ZN(G1347gat));
  AOI21_X1  g707(.A(new_n619), .B1(new_n798), .B2(new_n799), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(new_n417), .A3(new_n393), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n293), .A3(new_n652), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n619), .A2(new_n463), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n707), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n800), .A2(new_n652), .A3(new_n913), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n914), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT122), .B1(new_n914), .B2(G169gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n917), .B(new_n918), .ZN(G1348gat));
  AND2_X1   g718(.A1(new_n800), .A2(new_n913), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G176gat), .B1(new_n921), .B2(new_n617), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n910), .A2(new_n294), .A3(new_n616), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1349gat));
  OAI21_X1  g723(.A(new_n282), .B1(new_n921), .B2(new_n540), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n285), .A3(new_n648), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n286), .A3(new_n586), .ZN(new_n929));
  OAI21_X1  g728(.A(G190gat), .B1(new_n921), .B2(new_n660), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1351gat));
  NAND3_X1  g732(.A1(new_n909), .A2(new_n417), .A3(new_n861), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n361), .A3(new_n652), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n494), .A2(new_n912), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n881), .A2(new_n882), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n888), .A2(KEYINPUT124), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n937), .B1(new_n943), .B2(new_n279), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G197gat), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n943), .A2(new_n937), .A3(new_n279), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n936), .B1(new_n945), .B2(new_n946), .ZN(G1352gat));
  NAND3_X1  g746(.A1(new_n935), .A2(new_n362), .A3(new_n616), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(KEYINPUT62), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(KEYINPUT126), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(G204gat), .B1(new_n943), .B2(new_n617), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT62), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G1353gat));
  INV_X1    g754(.A(G211gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n935), .A2(new_n956), .A3(new_n648), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n888), .A2(new_n540), .A3(new_n938), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n958), .A2(KEYINPUT127), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(KEYINPUT127), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n959), .A2(KEYINPUT63), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n957), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  AOI21_X1  g762(.A(G218gat), .B1(new_n935), .B2(new_n586), .ZN(new_n964));
  INV_X1    g763(.A(new_n943), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n586), .A2(G218gat), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(G1355gat));
endmodule


