

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590;

  XNOR2_X1 U322 ( .A(n451), .B(n450), .ZN(n543) );
  XNOR2_X1 U323 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n408) );
  XNOR2_X1 U324 ( .A(n468), .B(n467), .ZN(n491) );
  XNOR2_X1 U325 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U326 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n362) );
  XNOR2_X1 U327 ( .A(n363), .B(n362), .ZN(n399) );
  NOR2_X1 U328 ( .A1(n553), .A2(n481), .ZN(n465) );
  XNOR2_X1 U329 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U330 ( .A(n411), .B(G218GAT), .ZN(n415) );
  XNOR2_X1 U331 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U332 ( .A(n415), .B(n441), .ZN(n416) );
  XNOR2_X1 U333 ( .A(n409), .B(n408), .ZN(n544) );
  INV_X1 U334 ( .A(n533), .ZN(n469) );
  XNOR2_X1 U335 ( .A(n477), .B(KEYINPUT41), .ZN(n533) );
  XNOR2_X1 U336 ( .A(n423), .B(n422), .ZN(n449) );
  XNOR2_X1 U337 ( .A(n446), .B(KEYINPUT58), .ZN(n447) );
  XNOR2_X1 U338 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n290) );
  XNOR2_X1 U340 ( .A(n290), .B(KEYINPUT88), .ZN(n291) );
  XOR2_X1 U341 ( .A(n291), .B(KEYINPUT89), .Z(n293) );
  XNOR2_X1 U342 ( .A(G141GAT), .B(KEYINPUT87), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n327) );
  XOR2_X1 U344 ( .A(G120GAT), .B(KEYINPUT83), .Z(n295) );
  XNOR2_X1 U345 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n433) );
  XOR2_X1 U347 ( .A(G85GAT), .B(n433), .Z(n297) );
  XOR2_X1 U348 ( .A(G113GAT), .B(G1GAT), .Z(n330) );
  XNOR2_X1 U349 ( .A(G29GAT), .B(n330), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n327), .B(n298), .ZN(n311) );
  XOR2_X1 U352 ( .A(G155GAT), .B(G148GAT), .Z(n300) );
  XNOR2_X1 U353 ( .A(G127GAT), .B(G162GAT), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U355 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n302) );
  XNOR2_X1 U356 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U358 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U359 ( .A(KEYINPUT6), .B(G57GAT), .Z(n306) );
  NAND2_X1 U360 ( .A1(G225GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U362 ( .A(KEYINPUT92), .B(n307), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n521) );
  INV_X1 U365 ( .A(n521), .ZN(n570) );
  XOR2_X1 U366 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n313) );
  NAND2_X1 U367 ( .A1(G228GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U369 ( .A(n314), .B(G78GAT), .Z(n319) );
  XOR2_X1 U370 ( .A(G162GAT), .B(KEYINPUT77), .Z(n316) );
  XNOR2_X1 U371 ( .A(G50GAT), .B(G218GAT), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n384) );
  XNOR2_X1 U373 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n317), .B(G148GAT), .ZN(n353) );
  XNOR2_X1 U375 ( .A(n384), .B(n353), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U377 ( .A(G204GAT), .B(G211GAT), .Z(n321) );
  XNOR2_X1 U378 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U380 ( .A(n323), .B(n322), .Z(n325) );
  XOR2_X1 U381 ( .A(G22GAT), .B(G155GAT), .Z(n376) );
  XOR2_X1 U382 ( .A(G197GAT), .B(KEYINPUT21), .Z(n410) );
  XNOR2_X1 U383 ( .A(n376), .B(n410), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n456) );
  AND2_X1 U386 ( .A1(n570), .A2(n456), .ZN(n425) );
  XOR2_X1 U387 ( .A(G29GAT), .B(G43GAT), .Z(n329) );
  XNOR2_X1 U388 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n329), .B(n328), .ZN(n385) );
  XOR2_X1 U390 ( .A(n385), .B(n330), .Z(n332) );
  NAND2_X1 U391 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U393 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n334) );
  XNOR2_X1 U394 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U396 ( .A(n336), .B(n335), .Z(n344) );
  XOR2_X1 U397 ( .A(G15GAT), .B(G50GAT), .Z(n338) );
  XNOR2_X1 U398 ( .A(G169GAT), .B(G36GAT), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U400 ( .A(G8GAT), .B(G197GAT), .Z(n340) );
  XNOR2_X1 U401 ( .A(G141GAT), .B(G22GAT), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n574) );
  XOR2_X1 U405 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n346) );
  XNOR2_X1 U406 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n361) );
  XOR2_X1 U408 ( .A(KEYINPUT13), .B(G57GAT), .Z(n348) );
  XNOR2_X1 U409 ( .A(G71GAT), .B(G78GAT), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n369) );
  XOR2_X1 U411 ( .A(G99GAT), .B(G85GAT), .Z(n392) );
  XOR2_X1 U412 ( .A(n369), .B(n392), .Z(n350) );
  NAND2_X1 U413 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n359) );
  XOR2_X1 U415 ( .A(G64GAT), .B(G92GAT), .Z(n352) );
  XNOR2_X1 U416 ( .A(G176GAT), .B(G204GAT), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n419) );
  XNOR2_X1 U418 ( .A(n353), .B(n419), .ZN(n357) );
  XOR2_X1 U419 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n355) );
  XNOR2_X1 U420 ( .A(KEYINPUT71), .B(KEYINPUT74), .ZN(n354) );
  XOR2_X1 U421 ( .A(n355), .B(n354), .Z(n356) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n477) );
  NOR2_X1 U423 ( .A1(n574), .A2(n533), .ZN(n363) );
  XOR2_X1 U424 ( .A(KEYINPUT15), .B(KEYINPUT82), .Z(n365) );
  NAND2_X1 U425 ( .A1(G231GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U427 ( .A(n366), .B(KEYINPUT81), .Z(n371) );
  XOR2_X1 U428 ( .A(KEYINPUT80), .B(G211GAT), .Z(n368) );
  XNOR2_X1 U429 ( .A(G8GAT), .B(G183GAT), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n418) );
  XNOR2_X1 U431 ( .A(n369), .B(n418), .ZN(n370) );
  XNOR2_X1 U432 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U433 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n373) );
  XNOR2_X1 U434 ( .A(G1GAT), .B(G64GAT), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U436 ( .A(n375), .B(n374), .Z(n378) );
  XOR2_X1 U437 ( .A(G15GAT), .B(G127GAT), .Z(n430) );
  XNOR2_X1 U438 ( .A(n430), .B(n376), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n553) );
  XOR2_X1 U440 ( .A(KEYINPUT113), .B(n553), .Z(n566) );
  XOR2_X1 U441 ( .A(G92GAT), .B(KEYINPUT79), .Z(n380) );
  XNOR2_X1 U442 ( .A(G134GAT), .B(G106GAT), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n396) );
  XOR2_X1 U444 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n382) );
  NAND2_X1 U445 ( .A1(G232GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U447 ( .A(n383), .B(KEYINPUT11), .Z(n387) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U450 ( .A(KEYINPUT78), .B(KEYINPUT68), .Z(n389) );
  XNOR2_X1 U451 ( .A(KEYINPUT65), .B(KEYINPUT9), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U453 ( .A(n391), .B(n390), .Z(n394) );
  XOR2_X1 U454 ( .A(G36GAT), .B(G190GAT), .Z(n417) );
  XNOR2_X1 U455 ( .A(n417), .B(n392), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n557) );
  INV_X1 U458 ( .A(n557), .ZN(n397) );
  OR2_X1 U459 ( .A1(n566), .A2(n397), .ZN(n398) );
  NOR2_X1 U460 ( .A1(n399), .A2(n398), .ZN(n401) );
  XNOR2_X1 U461 ( .A(KEYINPUT47), .B(KEYINPUT115), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n407) );
  XNOR2_X1 U463 ( .A(KEYINPUT36), .B(KEYINPUT101), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n402), .B(n557), .ZN(n586) );
  NAND2_X1 U465 ( .A1(n553), .A2(n586), .ZN(n403) );
  XNOR2_X1 U466 ( .A(KEYINPUT45), .B(n403), .ZN(n405) );
  INV_X1 U467 ( .A(n477), .ZN(n579) );
  NAND2_X1 U468 ( .A1(n579), .A2(n574), .ZN(n404) );
  NOR2_X1 U469 ( .A1(n405), .A2(n404), .ZN(n406) );
  NOR2_X1 U470 ( .A1(n407), .A2(n406), .ZN(n409) );
  XOR2_X1 U471 ( .A(KEYINPUT93), .B(n410), .Z(n411) );
  XOR2_X1 U472 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n413) );
  XNOR2_X1 U473 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U475 ( .A(G169GAT), .B(n414), .Z(n441) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n423) );
  XOR2_X1 U477 ( .A(n419), .B(n418), .Z(n421) );
  AND2_X1 U478 ( .A1(G226GAT), .A2(G233GAT), .ZN(n420) );
  NOR2_X1 U479 ( .A1(n544), .A2(n449), .ZN(n424) );
  XNOR2_X1 U480 ( .A(KEYINPUT54), .B(n424), .ZN(n569) );
  NAND2_X1 U481 ( .A1(n425), .A2(n569), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n426), .B(KEYINPUT55), .ZN(n444) );
  XOR2_X1 U483 ( .A(KEYINPUT66), .B(G99GAT), .Z(n428) );
  XNOR2_X1 U484 ( .A(G113GAT), .B(G190GAT), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U486 ( .A(n429), .B(G176GAT), .Z(n432) );
  XNOR2_X1 U487 ( .A(G43GAT), .B(n430), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n437) );
  XOR2_X1 U489 ( .A(G183GAT), .B(n433), .Z(n435) );
  NAND2_X1 U490 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U492 ( .A(n437), .B(n436), .Z(n443) );
  XOR2_X1 U493 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n439) );
  XNOR2_X1 U494 ( .A(KEYINPUT86), .B(G71GAT), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n531) );
  NAND2_X1 U498 ( .A1(n444), .A2(n531), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n445), .B(KEYINPUT122), .ZN(n565) );
  NOR2_X1 U500 ( .A1(n565), .A2(n557), .ZN(n448) );
  INV_X1 U501 ( .A(G190GAT), .ZN(n446) );
  INV_X1 U502 ( .A(G106GAT), .ZN(n476) );
  XOR2_X1 U503 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n474) );
  INV_X1 U504 ( .A(KEYINPUT109), .ZN(n471) );
  XNOR2_X1 U505 ( .A(KEYINPUT37), .B(KEYINPUT103), .ZN(n468) );
  INV_X1 U506 ( .A(KEYINPUT94), .ZN(n451) );
  INV_X1 U507 ( .A(n449), .ZN(n524) );
  XNOR2_X1 U508 ( .A(KEYINPUT27), .B(n524), .ZN(n458) );
  NAND2_X1 U509 ( .A1(n458), .A2(n521), .ZN(n450) );
  XNOR2_X1 U510 ( .A(KEYINPUT28), .B(n456), .ZN(n472) );
  NAND2_X1 U511 ( .A1(n543), .A2(n472), .ZN(n529) );
  XOR2_X1 U512 ( .A(KEYINPUT95), .B(n529), .Z(n452) );
  NOR2_X1 U513 ( .A1(n531), .A2(n452), .ZN(n464) );
  NAND2_X1 U514 ( .A1(n531), .A2(n524), .ZN(n453) );
  XNOR2_X1 U515 ( .A(KEYINPUT96), .B(n453), .ZN(n454) );
  NAND2_X1 U516 ( .A1(n454), .A2(n456), .ZN(n455) );
  XNOR2_X1 U517 ( .A(n455), .B(KEYINPUT25), .ZN(n460) );
  NOR2_X1 U518 ( .A1(n531), .A2(n456), .ZN(n457) );
  XNOR2_X1 U519 ( .A(KEYINPUT26), .B(n457), .ZN(n572) );
  AND2_X1 U520 ( .A1(n458), .A2(n572), .ZN(n459) );
  NOR2_X1 U521 ( .A1(n460), .A2(n459), .ZN(n461) );
  NOR2_X1 U522 ( .A1(n521), .A2(n461), .ZN(n462) );
  XOR2_X1 U523 ( .A(KEYINPUT97), .B(n462), .Z(n463) );
  NOR2_X1 U524 ( .A1(n464), .A2(n463), .ZN(n481) );
  XNOR2_X1 U525 ( .A(n465), .B(KEYINPUT102), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n466), .A2(n586), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n574), .A2(n469), .ZN(n509) );
  NOR2_X1 U528 ( .A1(n491), .A2(n509), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n471), .B(n470), .ZN(n526) );
  INV_X1 U530 ( .A(n472), .ZN(n516) );
  NAND2_X1 U531 ( .A1(n526), .A2(n516), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(G1339GAT) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n484) );
  NOR2_X1 U535 ( .A1(n574), .A2(n477), .ZN(n478) );
  XOR2_X1 U536 ( .A(KEYINPUT76), .B(n478), .Z(n492) );
  NAND2_X1 U537 ( .A1(n553), .A2(n557), .ZN(n479) );
  XNOR2_X1 U538 ( .A(KEYINPUT16), .B(n479), .ZN(n480) );
  NOR2_X1 U539 ( .A1(n481), .A2(n480), .ZN(n482) );
  XOR2_X1 U540 ( .A(KEYINPUT98), .B(n482), .Z(n510) );
  NOR2_X1 U541 ( .A1(n492), .A2(n510), .ZN(n489) );
  NAND2_X1 U542 ( .A1(n521), .A2(n489), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U544 ( .A1(n489), .A2(n524), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n485), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n487) );
  NAND2_X1 U547 ( .A1(n489), .A2(n531), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U549 ( .A(G15GAT), .B(n488), .Z(G1326GAT) );
  NAND2_X1 U550 ( .A1(n516), .A2(n489), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U552 ( .A1(n492), .A2(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(KEYINPUT38), .B(KEYINPUT104), .ZN(n494) );
  NAND2_X1 U554 ( .A1(n493), .A2(n494), .ZN(n498) );
  INV_X1 U555 ( .A(n493), .ZN(n496) );
  INV_X1 U556 ( .A(n494), .ZN(n495) );
  NAND2_X1 U557 ( .A1(n496), .A2(n495), .ZN(n497) );
  NAND2_X1 U558 ( .A1(n498), .A2(n497), .ZN(n506) );
  NAND2_X1 U559 ( .A1(n521), .A2(n506), .ZN(n500) );
  XOR2_X1 U560 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(n501), .ZN(G1328GAT) );
  NAND2_X1 U563 ( .A1(n524), .A2(n506), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(n502), .ZN(G1329GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n504) );
  NAND2_X1 U566 ( .A1(n506), .A2(n531), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n505), .ZN(G1330GAT) );
  NAND2_X1 U569 ( .A1(n516), .A2(n506), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n507), .B(KEYINPUT106), .ZN(n508) );
  XNOR2_X1 U571 ( .A(G50GAT), .B(n508), .ZN(G1331GAT) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n512) );
  NOR2_X1 U573 ( .A1(n510), .A2(n509), .ZN(n517) );
  NAND2_X1 U574 ( .A1(n521), .A2(n517), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(G1332GAT) );
  XOR2_X1 U576 ( .A(G64GAT), .B(KEYINPUT107), .Z(n514) );
  NAND2_X1 U577 ( .A1(n517), .A2(n524), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(G1333GAT) );
  NAND2_X1 U579 ( .A1(n517), .A2(n531), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n526), .A2(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n522), .B(KEYINPUT110), .ZN(n523) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n526), .A2(n524), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT111), .Z(n528) );
  NAND2_X1 U591 ( .A1(n526), .A2(n531), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1338GAT) );
  NOR2_X1 U593 ( .A1(n544), .A2(n529), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n539) );
  NOR2_X1 U595 ( .A1(n574), .A2(n539), .ZN(n532) );
  XOR2_X1 U596 ( .A(G113GAT), .B(n532), .Z(G1340GAT) );
  NOR2_X1 U597 ( .A1(n533), .A2(n539), .ZN(n535) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  INV_X1 U600 ( .A(n539), .ZN(n536) );
  NAND2_X1 U601 ( .A1(n536), .A2(n566), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U604 ( .A1(n557), .A2(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U608 ( .A1(n543), .A2(n572), .ZN(n545) );
  NOR2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n546), .B(KEYINPUT117), .ZN(n556) );
  NOR2_X1 U611 ( .A1(n574), .A2(n556), .ZN(n547) );
  XOR2_X1 U612 ( .A(G141GAT), .B(n547), .Z(G1344GAT) );
  NOR2_X1 U613 ( .A1(n533), .A2(n556), .ZN(n552) );
  XOR2_X1 U614 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n549) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(KEYINPUT53), .B(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  INV_X1 U619 ( .A(n553), .ZN(n583) );
  NOR2_X1 U620 ( .A1(n583), .A2(n556), .ZN(n554) );
  XOR2_X1 U621 ( .A(KEYINPUT120), .B(n554), .Z(n555) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n574), .A2(n565), .ZN(n560) );
  XOR2_X1 U627 ( .A(G169GAT), .B(n560), .Z(G1348GAT) );
  NOR2_X1 U628 ( .A1(n565), .A2(n533), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n562) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n561) );
  XNOR2_X1 U631 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  INV_X1 U633 ( .A(n565), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  AND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT124), .ZN(n585) );
  NOR2_X1 U639 ( .A1(n585), .A2(n574), .ZN(n578) );
  XOR2_X1 U640 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XNOR2_X1 U644 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n581) );
  NOR2_X1 U645 ( .A1(n579), .A2(n585), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n585), .A2(n583), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n589) );
  INV_X1 U651 ( .A(n585), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

