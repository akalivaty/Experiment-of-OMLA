//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n438, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1261, new_n1262,
    new_n1263;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G96), .ZN(new_n438));
  INV_X1    g013(.A(new_n438), .ZN(G221));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G132), .A4(new_n438), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT66), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n461), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n470), .B(G125), .C1(new_n462), .C2(new_n463), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n469), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n467), .B1(new_n475), .B2(G2105), .ZN(G160));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n461), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  OAI221_X1 g061(.A(new_n478), .B1(new_n483), .B2(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  AND2_X1   g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n462), .B2(new_n463), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n462), .B2(new_n463), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n497), .B(new_n500), .C1(new_n463), .C2(new_n462), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n495), .B1(new_n499), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G62), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(KEYINPUT70), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n508), .A2(new_n511), .A3(G62), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n503), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n513), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(G89), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT72), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n514), .A2(new_n527), .A3(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n529), .A2(G51), .B1(new_n508), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n525), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n533), .A2(new_n503), .B1(new_n534), .B2(new_n515), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(G52), .B2(new_n529), .ZN(G171));
  NAND2_X1  g111(.A1(new_n529), .A2(G43), .ZN(new_n537));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(new_n507), .ZN(new_n539));
  NOR2_X1   g114(.A1(KEYINPUT5), .A2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n508), .A2(new_n514), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n543), .A2(G651), .B1(new_n544), .B2(G81), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  AOI22_X1  g126(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n503), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(G65), .B1(new_n539), .B2(new_n540), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT74), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n554), .A2(new_n558), .B1(G91), .B2(new_n544), .ZN(new_n559));
  AND2_X1   g134(.A1(KEYINPUT6), .A2(G651), .ZN(new_n560));
  NOR2_X1   g135(.A1(KEYINPUT6), .A2(G651), .ZN(new_n561));
  OAI211_X1 g136(.A(G53), .B(G543), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n514), .A2(KEYINPUT73), .A3(G53), .A4(G543), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n562), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n559), .A2(new_n570), .ZN(G299));
  NOR2_X1   g146(.A1(G171), .A2(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n529), .A2(G52), .ZN(new_n573));
  NAND2_X1  g148(.A1(G77), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G64), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n541), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(new_n544), .B2(G90), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n572), .A2(new_n580), .ZN(G301));
  NAND2_X1  g156(.A1(new_n525), .A2(new_n531), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  OR2_X1    g158(.A1(new_n508), .A2(G74), .ZN(new_n584));
  INV_X1    g159(.A(new_n517), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n584), .A2(G651), .B1(new_n585), .B2(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n544), .A2(G87), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G288));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n506), .B2(new_n507), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n590), .B2(new_n591), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(G48), .A2(new_n585), .B1(new_n544), .B2(G86), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G305));
  XNOR2_X1  g173(.A(KEYINPUT77), .B(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n529), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G60), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n541), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(new_n544), .B2(G85), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(new_n529), .A2(G54), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n544), .A2(G92), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n607), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n515), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(new_n503), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n606), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  MUX2_X1   g190(.A(new_n615), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g191(.A(new_n615), .B(G301), .S(G868), .Z(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G299), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G168), .B2(new_n618), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(G168), .B2(new_n618), .ZN(G280));
  AND3_X1   g196(.A1(new_n606), .A2(new_n612), .A3(new_n614), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n537), .A2(new_n545), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n618), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n615), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n479), .A2(new_n465), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT13), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n635));
  INV_X1    g210(.A(G135), .ZN(new_n636));
  INV_X1    g211(.A(G123), .ZN(new_n637));
  OAI221_X1 g212(.A(new_n635), .B1(new_n483), .B2(new_n636), .C1(new_n637), .C2(new_n486), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n639), .A3(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(KEYINPUT15), .B(G2435), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT79), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n643), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(new_n656), .A3(G14), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT80), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  NOR3_X1   g238(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT81), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n660), .B(KEYINPUT82), .Z(new_n668));
  AOI21_X1  g243(.A(new_n661), .B1(new_n668), .B2(new_n663), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n663), .B(KEYINPUT17), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n669), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n668), .A2(new_n661), .A3(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n667), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n682), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n683), .A2(KEYINPUT20), .A3(new_n682), .ZN(new_n688));
  OAI221_X1 g263(.A(new_n684), .B1(new_n682), .B2(new_n680), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT84), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n693), .ZN(new_n696));
  AND3_X1   g271(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n695), .B1(new_n694), .B2(new_n696), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(G229));
  XNOR2_X1  g274(.A(KEYINPUT31), .B(G11), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G28), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(KEYINPUT93), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(G28), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n703), .B2(KEYINPUT93), .ZN(new_n706));
  OAI221_X1 g281(.A(new_n700), .B1(new_n704), .B2(new_n706), .C1(new_n638), .C2(new_n701), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NOR2_X1   g283(.A1(G286), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(KEYINPUT92), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G16), .B2(G21), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n710), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n707), .B1(new_n713), .B2(G1966), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n708), .A2(G5), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G171), .B2(new_n708), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT94), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G1961), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n714), .B(new_n718), .C1(G1966), .C2(new_n713), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT95), .Z(new_n720));
  INV_X1    g295(.A(G19), .ZN(new_n721));
  OR3_X1    g296(.A1(new_n721), .A2(KEYINPUT87), .A3(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(KEYINPUT87), .B1(new_n721), .B2(G16), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n722), .B(new_n723), .C1(new_n546), .C2(new_n708), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G1341), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n622), .A2(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G4), .B2(G16), .ZN(new_n727));
  INV_X1    g302(.A(G1348), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n701), .A2(G27), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G164), .B2(new_n701), .ZN(new_n731));
  INV_X1    g306(.A(G2078), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n725), .B(new_n729), .C1(KEYINPUT96), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n701), .A2(G35), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G162), .B2(new_n701), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT29), .B(G2090), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n727), .A2(new_n728), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n733), .A2(KEYINPUT96), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n734), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT26), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n465), .A2(G105), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n486), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G129), .ZN(new_n749));
  INV_X1    g324(.A(new_n483), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G141), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n749), .A2(G29), .A3(new_n751), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(KEYINPUT90), .C1(G29), .C2(G32), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT90), .B2(new_n752), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT27), .B(G1996), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT91), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n754), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n701), .A2(G33), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT25), .Z(new_n760));
  AOI22_X1  g335(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  INV_X1    g336(.A(G139), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n760), .B1(new_n461), .B2(new_n761), .C1(new_n483), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT88), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n758), .B1(new_n764), .B2(new_n701), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2072), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n708), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G1956), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n717), .A2(G1961), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n701), .A2(G26), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT28), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n750), .A2(G140), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n748), .A2(G128), .ZN(new_n777));
  OR2_X1    g352(.A1(G104), .A2(G2105), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n778), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n775), .B1(new_n780), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G34), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(G29), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G160), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2084), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n773), .A2(new_n783), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n742), .A2(new_n757), .A3(new_n772), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n720), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n708), .A2(G22), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G166), .B2(new_n708), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1971), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT85), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n708), .A2(G23), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n585), .A2(G49), .ZN(new_n798));
  OAI21_X1  g373(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n798), .A2(new_n587), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n797), .B1(new_n800), .B2(new_n708), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT33), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1976), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n794), .A2(new_n795), .ZN(new_n804));
  NOR2_X1   g379(.A1(G6), .A2(G16), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n596), .A2(new_n597), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(G16), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT32), .B(G1981), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n796), .A2(new_n803), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n750), .A2(G131), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n748), .A2(G119), .ZN(new_n814));
  OR2_X1    g389(.A1(G95), .A2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G29), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G25), .B2(G29), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  AND2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  MUX2_X1   g398(.A(G24), .B(G290), .S(G16), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1986), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(KEYINPUT86), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n811), .A2(new_n812), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n811), .A2(new_n812), .A3(new_n826), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT86), .B(KEYINPUT36), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n791), .A2(new_n829), .A3(new_n832), .ZN(G150));
  INV_X1    g408(.A(G150), .ZN(G311));
  NAND2_X1  g409(.A1(new_n529), .A2(G55), .ZN(new_n835));
  NAND2_X1  g410(.A1(G80), .A2(G543), .ZN(new_n836));
  INV_X1    g411(.A(G67), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n541), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n838), .A2(G651), .B1(new_n544), .B2(G93), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n835), .A2(KEYINPUT97), .A3(new_n839), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT99), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n625), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n840), .A2(new_n625), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n615), .A2(new_n623), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT98), .ZN(new_n856));
  INV_X1    g431(.A(G860), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n854), .B2(KEYINPUT39), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n847), .B1(new_n856), .B2(new_n858), .ZN(G145));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n764), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT88), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n763), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n763), .A2(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(KEYINPUT100), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n749), .A2(new_n751), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n479), .A2(new_n493), .B1(new_n869), .B2(new_n491), .ZN(new_n870));
  INV_X1    g445(.A(new_n501), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n500), .B1(new_n479), .B2(new_n497), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n749), .A2(G164), .A3(new_n751), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n780), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n780), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  OAI22_X1  g453(.A1(new_n861), .A2(new_n866), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n865), .A2(KEYINPUT100), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n764), .A2(new_n860), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n880), .A2(new_n881), .A3(new_n882), .A4(new_n876), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n879), .A2(new_n883), .A3(KEYINPUT102), .ZN(new_n887));
  OR2_X1    g462(.A1(G106), .A2(G2105), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n888), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n889));
  INV_X1    g464(.A(G142), .ZN(new_n890));
  INV_X1    g465(.A(G130), .ZN(new_n891));
  OAI221_X1 g466(.A(new_n889), .B1(new_n483), .B2(new_n890), .C1(new_n891), .C2(new_n486), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n631), .ZN(new_n893));
  INV_X1    g468(.A(new_n631), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n750), .A2(G142), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n748), .A2(G130), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .A4(new_n889), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n818), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n818), .B1(new_n893), .B2(new_n897), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n886), .A2(new_n887), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n638), .B(G160), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(G162), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n879), .A2(new_n883), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n893), .A2(new_n897), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n817), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n907), .A2(KEYINPUT101), .A3(new_n898), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT101), .B1(new_n907), .B2(new_n898), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n904), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n884), .A2(new_n910), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n884), .A2(new_n910), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n904), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g494(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n622), .A2(new_n559), .A3(new_n570), .ZN(new_n922));
  NAND2_X1  g497(.A1(G299), .A2(new_n615), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n627), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n848), .A2(new_n928), .A3(new_n850), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n546), .B1(new_n842), .B2(new_n843), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n627), .B1(new_n930), .B2(new_n849), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n922), .A2(new_n923), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT103), .B1(new_n933), .B2(new_n924), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n927), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n513), .B2(new_n519), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n513), .A2(new_n936), .A3(new_n519), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n806), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n939), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(G305), .A3(new_n937), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G290), .A2(G288), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n800), .A2(new_n600), .A3(new_n604), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n944), .B2(new_n945), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n940), .B(new_n942), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n922), .A2(new_n923), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n929), .A2(new_n931), .A3(new_n953), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n935), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n952), .B1(new_n935), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n920), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n935), .A2(new_n954), .ZN(new_n958));
  INV_X1    g533(.A(new_n952), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n935), .A2(new_n952), .A3(new_n954), .ZN(new_n961));
  INV_X1    g536(.A(new_n920), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(G868), .ZN(new_n965));
  INV_X1    g540(.A(new_n844), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(G868), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(G295));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n965), .A2(new_n970), .A3(new_n968), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n618), .B1(new_n957), .B2(new_n963), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT107), .B1(new_n972), .B2(new_n967), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(G331));
  XNOR2_X1  g549(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n927), .A2(new_n934), .ZN(new_n977));
  OAI21_X1  g552(.A(G168), .B1(new_n572), .B2(new_n580), .ZN(new_n978));
  AOI21_X1  g553(.A(G171), .B1(new_n525), .B2(new_n531), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n978), .B(new_n980), .C1(new_n930), .C2(new_n849), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n578), .A2(new_n579), .ZN(new_n982));
  NAND2_X1  g557(.A1(G171), .A2(KEYINPUT75), .ZN(new_n983));
  AOI21_X1  g558(.A(G286), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n848), .B(new_n850), .C1(new_n984), .C2(new_n979), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n977), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n985), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n933), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n952), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n917), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n953), .B1(new_n981), .B2(new_n985), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n977), .B2(new_n986), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n948), .A2(new_n951), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n948), .B2(new_n951), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n976), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n925), .A2(new_n926), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(new_n985), .A3(new_n981), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n989), .B2(KEYINPUT110), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n992), .A2(new_n1003), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n1002), .A2(new_n1004), .B1(new_n996), .B2(new_n995), .ZN(new_n1005));
  AOI21_X1  g580(.A(G37), .B1(new_n993), .B2(new_n952), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n975), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n999), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1003), .A2(new_n992), .B1(new_n986), .B2(new_n1000), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1004), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n997), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT43), .B1(new_n1012), .B2(new_n991), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1006), .B(new_n975), .C1(new_n993), .C2(new_n997), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1009), .A2(new_n1015), .ZN(G397));
  XOR2_X1   g591(.A(KEYINPUT111), .B(G1384), .Z(new_n1017));
  NAND2_X1  g592(.A1(new_n873), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n474), .A2(new_n471), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n470), .B1(new_n479), .B2(G125), .ZN(new_n1023));
  OAI21_X1  g598(.A(G2105), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n467), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(G40), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1021), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1996), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n867), .B(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n780), .A2(G2067), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n780), .A2(G2067), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n817), .B(new_n821), .Z(new_n1033));
  OR2_X1    g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G290), .B(G1986), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1027), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT122), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(G1384), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n873), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(new_n873), .B2(new_n1039), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G40), .ZN(new_n1044));
  AOI211_X1 g619(.A(new_n1044), .B(new_n467), .C1(new_n475), .C2(G2105), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1956), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n873), .A2(new_n1039), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1020), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n873), .A2(KEYINPUT45), .A3(new_n1017), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT56), .B(G2072), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1048), .A2(new_n1045), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n544), .A2(G91), .ZN(new_n1054));
  OAI21_X1  g629(.A(G651), .B1(new_n557), .B2(KEYINPUT74), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n552), .A2(new_n553), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1053), .B(KEYINPUT57), .C1(new_n1057), .C2(new_n569), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1053), .A2(KEYINPUT57), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1053), .A2(KEYINPUT57), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n559), .A2(new_n570), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1046), .A2(new_n1052), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1047), .A2(KEYINPUT50), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(new_n1045), .A3(new_n1040), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n770), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1066), .A2(new_n1051), .B1(new_n1061), .B2(new_n1058), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1037), .B(KEYINPUT61), .C1(new_n1063), .C2(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1069), .A2(new_n1037), .A3(new_n1066), .A4(new_n1051), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT61), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1062), .B1(new_n1046), .B2(new_n1052), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1070), .B(new_n1071), .C1(new_n1072), .C2(KEYINPUT122), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT120), .B1(new_n1026), .B2(new_n1047), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G164), .A2(G1384), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1076), .A2(new_n1077), .A3(G40), .A4(G160), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1079), .A2(new_n782), .B1(new_n728), .B2(new_n1065), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n622), .B1(new_n1080), .B2(KEYINPUT60), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n782), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1065), .A2(new_n728), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(KEYINPUT60), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(KEYINPUT123), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(new_n1080), .B2(KEYINPUT60), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1081), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT60), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n615), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1084), .A2(KEYINPUT123), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1080), .A2(new_n1086), .A3(KEYINPUT60), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT58), .B(G1341), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1048), .A2(new_n1045), .A3(new_n1049), .ZN(new_n1096));
  OAI22_X1  g671(.A1(new_n1079), .A2(new_n1095), .B1(G1996), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n546), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT59), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1100), .A3(new_n546), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1074), .A2(new_n1088), .A3(new_n1094), .A4(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1072), .B1(new_n1080), .B2(new_n615), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1069), .A2(new_n1066), .A3(new_n1051), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n615), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1104), .B(new_n1106), .C1(new_n1108), .C2(new_n1067), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1103), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n1113));
  INV_X1    g688(.A(G1961), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1065), .A2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(G164), .A2(G1384), .A3(new_n1019), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT45), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n873), .B2(new_n1039), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n732), .B(new_n1045), .C1(new_n1116), .C2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT53), .B1(new_n1119), .B2(KEYINPUT125), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n873), .A2(new_n1039), .A3(new_n1020), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT45), .B1(G164), .B2(G1384), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1026), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1121), .B1(new_n1124), .B2(new_n732), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1115), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(new_n1115), .C1(new_n1120), .C2(new_n1125), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1096), .B2(G2078), .ZN(new_n1132));
  AOI21_X1  g707(.A(G301), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1132), .A2(G301), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1131), .A2(G2078), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1021), .A2(new_n1045), .A3(new_n1049), .A4(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1115), .A2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1113), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(G1971), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1096), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(G2090), .B2(new_n1065), .ZN(new_n1142));
  NAND3_X1  g717(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT55), .ZN(new_n1144));
  INV_X1    g719(.A(G8), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(G166), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1142), .A2(G8), .A3(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT113), .B(G8), .Z(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1147), .B1(new_n1142), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1150), .B1(new_n1026), .B2(new_n1047), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT114), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT114), .B(new_n1150), .C1(new_n1026), .C2(new_n1047), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n586), .A2(G1976), .A3(new_n587), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT115), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT116), .ZN(new_n1160));
  AOI21_X1  g735(.A(G1976), .B1(new_n586), .B2(new_n587), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n1161), .B2(KEYINPUT52), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT52), .ZN(new_n1163));
  OAI211_X1 g738(.A(KEYINPUT116), .B(new_n1163), .C1(new_n800), .C2(G1976), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1157), .A2(KEYINPUT117), .A3(new_n1159), .A4(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1157), .A2(new_n1159), .A3(new_n1165), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT117), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(G305), .A2(G1981), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(G305), .A2(G1981), .ZN(new_n1172));
  OAI21_X1  g747(.A(KEYINPUT49), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1172), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT49), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1174), .A2(new_n1175), .A3(new_n1170), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1157), .A2(new_n1177), .B1(new_n1178), .B2(KEYINPUT52), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1152), .A2(new_n1166), .A3(new_n1169), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(G2084), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1064), .A2(new_n1045), .A3(new_n1181), .A4(new_n1040), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(new_n1124), .B2(G1966), .ZN(new_n1183));
  NAND2_X1  g758(.A1(G286), .A2(new_n1150), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT51), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1183), .A2(new_n1150), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT124), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1183), .A2(KEYINPUT124), .A3(new_n1150), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1183), .A2(G8), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1188), .B1(new_n1195), .B2(new_n1184), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1187), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1180), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1129), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1119), .A2(KEYINPUT125), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1123), .A2(new_n1122), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1202), .A2(new_n1121), .A3(new_n732), .A4(new_n1045), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1201), .A2(KEYINPUT53), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1128), .B1(new_n1204), .B2(new_n1115), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1134), .B1(new_n1200), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1130), .A2(KEYINPUT127), .A3(new_n1134), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1137), .A2(new_n1132), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1113), .B1(new_n1210), .B2(G171), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  AND4_X1   g787(.A1(new_n1112), .A2(new_n1139), .A3(new_n1199), .A4(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1196), .B1(new_n1193), .B2(new_n1192), .ZN(new_n1214));
  OAI21_X1  g789(.A(KEYINPUT62), .B1(new_n1214), .B2(new_n1187), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1193), .ZN(new_n1217));
  AOI21_X1  g792(.A(KEYINPUT124), .B1(new_n1183), .B2(new_n1150), .ZN(new_n1218));
  NOR3_X1   g793(.A1(new_n1217), .A2(new_n1218), .A3(new_n1189), .ZN(new_n1219));
  OAI211_X1 g794(.A(new_n1216), .B(new_n1186), .C1(new_n1219), .C2(new_n1196), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1177), .A2(new_n1157), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1178), .A2(KEYINPUT52), .ZN(new_n1222));
  NAND4_X1  g797(.A1(new_n1169), .A2(new_n1221), .A3(new_n1222), .A4(new_n1166), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1142), .A2(G8), .A3(new_n1147), .ZN(new_n1224));
  OR2_X1    g799(.A1(new_n1065), .A2(G2090), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1149), .B1(new_n1225), .B2(new_n1141), .ZN(new_n1226));
  OAI21_X1  g801(.A(new_n1224), .B1(new_n1226), .B2(new_n1147), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1223), .A2(new_n1227), .ZN(new_n1228));
  NAND4_X1  g803(.A1(new_n1215), .A2(new_n1220), .A3(new_n1228), .A4(new_n1133), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n1183), .A2(G168), .A3(new_n1150), .ZN(new_n1230));
  NOR3_X1   g805(.A1(new_n1223), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g806(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1147), .B1(new_n1142), .B2(G8), .ZN(new_n1233));
  NOR2_X1   g808(.A1(new_n1233), .A2(new_n1230), .ZN(new_n1234));
  NAND3_X1  g809(.A1(new_n1234), .A2(KEYINPUT63), .A3(new_n1224), .ZN(new_n1235));
  OAI22_X1  g810(.A1(new_n1231), .A2(new_n1232), .B1(new_n1223), .B2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g811(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1237));
  INV_X1    g812(.A(new_n1221), .ZN(new_n1238));
  OR2_X1    g813(.A1(G288), .A2(G1976), .ZN(new_n1239));
  OAI21_X1  g814(.A(new_n1174), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g815(.A(new_n1237), .B1(new_n1157), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g816(.A1(new_n1229), .A2(new_n1236), .A3(new_n1241), .ZN(new_n1242));
  OAI21_X1  g817(.A(new_n1036), .B1(new_n1213), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1034), .A2(new_n1027), .ZN(new_n1244));
  NOR2_X1   g819(.A1(G290), .A2(G1986), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1027), .A2(new_n1245), .ZN(new_n1246));
  XNOR2_X1  g821(.A(new_n1246), .B(KEYINPUT48), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n818), .A2(new_n821), .ZN(new_n1248));
  OAI21_X1  g823(.A(new_n1031), .B1(new_n1032), .B2(new_n1248), .ZN(new_n1249));
  AOI22_X1  g824(.A1(new_n1244), .A2(new_n1247), .B1(new_n1027), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1031), .A2(new_n1030), .ZN(new_n1251));
  OAI21_X1  g826(.A(new_n1027), .B1(new_n1251), .B2(new_n867), .ZN(new_n1252));
  NOR3_X1   g827(.A1(new_n1021), .A2(G1996), .A3(new_n1026), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1253), .A2(KEYINPUT46), .ZN(new_n1254));
  OR2_X1    g829(.A1(new_n1253), .A2(KEYINPUT46), .ZN(new_n1255));
  NAND3_X1  g830(.A1(new_n1252), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  XNOR2_X1  g831(.A(new_n1256), .B(KEYINPUT47), .ZN(new_n1257));
  AND2_X1   g832(.A1(new_n1250), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g833(.A1(new_n1243), .A2(new_n1258), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g834(.A1(new_n999), .A2(new_n1007), .ZN(new_n1261));
  NAND3_X1  g835(.A1(new_n675), .A2(G319), .A3(new_n657), .ZN(new_n1262));
  NOR3_X1   g836(.A1(new_n1262), .A2(new_n697), .A3(new_n698), .ZN(new_n1263));
  NAND3_X1  g837(.A1(new_n1261), .A2(new_n918), .A3(new_n1263), .ZN(G225));
  INV_X1    g838(.A(G225), .ZN(G308));
endmodule


