

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  NOR2_X1 U323 ( .A1(n513), .A2(n415), .ZN(n568) );
  XNOR2_X1 U324 ( .A(KEYINPUT109), .B(KEYINPUT46), .ZN(n367) );
  XNOR2_X1 U325 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U326 ( .A(n408), .B(n363), .ZN(n364) );
  XNOR2_X1 U327 ( .A(n365), .B(n364), .ZN(n393) );
  XNOR2_X1 U328 ( .A(n435), .B(KEYINPUT55), .ZN(n452) );
  INV_X1 U329 ( .A(G183GAT), .ZN(n456) );
  XNOR2_X1 U330 ( .A(n451), .B(n450), .ZN(n527) );
  XNOR2_X1 U331 ( .A(n456), .B(KEYINPUT118), .ZN(n457) );
  XNOR2_X1 U332 ( .A(n458), .B(n457), .ZN(G1350GAT) );
  XOR2_X1 U333 ( .A(G113GAT), .B(G36GAT), .Z(n292) );
  XOR2_X1 U334 ( .A(G169GAT), .B(G8GAT), .Z(n401) );
  XOR2_X1 U335 ( .A(G15GAT), .B(G22GAT), .Z(n343) );
  XNOR2_X1 U336 ( .A(n401), .B(n343), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U338 ( .A(n293), .B(G50GAT), .Z(n299) );
  XNOR2_X1 U339 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n294), .B(KEYINPUT7), .ZN(n382) );
  XOR2_X1 U341 ( .A(n382), .B(KEYINPUT67), .Z(n296) );
  NAND2_X1 U342 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n297), .B(G29GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n307) );
  XOR2_X1 U346 ( .A(KEYINPUT64), .B(G1GAT), .Z(n301) );
  XNOR2_X1 U347 ( .A(G141GAT), .B(G197GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U349 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n303) );
  XNOR2_X1 U350 ( .A(KEYINPUT30), .B(KEYINPUT65), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U352 ( .A(n305), .B(n304), .Z(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n528) );
  XOR2_X1 U354 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n309) );
  XNOR2_X1 U355 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n326) );
  XOR2_X1 U357 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n311) );
  XNOR2_X1 U358 ( .A(KEYINPUT6), .B(KEYINPUT94), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U360 ( .A(n312), .B(G85GAT), .Z(n314) );
  XOR2_X1 U361 ( .A(G1GAT), .B(G127GAT), .Z(n342) );
  XNOR2_X1 U362 ( .A(G162GAT), .B(n342), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n319) );
  XNOR2_X1 U364 ( .A(G120GAT), .B(G148GAT), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n315), .B(G57GAT), .ZN(n349) );
  XOR2_X1 U366 ( .A(G29GAT), .B(G134GAT), .Z(n377) );
  XOR2_X1 U367 ( .A(n349), .B(n377), .Z(n317) );
  NAND2_X1 U368 ( .A1(G225GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U370 ( .A(n319), .B(n318), .Z(n324) );
  XNOR2_X1 U371 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n320), .B(KEYINPUT84), .ZN(n436) );
  XOR2_X1 U373 ( .A(G155GAT), .B(KEYINPUT2), .Z(n322) );
  XNOR2_X1 U374 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n422) );
  XNOR2_X1 U376 ( .A(n436), .B(n422), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U378 ( .A(n326), .B(n325), .Z(n468) );
  XNOR2_X1 U379 ( .A(KEYINPUT95), .B(n468), .ZN(n513) );
  INV_X1 U380 ( .A(KEYINPUT54), .ZN(n414) );
  XOR2_X1 U381 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n328) );
  XNOR2_X1 U382 ( .A(KEYINPUT12), .B(KEYINPUT79), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n347) );
  XOR2_X1 U384 ( .A(G78GAT), .B(G211GAT), .Z(n330) );
  XNOR2_X1 U385 ( .A(G183GAT), .B(G155GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U387 ( .A(KEYINPUT14), .B(KEYINPUT78), .Z(n332) );
  XNOR2_X1 U388 ( .A(G8GAT), .B(G64GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U390 ( .A(n334), .B(n333), .Z(n339) );
  XOR2_X1 U391 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n336) );
  NAND2_X1 U392 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U394 ( .A(G57GAT), .B(n337), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n341) );
  XNOR2_X1 U396 ( .A(G71GAT), .B(KEYINPUT68), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n340), .B(KEYINPUT13), .ZN(n348) );
  XOR2_X1 U398 ( .A(n341), .B(n348), .Z(n345) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n533) );
  INV_X1 U402 ( .A(n533), .ZN(n578) );
  INV_X1 U403 ( .A(KEYINPUT41), .ZN(n366) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n355) );
  XOR2_X1 U405 ( .A(KEYINPUT70), .B(KEYINPUT31), .Z(n351) );
  NAND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n353) );
  INV_X1 U408 ( .A(KEYINPUT69), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U411 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n357) );
  XNOR2_X1 U412 ( .A(KEYINPUT73), .B(KEYINPUT71), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U414 ( .A(n359), .B(n358), .Z(n365) );
  XOR2_X1 U415 ( .A(G92GAT), .B(G64GAT), .Z(n361) );
  XNOR2_X1 U416 ( .A(G176GAT), .B(KEYINPUT72), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U418 ( .A(G204GAT), .B(n362), .Z(n408) );
  XOR2_X1 U419 ( .A(G106GAT), .B(G78GAT), .Z(n425) );
  XOR2_X1 U420 ( .A(G99GAT), .B(G85GAT), .Z(n376) );
  XNOR2_X1 U421 ( .A(n425), .B(n376), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n366), .B(n393), .ZN(n501) );
  OR2_X1 U423 ( .A1(n501), .A2(n528), .ZN(n368) );
  NOR2_X1 U424 ( .A1(n578), .A2(n369), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n370), .B(KEYINPUT110), .ZN(n389) );
  XOR2_X1 U426 ( .A(KEYINPUT76), .B(KEYINPUT74), .Z(n372) );
  XNOR2_X1 U427 ( .A(KEYINPUT11), .B(KEYINPUT75), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n388) );
  XOR2_X1 U429 ( .A(KEYINPUT9), .B(G92GAT), .Z(n374) );
  NAND2_X1 U430 ( .A1(G232GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U432 ( .A(G106GAT), .B(n375), .ZN(n386) );
  XOR2_X1 U433 ( .A(KEYINPUT10), .B(n376), .Z(n379) );
  XNOR2_X1 U434 ( .A(G218GAT), .B(n377), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n381) );
  XNOR2_X1 U436 ( .A(G36GAT), .B(G190GAT), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n380), .B(KEYINPUT77), .ZN(n404) );
  XOR2_X1 U438 ( .A(n381), .B(n404), .Z(n384) );
  XOR2_X1 U439 ( .A(G50GAT), .B(G162GAT), .Z(n426) );
  XNOR2_X1 U440 ( .A(n382), .B(n426), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U443 ( .A(n388), .B(n387), .Z(n551) );
  INV_X1 U444 ( .A(n551), .ZN(n561) );
  NAND2_X1 U445 ( .A1(n389), .A2(n561), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n390), .B(KEYINPUT47), .ZN(n397) );
  XOR2_X1 U447 ( .A(KEYINPUT36), .B(n561), .Z(n580) );
  NAND2_X1 U448 ( .A1(n580), .A2(n578), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n391), .B(KEYINPUT111), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n392), .B(KEYINPUT45), .ZN(n394) );
  NAND2_X1 U451 ( .A1(n394), .A2(n393), .ZN(n395) );
  INV_X1 U452 ( .A(n528), .ZN(n570) );
  NOR2_X1 U453 ( .A1(n395), .A2(n570), .ZN(n396) );
  NOR2_X1 U454 ( .A1(n397), .A2(n396), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n398), .B(KEYINPUT48), .ZN(n542) );
  XOR2_X1 U456 ( .A(G211GAT), .B(KEYINPUT21), .Z(n400) );
  XNOR2_X1 U457 ( .A(G197GAT), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n421) );
  XOR2_X1 U459 ( .A(KEYINPUT96), .B(n401), .Z(n403) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U462 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U463 ( .A(G183GAT), .B(KEYINPUT17), .Z(n407) );
  XNOR2_X1 U464 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n407), .B(n406), .ZN(n449) );
  XNOR2_X1 U466 ( .A(n449), .B(n408), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n421), .B(n411), .ZN(n515) );
  INV_X1 U469 ( .A(n515), .ZN(n412) );
  NOR2_X1 U470 ( .A1(n542), .A2(n412), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U472 ( .A(G148GAT), .B(G204GAT), .Z(n417) );
  XNOR2_X1 U473 ( .A(KEYINPUT90), .B(KEYINPUT88), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n434) );
  XOR2_X1 U475 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n419) );
  NAND2_X1 U476 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U478 ( .A(n420), .B(KEYINPUT24), .Z(n424) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U481 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n428) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U484 ( .A(n430), .B(n429), .Z(n432) );
  XNOR2_X1 U485 ( .A(G22GAT), .B(KEYINPUT86), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n471) );
  NAND2_X1 U488 ( .A1(n568), .A2(n471), .ZN(n435) );
  XOR2_X1 U489 ( .A(G134GAT), .B(n436), .Z(n438) );
  NAND2_X1 U490 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U492 ( .A(G127GAT), .B(KEYINPUT20), .Z(n440) );
  XNOR2_X1 U493 ( .A(G176GAT), .B(KEYINPUT85), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U495 ( .A(n442), .B(n441), .Z(n447) );
  XOR2_X1 U496 ( .A(G120GAT), .B(G190GAT), .Z(n444) );
  XNOR2_X1 U497 ( .A(G169GAT), .B(G99GAT), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U501 ( .A(n448), .B(G71GAT), .Z(n451) );
  XNOR2_X1 U502 ( .A(G15GAT), .B(n449), .ZN(n450) );
  NAND2_X1 U503 ( .A1(n452), .A2(n527), .ZN(n560) );
  NOR2_X1 U504 ( .A1(n528), .A2(n560), .ZN(n455) );
  INV_X1 U505 ( .A(G169GAT), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n453), .B(KEYINPUT116), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(G1348GAT) );
  NOR2_X1 U508 ( .A1(n533), .A2(n560), .ZN(n458) );
  NAND2_X1 U509 ( .A1(n570), .A2(n393), .ZN(n491) );
  NAND2_X1 U510 ( .A1(n561), .A2(n578), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n459), .B(KEYINPUT16), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT83), .ZN(n476) );
  NOR2_X1 U513 ( .A1(n527), .A2(n471), .ZN(n462) );
  XNOR2_X1 U514 ( .A(KEYINPUT26), .B(KEYINPUT98), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n462), .B(n461), .ZN(n567) );
  XNOR2_X1 U516 ( .A(n515), .B(KEYINPUT27), .ZN(n470) );
  NAND2_X1 U517 ( .A1(n567), .A2(n470), .ZN(n467) );
  AND2_X1 U518 ( .A1(n515), .A2(n527), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n463), .B(KEYINPUT99), .ZN(n464) );
  NAND2_X1 U520 ( .A1(n464), .A2(n471), .ZN(n465) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n465), .Z(n466) );
  NAND2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n469) );
  NAND2_X1 U523 ( .A1(n469), .A2(n468), .ZN(n475) );
  AND2_X1 U524 ( .A1(n513), .A2(n470), .ZN(n540) );
  XOR2_X1 U525 ( .A(KEYINPUT28), .B(n471), .Z(n519) );
  INV_X1 U526 ( .A(n519), .ZN(n472) );
  NAND2_X1 U527 ( .A1(n540), .A2(n472), .ZN(n525) );
  NOR2_X1 U528 ( .A1(n527), .A2(n525), .ZN(n473) );
  XNOR2_X1 U529 ( .A(KEYINPUT97), .B(n473), .ZN(n474) );
  NAND2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n488) );
  NAND2_X1 U531 ( .A1(n476), .A2(n488), .ZN(n502) );
  NOR2_X1 U532 ( .A1(n491), .A2(n502), .ZN(n484) );
  NAND2_X1 U533 ( .A1(n513), .A2(n484), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n477), .B(KEYINPUT34), .ZN(n478) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n478), .ZN(G1324GAT) );
  NAND2_X1 U536 ( .A1(n515), .A2(n484), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n479), .B(KEYINPUT100), .ZN(n480) );
  XNOR2_X1 U538 ( .A(G8GAT), .B(n480), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n482) );
  NAND2_X1 U540 ( .A1(n484), .A2(n527), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U542 ( .A(G15GAT), .B(n483), .Z(G1326GAT) );
  NAND2_X1 U543 ( .A1(n519), .A2(n484), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n487) );
  XNOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n494) );
  NAND2_X1 U548 ( .A1(n580), .A2(n488), .ZN(n489) );
  NOR2_X1 U549 ( .A1(n578), .A2(n489), .ZN(n490) );
  XNOR2_X1 U550 ( .A(KEYINPUT37), .B(n490), .ZN(n512) );
  NOR2_X1 U551 ( .A1(n512), .A2(n491), .ZN(n492) );
  XNOR2_X1 U552 ( .A(KEYINPUT38), .B(n492), .ZN(n498) );
  NAND2_X1 U553 ( .A1(n498), .A2(n513), .ZN(n493) );
  XOR2_X1 U554 ( .A(n494), .B(n493), .Z(G1328GAT) );
  NAND2_X1 U555 ( .A1(n515), .A2(n498), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(n495), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n498), .A2(n527), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n519), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(KEYINPUT104), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  INV_X1 U564 ( .A(n501), .ZN(n544) );
  NAND2_X1 U565 ( .A1(n544), .A2(n528), .ZN(n511) );
  NOR2_X1 U566 ( .A1(n511), .A2(n502), .ZN(n508) );
  NAND2_X1 U567 ( .A1(n508), .A2(n513), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n515), .A2(n508), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U571 ( .A(G71GAT), .B(KEYINPUT105), .Z(n507) );
  NAND2_X1 U572 ( .A1(n508), .A2(n527), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U575 ( .A1(n508), .A2(n519), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NOR2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n520), .A2(n513), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n515), .A2(n520), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(KEYINPUT106), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n520), .A2(n527), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(KEYINPUT107), .ZN(n524) );
  XOR2_X1 U586 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n522) );
  NAND2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n542), .A2(n525), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n537) );
  NOR2_X1 U592 ( .A1(n528), .A2(n537), .ZN(n529) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n529), .Z(G1340GAT) );
  NOR2_X1 U594 ( .A1(n501), .A2(n537), .ZN(n531) );
  XNOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT112), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(n532), .ZN(G1341GAT) );
  NOR2_X1 U598 ( .A1(n533), .A2(n537), .ZN(n535) );
  XNOR2_X1 U599 ( .A(KEYINPUT113), .B(KEYINPUT50), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  NOR2_X1 U602 ( .A1(n561), .A2(n537), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n567), .A2(n540), .ZN(n541) );
  NOR2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n552), .A2(n570), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n543), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT114), .ZN(n548) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  NAND2_X1 U611 ( .A1(n552), .A2(n544), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  XOR2_X1 U614 ( .A(G155GAT), .B(KEYINPUT115), .Z(n550) );
  NAND2_X1 U615 ( .A1(n552), .A2(n578), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U619 ( .A1(n560), .A2(n501), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT117), .Z(n555) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT119), .B(KEYINPUT58), .Z(n559) );
  XNOR2_X1 U625 ( .A(G190GAT), .B(KEYINPUT120), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n563) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(n563), .B(n562), .Z(G1351GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n565) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT122), .B(n566), .Z(n572) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT121), .B(n569), .Z(n573) );
  INV_X1 U635 ( .A(n573), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n581), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n393), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n575) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n585) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1355GAT) );
endmodule

