//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1262, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT64), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n214), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G20), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n202), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n217), .B1(KEYINPUT1), .B2(new_n224), .C1(new_n227), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  OAI211_X1 g0050(.A(G232), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  OAI211_X1 g0052(.A(G226), .B(new_n252), .C1(new_n249), .C2(new_n250), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G97), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n225), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT13), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n257), .A2(G274), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n257), .A2(G238), .A3(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n259), .A2(new_n260), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT73), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n259), .A2(new_n267), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT13), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n259), .A2(KEYINPUT73), .A3(new_n267), .A4(new_n260), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n270), .A2(new_n272), .A3(G190), .A4(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G13), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n275), .A2(new_n212), .A3(G1), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT74), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT12), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n276), .B(new_n228), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n278), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n228), .A2(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n212), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G77), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n282), .B1(new_n283), .B2(new_n284), .C1(new_n286), .C2(new_n201), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G1), .A2(G13), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(KEYINPUT11), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n211), .B2(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G68), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n281), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT11), .B1(new_n287), .B2(new_n290), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n259), .A2(new_n260), .A3(new_n267), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n260), .B1(new_n259), .B2(new_n267), .ZN(new_n298));
  OAI21_X1  g0098(.A(G200), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n274), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(new_n270), .A3(new_n273), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n272), .A2(new_n268), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT14), .B1(new_n305), .B2(G169), .ZN(new_n306));
  OAI211_X1 g0106(.A(KEYINPUT14), .B(G169), .C1(new_n297), .C2(new_n298), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n304), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n296), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n301), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT68), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n312), .A2(new_n313), .B1(G150), .B2(new_n285), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT8), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G58), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT67), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT8), .B(G58), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT67), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n314), .B1(new_n313), .B2(new_n312), .C1(new_n323), .C2(new_n283), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n290), .ZN(new_n325));
  OAI21_X1  g0125(.A(G50), .B1(new_n212), .B2(G1), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT69), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n276), .A2(new_n290), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n327), .A2(new_n328), .B1(new_n201), .B2(new_n276), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n257), .A2(new_n265), .ZN(new_n331));
  INV_X1    g0131(.A(G226), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n264), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OR2_X1    g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NAND2_X1  g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(G222), .A3(new_n252), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(G223), .A3(G1698), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n338), .C1(new_n284), .C2(new_n336), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n333), .B1(new_n339), .B2(new_n258), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n302), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n330), .B(new_n341), .C1(G169), .C2(new_n340), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT71), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n336), .A2(G238), .A3(G1698), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n249), .A2(new_n250), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G107), .ZN(new_n346));
  OAI211_X1 g0146(.A(G232), .B(new_n252), .C1(new_n249), .C2(new_n250), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n258), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n257), .A2(G244), .A3(new_n265), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n264), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n343), .B1(new_n353), .B2(G179), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n348), .B2(new_n258), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(KEYINPUT71), .A3(new_n302), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n359), .A2(new_n283), .B1(new_n212), .B2(new_n284), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n320), .A2(new_n286), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n290), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n276), .A2(new_n284), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n292), .A2(G77), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n354), .A2(new_n356), .A3(new_n358), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n355), .A2(G190), .ZN(new_n367));
  INV_X1    g0167(.A(new_n365), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT70), .B(G200), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n367), .B(new_n368), .C1(new_n369), .C2(new_n355), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n342), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT9), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n330), .B(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n340), .A2(new_n369), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n374), .A2(KEYINPUT72), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n374), .A2(KEYINPUT72), .B1(G190), .B2(new_n340), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n373), .A2(new_n377), .A3(KEYINPUT10), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT10), .B1(new_n373), .B2(new_n377), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n371), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n229), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G20), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT75), .ZN(new_n386));
  INV_X1    g0186(.A(G159), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n385), .B(new_n386), .C1(new_n387), .C2(new_n286), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n286), .A2(new_n387), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n212), .B1(new_n229), .B2(new_n383), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT75), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n336), .B2(G20), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n345), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n228), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n382), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n336), .A2(new_n393), .A3(G20), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT7), .B1(new_n345), .B2(new_n212), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n400), .A2(KEYINPUT16), .A3(new_n388), .A4(new_n391), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n290), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n275), .A2(G1), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G20), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n323), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n290), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(G1), .B2(new_n212), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n319), .A3(new_n322), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n405), .A2(new_n408), .A3(KEYINPUT76), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT76), .B1(new_n405), .B2(new_n408), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n402), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n332), .A2(G1698), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n413), .B1(G223), .B2(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n257), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n257), .A2(G232), .A3(new_n265), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n264), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  MUX2_X1   g0219(.A(G169), .B(G179), .S(new_n419), .Z(new_n420));
  NAND2_X1  g0220(.A1(new_n412), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n402), .A2(new_n411), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n414), .A2(new_n415), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n258), .ZN(new_n425));
  INV_X1    g0225(.A(new_n418), .ZN(new_n426));
  INV_X1    g0226(.A(G190), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G200), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n416), .B2(new_n418), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(KEYINPUT77), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT77), .B1(new_n428), .B2(new_n430), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n423), .A2(KEYINPUT17), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n428), .A2(new_n430), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT77), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n402), .A2(new_n438), .A3(new_n431), .A4(new_n411), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n412), .A2(new_n420), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n422), .A2(new_n435), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT78), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n444), .A2(KEYINPUT78), .ZN(new_n446));
  AND4_X1   g0246(.A1(new_n311), .A2(new_n381), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(G257), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n449));
  OAI211_X1 g0249(.A(G250), .B(new_n252), .C1(new_n249), .C2(new_n250), .ZN(new_n450));
  INV_X1    g0250(.A(G33), .ZN(new_n451));
  INV_X1    g0251(.A(G294), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n449), .B(new_n450), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n258), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n211), .B(G45), .C1(new_n261), .C2(KEYINPUT5), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G41), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n459), .A2(KEYINPUT79), .A3(new_n211), .A4(G45), .ZN(new_n460));
  INV_X1    g0260(.A(G274), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n225), .B2(new_n256), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n458), .A2(G41), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n457), .A2(new_n460), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n257), .B(G264), .C1(new_n455), .C2(new_n463), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n454), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n357), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(G179), .B2(new_n467), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT24), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT23), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n212), .B2(G107), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G116), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n451), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n212), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n212), .B(G87), .C1(new_n249), .C2(new_n250), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT22), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT22), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n336), .A2(new_n481), .A3(new_n212), .A4(G87), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n478), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n470), .B1(new_n483), .B2(KEYINPUT82), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(KEYINPUT82), .B2(new_n483), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n483), .A2(KEYINPUT82), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n406), .B1(new_n486), .B2(new_n470), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n276), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT25), .B1(new_n276), .B2(new_n206), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n211), .A2(G33), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n406), .A2(new_n404), .A3(new_n491), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n489), .A2(new_n490), .B1(new_n492), .B2(new_n206), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n469), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n493), .B1(new_n485), .B2(new_n487), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT83), .B1(new_n467), .B2(G190), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n467), .A2(new_n429), .ZN(new_n499));
  INV_X1    g0299(.A(new_n466), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n258), .B2(new_n453), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT83), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(new_n427), .A4(new_n465), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n498), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n406), .A2(new_n404), .A3(new_n491), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(KEYINPUT81), .A3(G116), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT81), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n492), .B2(new_n475), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n212), .C1(G33), .C2(new_n205), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n475), .A2(G20), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n290), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT20), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n290), .A4(new_n514), .ZN(new_n518));
  INV_X1    g0318(.A(new_n514), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n517), .A2(new_n518), .B1(new_n403), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G264), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n522));
  OAI211_X1 g0322(.A(G257), .B(new_n252), .C1(new_n249), .C2(new_n250), .ZN(new_n523));
  INV_X1    g0323(.A(G303), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n522), .B(new_n523), .C1(new_n524), .C2(new_n336), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n258), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n257), .B(G270), .C1(new_n455), .C2(new_n463), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n465), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G200), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n521), .B(new_n529), .C1(new_n427), .C2(new_n528), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT21), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(G169), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n531), .B1(new_n521), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n511), .A2(new_n520), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n534), .A2(KEYINPUT21), .A3(G169), .A4(new_n528), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n526), .A2(G179), .A3(new_n465), .A4(new_n527), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n534), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n530), .A2(new_n533), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  AND2_X1   g0339(.A1(KEYINPUT4), .A2(G244), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n252), .B(new_n540), .C1(new_n249), .C2(new_n250), .ZN(new_n541));
  INV_X1    g0341(.A(G244), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n334), .B2(new_n335), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n541), .B(new_n512), .C1(new_n543), .C2(KEYINPUT4), .ZN(new_n544));
  OAI21_X1  g0344(.A(G250), .B1(new_n249), .B2(new_n250), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n252), .B1(new_n545), .B2(KEYINPUT4), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n258), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n257), .B(G257), .C1(new_n455), .C2(new_n463), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n465), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G190), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n552), .A2(new_n205), .A3(G107), .ZN(new_n553));
  XNOR2_X1  g0353(.A(G97), .B(G107), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n555), .A2(new_n212), .B1(new_n284), .B2(new_n286), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n206), .B1(new_n394), .B2(new_n395), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n290), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n404), .A2(G97), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n507), .B2(G97), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n547), .A2(new_n549), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G200), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n551), .A2(new_n558), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n550), .A2(new_n302), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n558), .A2(new_n560), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n357), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n336), .A2(new_n212), .A3(G68), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT19), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n212), .B1(new_n254), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G87), .B2(new_n207), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n283), .B2(new_n205), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n569), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n290), .B1(new_n276), .B2(new_n359), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n507), .A2(G87), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n211), .A2(new_n461), .A3(G45), .ZN(new_n578));
  INV_X1    g0378(.A(G250), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n262), .B2(G1), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n257), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(G244), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n583));
  OAI211_X1 g0383(.A(G238), .B(new_n252), .C1(new_n249), .C2(new_n250), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n583), .B(new_n584), .C1(new_n451), .C2(new_n475), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n582), .B1(new_n585), .B2(new_n258), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G190), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n577), .B(new_n587), .C1(new_n369), .C2(new_n586), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT80), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n492), .B2(new_n359), .ZN(new_n590));
  INV_X1    g0390(.A(new_n359), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n507), .A2(KEYINPUT80), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n575), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n585), .A2(new_n258), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n581), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n357), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n593), .B(new_n596), .C1(G179), .C2(new_n595), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n588), .A2(new_n597), .ZN(new_n598));
  OR3_X1    g0398(.A1(new_n539), .A2(new_n568), .A3(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n448), .A2(new_n506), .A3(new_n599), .ZN(G372));
  INV_X1    g0400(.A(KEYINPUT86), .ZN(new_n601));
  INV_X1    g0401(.A(new_n380), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n378), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n379), .A2(KEYINPUT86), .A3(new_n380), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n412), .A2(new_n442), .A3(new_n420), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n442), .B1(new_n412), .B2(new_n420), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n309), .A2(new_n310), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n301), .B2(new_n366), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n439), .B(KEYINPUT17), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n605), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n614), .A2(new_n342), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT84), .ZN(new_n616));
  INV_X1    g0416(.A(new_n369), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n595), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT84), .B1(new_n586), .B2(new_n369), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n577), .A2(new_n618), .A3(new_n587), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n597), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n622), .A2(new_n505), .A3(new_n567), .A4(new_n563), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n495), .A2(KEYINPUT85), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT85), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n497), .B2(new_n469), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n533), .A2(new_n535), .A3(new_n538), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n623), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n621), .A2(new_n567), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT26), .B1(new_n598), .B2(new_n567), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n597), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n615), .B1(new_n448), .B2(new_n636), .ZN(G369));
  NAND2_X1  g0437(.A1(new_n403), .A2(new_n212), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n497), .A2(new_n644), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n506), .A2(new_n645), .B1(new_n496), .B2(new_n644), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT88), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT88), .ZN(new_n648));
  OAI221_X1 g0448(.A(new_n648), .B1(new_n496), .B2(new_n644), .C1(new_n506), .C2(new_n645), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n628), .A2(new_n644), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n627), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n650), .A2(new_n652), .B1(new_n653), .B2(new_n644), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n534), .A2(new_n643), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT87), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n629), .A2(new_n530), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n629), .B2(new_n656), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G330), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n650), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0463(.A(new_n215), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G1), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n230), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT28), .ZN(new_n670));
  INV_X1    g0470(.A(G330), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT31), .B1(new_n599), .B2(new_n506), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n586), .A2(G179), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n561), .A2(KEYINPUT93), .A3(new_n467), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT93), .B1(new_n561), .B2(new_n467), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n528), .B(new_n673), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT90), .B1(new_n501), .B2(new_n586), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n677), .A2(new_n536), .A3(new_n561), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n501), .A2(new_n586), .A3(KEYINPUT90), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(KEYINPUT30), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT94), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n561), .A2(new_n536), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n501), .A2(new_n586), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT90), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n683), .A2(new_n686), .A3(KEYINPUT91), .A4(new_n679), .ZN(new_n687));
  XOR2_X1   g0487(.A(KEYINPUT92), .B(KEYINPUT30), .Z(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT91), .B1(new_n678), .B2(new_n679), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n682), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n683), .A2(new_n679), .A3(new_n686), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT91), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(KEYINPUT94), .A3(new_n687), .A4(new_n688), .ZN(new_n695));
  AOI211_X1 g0495(.A(KEYINPUT31), .B(new_n681), .C1(new_n691), .C2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n672), .B1(new_n696), .B2(new_n644), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n643), .A2(KEYINPUT31), .ZN(new_n698));
  INV_X1    g0498(.A(new_n681), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n694), .A2(new_n687), .A3(new_n688), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n671), .B1(new_n697), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT96), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n568), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n563), .A2(new_n567), .A3(KEYINPUT96), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n622), .B(new_n505), .C1(new_n628), .C2(new_n495), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n567), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n632), .A3(new_n588), .A4(new_n597), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n712), .B(new_n597), .C1(new_n631), .C2(new_n632), .ZN(new_n713));
  OAI211_X1 g0513(.A(KEYINPUT29), .B(new_n644), .C1(new_n710), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n636), .A2(new_n643), .ZN(new_n715));
  XOR2_X1   g0515(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n704), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n670), .B1(new_n718), .B2(G1), .ZN(G364));
  NOR2_X1   g0519(.A1(new_n275), .A2(G20), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n211), .B1(new_n720), .B2(G45), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n665), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n660), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(G330), .B2(new_n658), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n215), .A2(new_n336), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n209), .A2(new_n726), .B1(G116), .B2(new_n215), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n244), .A2(G45), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n664), .A2(new_n336), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n230), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n730), .B1(new_n262), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n727), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n212), .B1(KEYINPUT97), .B2(new_n357), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n357), .A2(KEYINPUT97), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n289), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT98), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n723), .B1(new_n733), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n212), .A2(G190), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n617), .A2(new_n302), .A3(new_n743), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT102), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(KEYINPUT102), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G107), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n212), .B1(new_n750), .B2(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n205), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n743), .A2(new_n750), .ZN(new_n753));
  XNOR2_X1  g0553(.A(KEYINPUT100), .B(G159), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT101), .B(KEYINPUT32), .Z(new_n756));
  NAND3_X1  g0556(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n427), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n755), .A2(new_n756), .B1(new_n201), .B2(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n752), .B(new_n760), .C1(new_n755), .C2(new_n756), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n302), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n743), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT99), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G77), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n212), .A2(new_n427), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n762), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n757), .A2(G190), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n336), .B1(new_n772), .B2(new_n202), .C1(new_n228), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n771), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n776), .A2(new_n369), .A3(G179), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(G87), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n749), .A2(new_n761), .A3(new_n770), .A4(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G329), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n345), .B1(new_n753), .B2(new_n780), .C1(new_n772), .C2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n769), .B2(G311), .ZN(new_n783));
  INV_X1    g0583(.A(G326), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n759), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g0585(.A1(KEYINPUT33), .A2(G317), .ZN(new_n786));
  NAND2_X1  g0586(.A1(KEYINPUT33), .A2(G317), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n774), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n751), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n785), .B(new_n788), .C1(G294), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n777), .A2(G303), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n783), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n747), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n779), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n742), .B1(new_n795), .B2(new_n736), .ZN(new_n796));
  INV_X1    g0596(.A(new_n739), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n658), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n725), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  NOR2_X1   g0600(.A1(new_n759), .A2(new_n524), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n752), .B(new_n801), .C1(G283), .C2(new_n773), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n748), .A2(G87), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n777), .A2(G107), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n345), .B1(new_n753), .B2(new_n805), .C1(new_n772), .C2(new_n452), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n769), .B2(G116), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n802), .A2(new_n803), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT103), .ZN(new_n809));
  INV_X1    g0609(.A(G150), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n774), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  INV_X1    g0612(.A(G143), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n759), .A2(new_n812), .B1(new_n772), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n754), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n811), .B(new_n814), .C1(new_n769), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n748), .A2(G68), .ZN(new_n819));
  INV_X1    g0619(.A(G132), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n336), .B1(new_n751), .B2(new_n202), .C1(new_n820), .C2(new_n753), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G50), .B2(new_n777), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n818), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n809), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n808), .A2(KEYINPUT103), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n736), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n723), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n736), .A2(new_n737), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(new_n828), .B2(new_n284), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n643), .A2(new_n365), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n366), .B2(new_n370), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n358), .A2(new_n356), .A3(new_n365), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n830), .B1(new_n833), .B2(new_n354), .ZN(new_n834));
  OAI21_X1  g0634(.A(KEYINPUT104), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n358), .A2(new_n356), .A3(new_n365), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT71), .B1(new_n355), .B2(new_n302), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n370), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n830), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT104), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n366), .A2(new_n831), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n835), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n826), .B(new_n829), .C1(new_n843), .C2(new_n738), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n715), .B(new_n843), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n723), .B1(new_n845), .B2(new_n704), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n704), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n844), .B1(new_n847), .B2(new_n848), .ZN(G384));
  NOR2_X1   g0649(.A1(new_n720), .A2(new_n211), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT40), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n405), .A2(new_n408), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n402), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n641), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n444), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n412), .A2(new_n854), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n421), .A2(new_n858), .A3(new_n859), .A4(new_n439), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n853), .A2(new_n420), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n855), .A2(new_n861), .A3(new_n439), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n860), .B1(new_n862), .B2(new_n859), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n857), .A2(new_n863), .A3(KEYINPUT38), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n857), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT107), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n423), .A2(new_n434), .B1(new_n853), .B2(new_n420), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n859), .B1(new_n868), .B2(new_n855), .ZN(new_n869));
  INV_X1    g0669(.A(new_n860), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n855), .B1(new_n612), .B2(new_n608), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT107), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n857), .A2(new_n863), .A3(KEYINPUT38), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n866), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n681), .B1(new_n691), .B2(new_n695), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n878), .A2(new_n698), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT31), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n644), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n539), .A2(new_n568), .A3(new_n598), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n495), .B1(new_n497), .B2(new_n504), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n879), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(G169), .B1(new_n297), .B2(new_n298), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT14), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n270), .A2(new_n273), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n888), .A2(new_n307), .B1(new_n889), .B2(new_n303), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n310), .A2(new_n643), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n300), .B(new_n891), .C1(new_n890), .C2(new_n296), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT105), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT105), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n610), .A2(new_n895), .A3(new_n300), .A4(new_n891), .ZN(new_n896));
  AOI211_X1 g0696(.A(KEYINPUT106), .B(new_n892), .C1(new_n894), .C2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT106), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n894), .A2(new_n896), .ZN(new_n899));
  INV_X1    g0699(.A(new_n892), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n885), .B(new_n843), .C1(new_n897), .C2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n851), .B1(new_n877), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n858), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n444), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n421), .A2(new_n858), .A3(new_n439), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT37), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n860), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n867), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n875), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT40), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n903), .B1(new_n902), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT109), .ZN(new_n914));
  INV_X1    g0714(.A(new_n885), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n448), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n671), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n914), .B2(new_n916), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n644), .B(new_n843), .C1(new_n630), .C2(new_n635), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n366), .A2(new_n643), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n897), .B2(new_n901), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n877), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n905), .B2(new_n908), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(new_n864), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n873), .A2(KEYINPUT39), .A3(new_n875), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n309), .A2(new_n310), .A3(new_n644), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT108), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n929), .A2(new_n932), .B1(new_n608), .B2(new_n854), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n924), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n447), .B(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n615), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n934), .B(new_n936), .Z(new_n937));
  AOI21_X1  g0737(.A(new_n850), .B1(new_n918), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n937), .B2(new_n918), .ZN(new_n939));
  INV_X1    g0739(.A(new_n555), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n940), .A2(KEYINPUT35), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(KEYINPUT35), .ZN(new_n942));
  NOR4_X1   g0742(.A1(new_n941), .A2(new_n942), .A3(new_n475), .A4(new_n227), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT36), .Z(new_n944));
  NAND3_X1  g0744(.A1(new_n731), .A2(G77), .A3(new_n383), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n201), .A2(G68), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(G1), .A3(new_n275), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n939), .A2(new_n944), .A3(new_n948), .ZN(G367));
  AOI21_X1  g0749(.A(new_n651), .B1(new_n647), .B2(new_n649), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n567), .A2(new_n644), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT111), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n565), .A2(new_n643), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n706), .A2(new_n707), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT42), .ZN(new_n957));
  INV_X1    g0757(.A(new_n955), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n567), .B1(new_n958), .B2(new_n496), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n957), .B1(new_n644), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n577), .A2(new_n644), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n622), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n597), .B2(new_n961), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT110), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n960), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n960), .B2(new_n967), .ZN(new_n971));
  INV_X1    g0771(.A(new_n661), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n955), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n971), .B(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n665), .B(KEYINPUT41), .Z(new_n975));
  INV_X1    g0775(.A(new_n654), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(KEYINPUT44), .A3(new_n958), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n654), .B2(new_n955), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n654), .A2(new_n955), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n654), .A2(KEYINPUT45), .A3(new_n955), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n972), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n650), .A2(new_n652), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n988), .A2(new_n659), .A3(new_n950), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n659), .B1(new_n988), .B2(new_n950), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n991), .A2(new_n718), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n980), .A2(new_n985), .A3(new_n661), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n987), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT112), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n987), .A2(new_n992), .A3(KEYINPUT112), .A4(new_n993), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n975), .B1(new_n998), .B2(new_n718), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n974), .B1(new_n999), .B2(new_n722), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n768), .A2(new_n201), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n777), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n1002), .A2(new_n202), .B1(new_n284), .B2(new_n744), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n789), .A2(G68), .B1(G143), .B2(new_n758), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n754), .B2(new_n774), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n336), .B1(new_n753), .B2(new_n812), .C1(new_n772), .C2(new_n810), .ZN(new_n1006));
  NOR4_X1   g0806(.A1(new_n1001), .A2(new_n1003), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT113), .Z(new_n1008));
  NAND2_X1  g0808(.A1(new_n777), .A2(G116), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT46), .Z(new_n1010));
  OAI22_X1  g0810(.A1(new_n774), .A2(new_n452), .B1(new_n751), .B2(new_n206), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G311), .B2(new_n758), .ZN(new_n1012));
  INV_X1    g0812(.A(G317), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n345), .B1(new_n753), .B2(new_n1013), .C1(new_n772), .C2(new_n524), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n769), .B2(G283), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1012), .B(new_n1015), .C1(new_n205), .C2(new_n744), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1008), .B1(new_n1010), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT47), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n736), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n741), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n729), .A2(new_n239), .B1(new_n664), .B2(new_n591), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n827), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1019), .B(new_n1022), .C1(new_n797), .C2(new_n963), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1000), .A2(new_n1023), .ZN(G387));
  NOR2_X1   g0824(.A1(new_n992), .A2(new_n666), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n718), .B2(new_n991), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n650), .A2(new_n797), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n726), .A2(new_n667), .B1(G107), .B2(new_n215), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n236), .A2(new_n262), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n667), .ZN(new_n1030));
  AOI211_X1 g0830(.A(G45), .B(new_n1030), .C1(G68), .C2(G77), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n320), .A2(G50), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n730), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1028), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n723), .B1(new_n1035), .B2(new_n741), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n777), .A2(G77), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n810), .B2(new_n753), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT115), .Z(new_n1039));
  OAI221_X1 g0839(.A(new_n336), .B1(new_n387), .B2(new_n759), .C1(new_n768), .C2(new_n228), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n323), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1040), .B1(new_n1041), .B2(new_n773), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n789), .A2(new_n591), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n201), .B2(new_n772), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT116), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n748), .A2(G97), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1039), .A2(new_n1042), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n772), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1048), .A2(G317), .B1(G311), .B2(new_n773), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n781), .B2(new_n759), .C1(new_n768), .C2(new_n524), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n777), .A2(G294), .B1(G283), .B2(new_n789), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT49), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n345), .B1(new_n784), .B2(new_n753), .C1(new_n744), .C2(new_n475), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1047), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1036), .B1(new_n1061), .B2(new_n736), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT117), .ZN(new_n1063));
  AOI21_X1  g0863(.A(KEYINPUT114), .B1(new_n991), .B2(new_n722), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n991), .A2(KEYINPUT114), .A3(new_n722), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1026), .B1(new_n1027), .B2(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(G393));
  AOI21_X1  g0866(.A(new_n992), .B1(new_n987), .B2(new_n993), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n666), .B(new_n1067), .C1(new_n996), .C2(new_n997), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n987), .A2(new_n722), .A3(new_n993), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n759), .A2(new_n810), .B1(new_n772), .B2(new_n387), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT51), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n751), .A2(new_n284), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n336), .B1(new_n753), .B2(new_n813), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(G50), .C2(new_n773), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n769), .A2(new_n318), .B1(G68), .B2(new_n777), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n803), .A2(new_n1071), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n345), .B1(new_n753), .B2(new_n781), .C1(new_n774), .C2(new_n524), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G116), .B2(new_n789), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n769), .A2(G294), .B1(G283), .B2(new_n777), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n749), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1048), .A2(G311), .B1(G317), .B2(new_n758), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1076), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n736), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n729), .A2(new_n247), .B1(G97), .B2(new_n664), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n827), .B1(new_n1020), .B2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(new_n955), .C2(new_n797), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1069), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1068), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(G390));
  AOI21_X1  g0890(.A(new_n931), .B1(new_n910), .B2(new_n875), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n901), .A2(new_n897), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n843), .B(new_n644), .C1(new_n710), .C2(new_n713), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(new_n921), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n895), .B1(new_n311), .B2(new_n891), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n893), .A2(KEYINPUT105), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n900), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT106), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n899), .A2(new_n898), .A3(new_n900), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n703), .A2(new_n1101), .A3(new_n843), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n931), .B1(new_n1101), .B2(new_n922), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n927), .A2(new_n928), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1095), .B(new_n1102), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT118), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1099), .A2(new_n1100), .B1(new_n919), .B2(new_n921), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n929), .B1(new_n1107), .B2(new_n931), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT118), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n1095), .A4(new_n1102), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n885), .A2(G330), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n843), .B1(new_n901), .B2(new_n897), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n923), .A2(new_n932), .B1(new_n927), .B2(new_n928), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1095), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1106), .A2(new_n1110), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n929), .A2(new_n737), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n828), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n723), .B1(new_n1119), .B2(new_n1041), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n759), .A2(new_n793), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1072), .B(new_n1121), .C1(G107), .C2(new_n773), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n769), .A2(G97), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n345), .B1(new_n753), .B2(new_n452), .C1(new_n772), .C2(new_n475), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G87), .B2(new_n777), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n819), .A2(new_n1122), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n777), .A2(G150), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT53), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n774), .A2(new_n812), .B1(new_n751), .B2(new_n387), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G128), .B2(new_n758), .ZN(new_n1130));
  INV_X1    g0930(.A(G125), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n336), .B1(new_n753), .B2(new_n1131), .C1(new_n772), .C2(new_n820), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT54), .B(G143), .Z(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n769), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1130), .B(new_n1134), .C1(new_n201), .C2(new_n744), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1126), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1120), .B1(new_n1136), .B2(new_n736), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1117), .A2(new_n722), .B1(new_n1118), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1106), .A2(new_n1116), .A3(new_n1110), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1101), .B1(new_n703), .B2(new_n843), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n922), .B1(new_n1140), .B2(new_n1113), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n843), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1092), .B1(new_n1111), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n1094), .A3(new_n1102), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n671), .B1(new_n697), .B2(new_n879), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n447), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n615), .A2(new_n935), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n666), .B1(new_n1139), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT119), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1148), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1153), .A2(new_n1110), .A3(new_n1116), .A4(new_n1106), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1152), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1138), .B1(new_n1155), .B2(new_n1156), .ZN(G378));
  INV_X1    g0957(.A(KEYINPUT123), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n603), .A2(new_n604), .A3(new_n342), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n330), .A2(new_n854), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1160), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n605), .A2(new_n342), .A3(new_n1162), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n1168), .A3(new_n1159), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1112), .A2(new_n915), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n866), .A2(new_n876), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT40), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(G330), .B1(new_n902), .B2(new_n912), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1170), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n912), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n671), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n903), .A3(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1175), .A2(new_n934), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n934), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT57), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1148), .B(KEYINPUT122), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1117), .B2(new_n1153), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1158), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1175), .A2(new_n1179), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n934), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1175), .A2(new_n1179), .A3(new_n934), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1183), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1154), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1190), .A2(new_n1192), .A3(KEYINPUT123), .A4(KEYINPUT57), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1185), .A2(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1189), .A2(new_n1188), .B1(new_n1154), .B2(new_n1191), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n665), .B1(new_n1195), .B2(KEYINPUT57), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1190), .A2(new_n722), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n723), .B1(new_n1119), .B2(G50), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n336), .A2(G41), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G50), .B(new_n1200), .C1(new_n451), .C2(new_n261), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1037), .A2(new_n1200), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1202), .A2(KEYINPUT120), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n744), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n769), .A2(new_n591), .B1(new_n1204), .B2(G58), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n772), .A2(new_n206), .B1(new_n753), .B2(new_n793), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n774), .A2(new_n205), .B1(new_n759), .B2(new_n475), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G68), .C2(new_n789), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1202), .A2(KEYINPUT120), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1203), .A2(new_n1205), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT58), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1201), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n769), .A2(G137), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1048), .A2(G128), .B1(new_n789), .B2(G150), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G125), .A2(new_n758), .B1(new_n773), .B2(G132), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n777), .A2(new_n1133), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  INV_X1    g1018(.A(G124), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n451), .B(new_n261), .C1(new_n753), .C2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1204), .B2(new_n815), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1212), .B1(new_n1211), .B2(new_n1210), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1199), .B1(new_n1224), .B2(new_n736), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1178), .B2(new_n738), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT121), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1198), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1197), .A2(new_n1229), .ZN(G375));
  NOR2_X1   g1030(.A1(new_n1153), .A2(new_n975), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1149), .B2(new_n1145), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1092), .A2(new_n737), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n723), .B1(new_n1119), .B2(G68), .ZN(new_n1234));
  INV_X1    g1034(.A(G128), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n336), .B1(new_n753), .B2(new_n1235), .C1(new_n772), .C2(new_n812), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G58), .B2(new_n1204), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1237), .B1(new_n810), .B2(new_n768), .C1(new_n387), .C2(new_n1002), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1133), .A2(new_n773), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n201), .B2(new_n751), .C1(new_n759), .C2(new_n820), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1043), .B1(new_n759), .B2(new_n452), .C1(new_n475), .C2(new_n774), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n345), .B1(new_n753), .B2(new_n524), .C1(new_n772), .C2(new_n793), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G97), .B2(new_n777), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1242), .B(new_n1244), .C1(new_n206), .C2(new_n768), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n747), .A2(new_n284), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1238), .A2(new_n1240), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1234), .B1(new_n1247), .B2(new_n736), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT124), .Z(new_n1249));
  AOI22_X1  g1049(.A1(new_n1145), .A2(new_n722), .B1(new_n1233), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1232), .A2(new_n1250), .ZN(G381));
  NOR2_X1   g1051(.A1(G387), .A2(G390), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(KEYINPUT125), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(KEYINPUT125), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1257), .A2(new_n1138), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(G375), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1255), .A2(new_n1256), .A3(new_n1260), .ZN(G407));
  INV_X1    g1061(.A(G213), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1260), .B2(new_n642), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G407), .A2(new_n1263), .ZN(G409));
  INV_X1    g1064(.A(KEYINPUT126), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G378), .B(new_n1229), .C1(new_n1194), .C2(new_n1196), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1190), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1267), .A2(new_n975), .A3(new_n1184), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1258), .B1(new_n1268), .B2(new_n1228), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(KEYINPUT60), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1141), .A2(new_n1272), .A3(new_n1144), .A4(new_n1148), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1153), .A2(new_n666), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(G384), .A3(new_n1250), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1276), .B2(new_n1250), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1262), .A2(G343), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  AND4_X1   g1082(.A1(new_n1265), .A2(new_n1270), .A3(new_n1280), .A4(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1265), .B1(new_n1284), .B2(new_n1280), .ZN(new_n1285));
  OR3_X1    g1085(.A1(new_n1283), .A2(new_n1285), .A3(KEYINPUT63), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1089), .B1(new_n1000), .B2(new_n1023), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1252), .A2(new_n1287), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(G393), .B(new_n799), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1252), .A2(new_n1289), .A3(new_n1287), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  INV_X1    g1094(.A(G2897), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1282), .A2(new_n1295), .ZN(new_n1296));
  OR3_X1    g1096(.A1(new_n1278), .A2(new_n1279), .A3(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1294), .B1(new_n1284), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1284), .A2(KEYINPUT63), .A3(new_n1280), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1286), .A2(new_n1293), .A3(new_n1301), .A4(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1284), .B2(new_n1280), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1300), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1305), .A2(KEYINPUT127), .A3(new_n1307), .ZN(new_n1308));
  OR2_X1    g1108(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT127), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1303), .B1(new_n1310), .B2(new_n1311), .ZN(G405));
  AOI21_X1  g1112(.A(new_n1259), .B1(new_n1197), .B2(new_n1229), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1266), .ZN(new_n1314));
  OR3_X1    g1114(.A1(new_n1313), .A2(new_n1280), .A3(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1280), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1309), .B(new_n1317), .ZN(G402));
endmodule


