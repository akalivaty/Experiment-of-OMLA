//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G227), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT77), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT82), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT78), .A2(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT78), .A2(G107), .ZN(new_n195));
  AOI21_X1  g009(.A(G104), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G104), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(G101), .B1(new_n196), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  AOI21_X1  g016(.A(G101), .B1(new_n202), .B2(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n194), .A2(new_n195), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n202), .A2(KEYINPUT3), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n201), .B(new_n203), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  AOI21_X1  g025(.A(G128), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(KEYINPUT1), .A3(G146), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT67), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n216), .B(new_n213), .C1(new_n217), .C2(G128), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n220), .A3(G128), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n207), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n209), .A2(new_n211), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n225), .A3(new_n213), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n206), .A3(new_n200), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n222), .A2(KEYINPUT81), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT81), .B1(new_n222), .B2(new_n227), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT11), .A3(G134), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(G137), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  INV_X1    g051(.A(G131), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n232), .A2(new_n234), .A3(new_n238), .A4(new_n235), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n228), .A2(new_n229), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n193), .B1(new_n242), .B2(KEYINPUT12), .ZN(new_n243));
  INV_X1    g057(.A(new_n229), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n222), .A2(KEYINPUT81), .A3(new_n227), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n240), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT12), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(KEYINPUT82), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n222), .A2(new_n227), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n241), .A2(new_n247), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n243), .A2(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n201), .B1(new_n204), .B2(new_n205), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n197), .A2(G104), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n252), .B(G101), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT0), .A4(G128), .ZN(new_n256));
  OR2_X1    g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n256), .B(KEYINPUT64), .C1(new_n217), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT64), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n223), .A2(new_n261), .A3(new_n258), .A4(new_n257), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G101), .ZN(new_n264));
  AND2_X1   g078(.A1(KEYINPUT78), .A2(G107), .ZN(new_n265));
  NOR2_X1   g079(.A1(KEYINPUT78), .A2(G107), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n202), .A2(KEYINPUT3), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n267), .A2(new_n268), .B1(KEYINPUT3), .B2(new_n198), .ZN(new_n269));
  INV_X1    g083(.A(new_n254), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n206), .A2(KEYINPUT4), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n255), .B(new_n263), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n216), .B1(new_n225), .B2(new_n213), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n212), .A2(KEYINPUT67), .A3(new_n214), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n221), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n202), .B1(new_n265), .B2(new_n266), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n198), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n269), .A2(new_n203), .B1(new_n278), .B2(G101), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n276), .A2(KEYINPUT10), .A3(new_n279), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n281));
  NAND2_X1  g095(.A1(new_n227), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(KEYINPUT80), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT80), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(new_n227), .B2(new_n281), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n273), .B(new_n280), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(new_n240), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n192), .B1(new_n251), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n282), .B(KEYINPUT80), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n280), .A2(new_n273), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n241), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT83), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n191), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n286), .A2(new_n240), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n191), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT83), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n288), .A2(G469), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G469), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT72), .B(G902), .Z(new_n301));
  NAND2_X1  g115(.A1(new_n243), .A2(new_n248), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n249), .A2(new_n250), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n296), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n191), .B1(new_n294), .B2(new_n291), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n300), .B(new_n301), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(G469), .A2(G902), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n299), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G221), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT9), .B(G234), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT16), .ZN(new_n316));
  AND2_X1   g130(.A1(KEYINPUT74), .A2(G125), .ZN(new_n317));
  NOR2_X1   g131(.A1(KEYINPUT74), .A2(G125), .ZN(new_n318));
  OAI21_X1  g132(.A(G140), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(G125), .A2(G140), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n316), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT74), .B(G125), .ZN(new_n323));
  NOR2_X1   g137(.A1(KEYINPUT16), .A2(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n208), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n320), .B1(new_n323), .B2(G140), .ZN(new_n328));
  OAI211_X1 g142(.A(G146), .B(new_n325), .C1(new_n328), .C2(new_n316), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT92), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G237), .ZN(new_n333));
  AND4_X1   g147(.A1(G143), .A2(new_n333), .A3(new_n187), .A4(G214), .ZN(new_n334));
  NOR2_X1   g148(.A1(G237), .A2(G953), .ZN(new_n335));
  AOI21_X1  g149(.A(G143), .B1(new_n335), .B2(G214), .ZN(new_n336));
  OAI21_X1  g150(.A(G131), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n187), .A3(G214), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n210), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(G143), .A3(G214), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n238), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  MUX2_X1   g156(.A(new_n342), .B(new_n337), .S(KEYINPUT17), .Z(new_n343));
  NAND3_X1  g157(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT92), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n332), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G113), .B(G122), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(new_n202), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n319), .A2(G146), .A3(new_n321), .ZN(new_n348));
  XNOR2_X1  g162(.A(G125), .B(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n208), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g165(.A1(KEYINPUT18), .A2(G131), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n334), .A2(new_n336), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT89), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND4_X1   g169(.A1(new_n354), .A2(new_n339), .A3(new_n352), .A4(new_n340), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n345), .A2(new_n347), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n347), .B1(new_n345), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n312), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G475), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n328), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n319), .A2(KEYINPUT19), .A3(new_n321), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT19), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT90), .B1(new_n349), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(G146), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n329), .A2(new_n342), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n357), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT91), .ZN(new_n371));
  INV_X1    g185(.A(new_n347), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT91), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n357), .B(new_n373), .C1(new_n368), .C2(new_n369), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n345), .A2(new_n347), .A3(new_n357), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(G475), .A2(G902), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n362), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n378), .ZN(new_n380));
  AOI211_X1 g194(.A(KEYINPUT20), .B(new_n380), .C1(new_n375), .C2(new_n376), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n361), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT93), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n361), .B(KEYINPUT93), .C1(new_n379), .C2(new_n381), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G214), .B1(G237), .B2(G902), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G210), .B1(G237), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n263), .A2(new_n323), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n223), .A2(KEYINPUT1), .A3(new_n224), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n215), .B2(new_n218), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n393), .B2(new_n323), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n187), .A2(G224), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n394), .B(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT2), .ZN(new_n398));
  INV_X1    g212(.A(G113), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT69), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT69), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(KEYINPUT2), .B2(G113), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT2), .A2(G113), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT70), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT70), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT2), .A3(G113), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G116), .B(G119), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n403), .A2(new_n408), .A3(new_n410), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n414), .B(new_n255), .C1(new_n271), .C2(new_n272), .ZN(new_n415));
  XNOR2_X1  g229(.A(G110), .B(G122), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT86), .ZN(new_n417));
  INV_X1    g231(.A(G119), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G116), .ZN(new_n419));
  INV_X1    g233(.A(G116), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G119), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n421), .A3(KEYINPUT5), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT5), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(new_n418), .A3(G116), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n423), .A2(new_n418), .A3(KEYINPUT84), .A4(G116), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n422), .A2(new_n426), .A3(G113), .A4(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n428), .A2(new_n413), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT85), .B1(new_n429), .B2(new_n279), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n200), .A2(new_n428), .A3(new_n206), .A4(new_n413), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n415), .B(new_n417), .C1(new_n430), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT6), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n415), .B1(new_n430), .B2(new_n433), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n417), .B(KEYINPUT87), .Z(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n397), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT88), .A2(KEYINPUT7), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n394), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n395), .A2(KEYINPUT7), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n417), .B(KEYINPUT8), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n429), .A2(new_n279), .ZN(new_n447));
  INV_X1    g261(.A(new_n431), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n444), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n393), .A2(new_n323), .ZN(new_n451));
  INV_X1    g265(.A(new_n323), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(new_n260), .B2(new_n262), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n450), .B(new_n442), .C1(new_n451), .C2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n445), .A2(new_n434), .A3(new_n449), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n312), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n390), .B1(new_n441), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n397), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n434), .A2(KEYINPUT6), .B1(new_n436), .B2(new_n437), .ZN(new_n459));
  INV_X1    g273(.A(new_n440), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n454), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n450), .B1(new_n394), .B2(new_n442), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n434), .A2(new_n449), .ZN(new_n465));
  AOI21_X1  g279(.A(G902), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n461), .A2(new_n466), .A3(new_n389), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n388), .B1(new_n457), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT96), .B(G952), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(G953), .ZN(new_n470));
  NAND2_X1  g284(.A1(G234), .A2(G237), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n301), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(G953), .A3(new_n471), .ZN(new_n474));
  XOR2_X1   g288(.A(KEYINPUT21), .B(G898), .Z(new_n475));
  OAI21_X1  g289(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT94), .B1(new_n420), .B2(G122), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n478));
  INV_X1    g292(.A(G122), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n479), .A3(G116), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n420), .A2(G122), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n477), .A2(new_n480), .B1(new_n481), .B2(KEYINPUT14), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT95), .ZN(new_n483));
  OAI22_X1  g297(.A1(new_n482), .A2(new_n483), .B1(KEYINPUT14), .B2(new_n481), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n482), .A2(new_n483), .ZN(new_n485));
  OAI21_X1  g299(.A(G107), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n477), .A2(new_n480), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n267), .A3(new_n481), .ZN(new_n488));
  XNOR2_X1  g302(.A(G128), .B(G143), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n489), .A2(G134), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(G134), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n481), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n204), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n488), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT13), .B1(new_n224), .B2(G143), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(new_n231), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n489), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G217), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n310), .A2(new_n502), .A3(G953), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n486), .A2(new_n492), .B1(new_n496), .B2(new_n499), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n503), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n301), .ZN(new_n509));
  INV_X1    g323(.A(G478), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n509), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n386), .A2(new_n468), .A3(new_n476), .A4(new_n513), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n315), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G472), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT65), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n231), .B2(G137), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n233), .A2(G134), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n233), .A2(G134), .ZN(new_n521));
  OAI21_X1  g335(.A(G131), .B1(new_n521), .B2(new_n517), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT66), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT66), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n231), .A2(G137), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n238), .B1(new_n525), .B2(KEYINPUT65), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n521), .A2(new_n235), .A3(new_n517), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n239), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT68), .B1(new_n529), .B2(new_n393), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT68), .ZN(new_n531));
  INV_X1    g345(.A(new_n239), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT66), .B1(new_n520), .B2(new_n522), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n526), .A2(new_n524), .A3(new_n527), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n276), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n263), .A2(new_n240), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n530), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n537), .B(KEYINPUT30), .C1(new_n529), .C2(new_n393), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n414), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n276), .A2(new_n535), .ZN(new_n543));
  INV_X1    g357(.A(new_n414), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n537), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n335), .A2(G210), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n547), .B(KEYINPUT27), .Z(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT26), .B(G101), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n548), .B(new_n549), .Z(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT29), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT71), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n538), .A2(new_n553), .A3(new_n414), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n545), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n538), .B2(new_n414), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT28), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n545), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(KEYINPUT28), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n552), .B1(new_n561), .B2(new_n551), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n544), .B1(new_n543), .B2(new_n537), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n559), .B1(new_n564), .B2(KEYINPUT28), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n550), .A2(KEYINPUT29), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n473), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n516), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT32), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n561), .A2(new_n551), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n542), .A2(new_n545), .A3(new_n550), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT31), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n542), .A2(KEYINPUT31), .A3(new_n545), .A4(new_n550), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G472), .A2(G902), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n570), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n578), .ZN(new_n580));
  AOI211_X1 g394(.A(KEYINPUT32), .B(new_n580), .C1(new_n571), .C2(new_n576), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n569), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n502), .B1(new_n301), .B2(G234), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT22), .B(G137), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(G119), .B(G128), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT24), .B(G110), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT73), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT23), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n418), .B2(G128), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n595), .B(new_n596), .C1(G119), .C2(new_n224), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n597), .A2(G110), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n593), .A2(new_n598), .B1(new_n208), .B2(new_n349), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n589), .B(KEYINPUT73), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n600), .A2(new_n587), .B1(G110), .B2(new_n597), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n599), .A2(new_n329), .B1(new_n330), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n586), .B1(new_n602), .B2(KEYINPUT75), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n599), .A2(new_n329), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n330), .A2(new_n601), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT75), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n602), .A2(KEYINPUT75), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n603), .B1(new_n610), .B2(new_n586), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT25), .B1(new_n611), .B2(new_n301), .ZN(new_n612));
  INV_X1    g426(.A(new_n586), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n608), .B2(new_n609), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT25), .ZN(new_n615));
  NOR4_X1   g429(.A1(new_n614), .A2(new_n615), .A3(new_n473), .A4(new_n603), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n583), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n583), .A2(G902), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n582), .A2(KEYINPUT76), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT76), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n561), .A2(new_n551), .B1(new_n574), .B2(new_n575), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT32), .B1(new_n624), .B2(new_n580), .ZN(new_n625));
  INV_X1    g439(.A(new_n541), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n539), .B2(new_n538), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n558), .B1(new_n627), .B2(new_n414), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT31), .B1(new_n628), .B2(new_n550), .ZN(new_n629));
  INV_X1    g443(.A(new_n575), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n550), .B1(new_n557), .B2(new_n560), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n570), .B(new_n578), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n568), .B1(new_n625), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n623), .B1(new_n634), .B2(new_n620), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n515), .B1(new_n622), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n264), .ZN(G3));
  AOI21_X1  g451(.A(new_n473), .B1(new_n571), .B2(new_n576), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n638), .A2(KEYINPUT97), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n516), .B1(new_n638), .B2(KEYINPUT97), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n639), .A2(new_n640), .B1(new_n578), .B2(new_n577), .ZN(new_n641));
  INV_X1    g455(.A(new_n315), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n641), .A2(new_n642), .A3(new_n621), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(KEYINPUT98), .Z(new_n644));
  NOR2_X1   g458(.A1(new_n473), .A2(new_n510), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT33), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n505), .A2(new_n646), .A3(new_n507), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n646), .B1(new_n505), .B2(new_n507), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT99), .B(G478), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n508), .B2(new_n301), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n650), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n645), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n506), .A2(new_n503), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n493), .A2(new_n500), .A3(new_n503), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT33), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n656), .B1(new_n659), .B2(new_n647), .ZN(new_n660));
  OAI21_X1  g474(.A(KEYINPUT100), .B1(new_n660), .B2(new_n653), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n384), .A2(new_n662), .A3(new_n385), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n468), .A2(new_n476), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n644), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT101), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  NOR3_X1   g483(.A1(new_n664), .A2(new_n513), .A3(new_n382), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n644), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NOR2_X1   g487(.A1(new_n315), .A2(new_n514), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n613), .A2(KEYINPUT36), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n606), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n618), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n617), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n674), .A2(new_n641), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT37), .B(G110), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n468), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n582), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n472), .B1(new_n474), .B2(G900), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n513), .A2(new_n382), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n308), .A2(new_n314), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n682), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n625), .A2(new_n633), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n683), .B1(new_n691), .B2(new_n569), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n308), .A2(new_n314), .A3(new_n688), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(KEYINPUT102), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  XNOR2_X1  g510(.A(new_n686), .B(KEYINPUT39), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n642), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT40), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n642), .A2(new_n700), .A3(new_n697), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n564), .A2(new_n551), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT103), .ZN(new_n703));
  INV_X1    g517(.A(new_n572), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n312), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G472), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n691), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n678), .A2(new_n388), .A3(new_n513), .ZN(new_n708));
  INV_X1    g522(.A(new_n457), .ZN(new_n709));
  INV_X1    g523(.A(new_n467), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT38), .ZN(new_n712));
  INV_X1    g526(.A(new_n386), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(KEYINPUT38), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n708), .A2(new_n712), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n699), .A2(new_n701), .A3(new_n707), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G143), .ZN(G45));
  AND4_X1   g532(.A1(new_n384), .A2(new_n662), .A3(new_n385), .A4(new_n686), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n719), .A2(new_n314), .A3(new_n308), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n692), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G146), .ZN(G48));
  NOR3_X1   g536(.A1(new_n242), .A2(new_n193), .A3(KEYINPUT12), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT82), .B1(new_n246), .B2(new_n247), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n303), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n296), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n305), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(G469), .B1(new_n727), .B2(new_n473), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n728), .A2(new_n314), .A3(new_n306), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n582), .A2(new_n621), .A3(new_n665), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND4_X1  g546(.A1(new_n582), .A2(new_n621), .A3(new_n670), .A4(new_n729), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  NAND4_X1  g548(.A1(new_n386), .A2(new_n678), .A3(new_n476), .A4(new_n513), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n728), .A2(new_n314), .A3(new_n306), .A4(new_n468), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(new_n582), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n634), .A2(new_n735), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(KEYINPUT104), .A3(new_n738), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  NOR3_X1   g559(.A1(new_n664), .A2(new_n386), .A3(new_n513), .ZN(new_n746));
  INV_X1    g560(.A(new_n638), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n576), .B1(new_n550), .B2(new_n565), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n747), .A2(G472), .B1(new_n578), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n746), .A2(new_n749), .A3(new_n621), .A4(new_n729), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  NOR2_X1   g565(.A1(new_n565), .A2(new_n550), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n578), .B1(new_n631), .B2(new_n752), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(new_n678), .C1(new_n638), .C2(new_n516), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n384), .A2(new_n662), .A3(new_n385), .A4(new_n686), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n738), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  NOR2_X1   g572(.A1(new_n634), .A2(new_n620), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n457), .A2(new_n387), .A3(new_n467), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n457), .A2(new_n467), .A3(KEYINPUT106), .A4(new_n387), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n762), .A2(new_n314), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n307), .B(KEYINPUT105), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n299), .A2(new_n306), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT107), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n299), .A2(new_n306), .A3(new_n765), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n762), .A2(new_n314), .A3(new_n763), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n759), .B(new_n719), .C1(new_n767), .C2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n764), .A2(KEYINPUT107), .A3(new_n766), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n770), .B1(new_n768), .B2(new_n769), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(KEYINPUT42), .A3(new_n759), .A4(new_n719), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G131), .ZN(G33));
  OAI211_X1 g594(.A(new_n759), .B(new_n688), .C1(new_n767), .C2(new_n771), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT108), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n777), .A2(new_n783), .A3(new_n759), .A4(new_n688), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  AOI21_X1  g600(.A(KEYINPUT45), .B1(new_n288), .B2(new_n298), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT109), .B1(new_n787), .B2(new_n300), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n725), .A2(new_n291), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n790), .A2(new_n192), .B1(new_n295), .B2(new_n297), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n789), .B(G469), .C1(new_n791), .C2(KEYINPUT45), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(KEYINPUT45), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n788), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT46), .B1(new_n794), .B2(new_n765), .ZN(new_n795));
  INV_X1    g609(.A(new_n306), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n765), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n313), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n386), .A2(new_n662), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT43), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT43), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n386), .A2(new_n803), .A3(new_n662), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n678), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n800), .B1(new_n805), .B2(new_n641), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT110), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n808), .B(new_n800), .C1(new_n805), .C2(new_n641), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n762), .A2(new_n763), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n805), .A2(new_n641), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n811), .B1(new_n812), .B2(KEYINPUT44), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n799), .A2(new_n810), .A3(new_n697), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  INV_X1    g629(.A(new_n811), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n620), .A3(new_n719), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n582), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n799), .A2(KEYINPUT47), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT47), .ZN(new_n821));
  INV_X1    g635(.A(new_n798), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n796), .A3(new_n795), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n823), .B2(new_n313), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n819), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(G140), .Z(G42));
  NAND2_X1  g640(.A1(new_n712), .A2(new_n714), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n314), .A3(new_n387), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n728), .A2(new_n306), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n801), .B(new_n828), .C1(KEYINPUT49), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n707), .A2(new_n620), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n830), .B(new_n831), .C1(KEYINPUT49), .C2(new_n829), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n756), .B1(new_n767), .B2(new_n771), .ZN(new_n834));
  INV_X1    g648(.A(new_n678), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n513), .A2(new_n686), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n811), .A2(new_n835), .A3(new_n382), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n642), .A3(new_n582), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n833), .B(new_n839), .C1(new_n784), .C2(new_n782), .ZN(new_n840));
  INV_X1    g654(.A(new_n839), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT111), .B1(new_n785), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n692), .A2(new_n720), .B1(new_n756), .B2(new_n738), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n713), .A2(new_n468), .A3(new_n512), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n314), .A2(new_n617), .A3(new_n677), .A4(new_n686), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n847), .A2(new_n766), .A3(KEYINPUT112), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT112), .B1(new_n847), .B2(new_n766), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n707), .B(new_n846), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n689), .A2(new_n634), .A3(new_n682), .A4(new_n683), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT102), .B1(new_n692), .B2(new_n693), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n844), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n695), .A2(KEYINPUT52), .A3(new_n844), .A4(new_n850), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT104), .B1(new_n742), .B2(new_n738), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n634), .A2(new_n735), .A3(new_n737), .A4(new_n740), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n386), .A2(new_n662), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n512), .B1(new_n384), .B2(new_n385), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n861), .A2(new_n862), .A3(new_n664), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n641), .A2(new_n863), .A3(new_n642), .A4(new_n621), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n679), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n730), .A2(new_n733), .A3(new_n750), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n860), .A2(new_n865), .A3(new_n636), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n857), .A2(new_n867), .A3(new_n779), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n843), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n866), .B1(new_n741), .B2(new_n743), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n865), .A2(new_n636), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n779), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n855), .B2(new_n856), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n582), .A2(new_n621), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n776), .B2(new_n775), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n783), .B1(new_n876), .B2(new_n688), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n783), .A2(new_n777), .A3(new_n759), .A4(new_n688), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n841), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n833), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n785), .A2(KEYINPUT111), .A3(new_n841), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT53), .B1(new_n874), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT54), .B1(new_n870), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n869), .B1(new_n843), .B2(new_n868), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT76), .B1(new_n582), .B2(new_n621), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n634), .A2(new_n623), .A3(new_n620), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n674), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(KEYINPUT53), .A3(new_n679), .A4(new_n864), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n774), .B2(new_n778), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT113), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n860), .B2(new_n866), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n730), .A2(new_n733), .A3(new_n750), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(new_n744), .A3(KEYINPUT113), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n890), .A2(new_n857), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n882), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n885), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n884), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT114), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n729), .A2(new_n901), .A3(new_n816), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n728), .A2(new_n314), .A3(new_n306), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT114), .B1(new_n903), .B2(new_n811), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n472), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n802), .A2(new_n804), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n908), .A2(new_n909), .A3(new_n754), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n909), .B1(new_n908), .B2(new_n754), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n905), .A2(new_n906), .A3(new_n831), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n713), .A2(new_n662), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n910), .A2(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND4_X1   g730(.A1(new_n906), .A2(new_n907), .A3(new_n621), .A4(new_n749), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n820), .A2(new_n824), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n829), .A2(new_n314), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n816), .B(new_n917), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT51), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n914), .B2(new_n915), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n827), .A2(new_n388), .A3(new_n729), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT50), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n916), .A2(new_n920), .A3(new_n922), .A4(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n908), .A2(new_n875), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT48), .Z(new_n930));
  NAND3_X1  g744(.A1(new_n912), .A2(new_n713), .A3(new_n662), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n917), .A2(new_n738), .ZN(new_n932));
  AND4_X1   g746(.A1(new_n470), .A2(new_n930), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n920), .A2(new_n914), .A3(new_n927), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n928), .B(new_n933), .C1(new_n934), .C2(KEYINPUT51), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n900), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(G952), .A2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n832), .B1(new_n936), .B2(new_n937), .ZN(G75));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n439), .A2(new_n440), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT117), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT55), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n397), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n874), .A2(new_n882), .ZN(new_n945));
  AOI22_X1  g759(.A1(new_n945), .A2(new_n869), .B1(new_n896), .B2(new_n882), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n301), .A2(new_n389), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n939), .B(new_n944), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n187), .A2(G952), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n948), .B1(new_n885), .B2(new_n897), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n943), .B1(new_n953), .B2(KEYINPUT56), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT118), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(KEYINPUT118), .B(new_n943), .C1(new_n953), .C2(KEYINPUT56), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(G51));
  XOR2_X1   g772(.A(new_n765), .B(KEYINPUT57), .Z(new_n959));
  NAND3_X1  g773(.A1(new_n890), .A2(new_n857), .A3(new_n895), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n843), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n883), .A2(new_n961), .A3(KEYINPUT54), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n898), .B1(new_n885), .B2(new_n897), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n727), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OR3_X1    g780(.A1(new_n946), .A2(new_n301), .A3(new_n794), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n950), .B1(new_n966), .B2(new_n967), .ZN(G54));
  NAND2_X1  g782(.A1(new_n885), .A2(new_n897), .ZN(new_n969));
  AND2_X1   g783(.A1(KEYINPUT58), .A2(G475), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n473), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n971), .A2(new_n376), .A3(new_n375), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n969), .A2(new_n473), .A3(new_n377), .A4(new_n970), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n972), .A2(new_n951), .A3(new_n973), .ZN(G60));
  NOR2_X1   g788(.A1(new_n648), .A2(new_n649), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  XOR2_X1   g790(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n977));
  NOR2_X1   g791(.A1(new_n510), .A2(new_n312), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n900), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n976), .A2(new_n979), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n962), .B2(new_n963), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n951), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n980), .A2(new_n983), .ZN(G63));
  INV_X1    g798(.A(KEYINPUT61), .ZN(new_n985));
  NAND2_X1  g799(.A1(G217), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT120), .Z(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT60), .Z(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n885), .B2(new_n897), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n611), .B(KEYINPUT121), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n951), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n969), .A2(new_n676), .A3(new_n988), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n985), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n991), .B1(new_n946), .B2(new_n989), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n990), .A2(new_n676), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n996), .A2(new_n997), .A3(KEYINPUT61), .A4(new_n951), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(G66));
  AOI21_X1  g813(.A(new_n187), .B1(new_n475), .B2(G224), .ZN(new_n1000));
  INV_X1    g814(.A(new_n867), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(new_n187), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n941), .B1(G898), .B2(new_n187), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT122), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1002), .B(new_n1004), .ZN(G69));
  NAND2_X1  g819(.A1(G227), .A2(G900), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n875), .A2(new_n845), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n799), .A2(new_n697), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n844), .B1(new_n851), .B2(new_n852), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(new_n774), .B2(new_n778), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n814), .A2(new_n785), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n187), .B1(new_n1011), .B2(new_n825), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n187), .A2(G900), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT124), .Z(new_n1014));
  NAND2_X1  g828(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(KEYINPUT125), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT125), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1012), .A2(new_n1017), .A3(new_n1014), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n363), .A2(new_n367), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n627), .B(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  OAI211_X1 g836(.A(G953), .B(new_n1006), .C1(new_n1019), .C2(new_n1022), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n1012), .A2(new_n1017), .A3(new_n1014), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1017), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1006), .A2(G953), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n717), .A2(new_n695), .A3(new_n844), .ZN(new_n1028));
  OR3_X1    g842(.A1(new_n1028), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1029));
  OAI21_X1  g843(.A(KEYINPUT123), .B1(new_n1028), .B2(KEYINPUT62), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(new_n825), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n622), .A2(new_n635), .ZN(new_n1033));
  NOR4_X1   g847(.A1(new_n698), .A2(new_n862), .A3(new_n811), .A4(new_n861), .ZN(new_n1034));
  AOI22_X1  g848(.A1(new_n1028), .A2(KEYINPUT62), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1031), .A2(new_n1032), .A3(new_n814), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1022), .B1(new_n1037), .B2(G953), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1026), .A2(new_n1027), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1023), .A2(new_n1039), .ZN(G72));
  NAND2_X1  g854(.A1(G472), .A2(G902), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT63), .Z(new_n1042));
  OAI21_X1  g856(.A(new_n1042), .B1(new_n1036), .B2(new_n1001), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n546), .B(KEYINPUT126), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n1044), .A2(new_n551), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n546), .A2(new_n551), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1047), .A2(new_n572), .ZN(new_n1048));
  OAI211_X1 g862(.A(new_n1042), .B(new_n1048), .C1(new_n870), .C2(new_n883), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1046), .A2(new_n951), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1044), .A2(new_n551), .ZN(new_n1051));
  OR2_X1    g865(.A1(new_n1011), .A2(new_n825), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1042), .B1(new_n1052), .B2(new_n1001), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1053), .A2(KEYINPUT127), .ZN(new_n1054));
  INV_X1    g868(.A(KEYINPUT127), .ZN(new_n1055));
  OAI211_X1 g869(.A(new_n1055), .B(new_n1042), .C1(new_n1052), .C2(new_n1001), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1051), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n1050), .A2(new_n1057), .ZN(G57));
endmodule


