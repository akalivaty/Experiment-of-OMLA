//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  NOR3_X1   g002(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT27), .B(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(KEYINPUT28), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT28), .B1(new_n209), .B2(new_n210), .ZN(new_n213));
  OAI221_X1 g012(.A(new_n203), .B1(new_n204), .B2(new_n208), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n216), .B1(new_n203), .B2(KEYINPUT65), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n218));
  AOI211_X1 g017(.A(new_n215), .B(new_n217), .C1(new_n218), .C2(KEYINPUT65), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n205), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT25), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n203), .A2(new_n216), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n224), .A2(new_n218), .A3(new_n215), .ZN(new_n225));
  OR3_X1    g024(.A1(new_n222), .A2(new_n225), .A3(KEYINPUT25), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n214), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G113gat), .B(G120gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  XOR2_X1   g028(.A(G127gat), .B(G134gat), .Z(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n227), .A2(new_n232), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n237), .B(KEYINPUT64), .Z(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n233), .B2(new_n234), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT66), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT32), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n240), .A2(new_n242), .B1(new_n243), .B2(KEYINPUT33), .ZN(new_n244));
  XNOR2_X1  g043(.A(G71gat), .B(G99gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XNOR2_X1  g045(.A(G15gat), .B(G43gat), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n246), .B(new_n247), .Z(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n202), .B1(new_n244), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(KEYINPUT33), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n241), .A2(KEYINPUT66), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n241), .A2(KEYINPUT66), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(KEYINPUT68), .A3(new_n248), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n248), .A2(KEYINPUT33), .ZN(new_n257));
  OAI211_X1 g056(.A(KEYINPUT32), .B(new_n257), .C1(new_n252), .C2(new_n253), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n239), .A2(KEYINPUT34), .ZN(new_n261));
  OR3_X1    g060(.A1(new_n235), .A2(KEYINPUT70), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n237), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT34), .B1(new_n235), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT70), .B1(new_n235), .B2(new_n261), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n260), .B1(new_n266), .B2(KEYINPUT71), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n258), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n269), .B1(new_n250), .B2(new_n255), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT71), .B1(new_n270), .B2(new_n260), .ZN(new_n271));
  INV_X1    g070(.A(new_n266), .ZN(new_n272));
  OAI211_X1 g071(.A(KEYINPUT36), .B(new_n268), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n259), .A2(new_n266), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT36), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n270), .A2(new_n272), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279));
  INV_X1    g078(.A(G155gat), .ZN(new_n280));
  INV_X1    g079(.A(G162gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G141gat), .B(G148gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT74), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT75), .B(KEYINPUT2), .Z(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n283), .A2(KEYINPUT74), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n279), .B(new_n282), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT76), .ZN(new_n289));
  OR3_X1    g088(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n283), .A2(new_n289), .B1(new_n290), .B2(new_n279), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(new_n289), .B2(new_n283), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G197gat), .B(G204gat), .ZN(new_n294));
  AND2_X1   g093(.A1(G211gat), .A2(G218gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n294), .B1(KEYINPUT22), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G211gat), .B(G218gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT29), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n299), .A2(KEYINPUT81), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT3), .B1(new_n299), .B2(KEYINPUT81), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n293), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n292), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n305));
  XOR2_X1   g104(.A(KEYINPUT73), .B(KEYINPUT29), .Z(new_n306));
  OAI21_X1  g105(.A(new_n298), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G228gat), .ZN(new_n308));
  INV_X1    g107(.A(G233gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n303), .A2(new_n307), .A3(KEYINPUT82), .A4(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT82), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(new_n310), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(new_n302), .ZN(new_n314));
  INV_X1    g113(.A(new_n307), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n304), .A2(KEYINPUT77), .ZN(new_n316));
  INV_X1    g115(.A(new_n298), .ZN(new_n317));
  INV_X1    g116(.A(new_n306), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT3), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT77), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  OAI22_X1  g120(.A1(new_n315), .A2(new_n321), .B1(new_n308), .B2(new_n309), .ZN(new_n322));
  INV_X1    g121(.A(G22gat), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n311), .A2(new_n314), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT83), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n311), .A2(new_n314), .A3(new_n322), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G22gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT80), .B(G50gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT31), .ZN(new_n329));
  XOR2_X1   g128(.A(G78gat), .B(G106gat), .Z(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  AND4_X1   g130(.A1(new_n324), .A2(new_n325), .A3(new_n327), .A4(new_n331), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n325), .A2(new_n331), .B1(new_n327), .B2(new_n324), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335));
  INV_X1    g134(.A(G85gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  OAI21_X1  g138(.A(new_n231), .B1(new_n316), .B2(new_n320), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n305), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n232), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n293), .A2(new_n231), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(KEYINPUT5), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n304), .A2(new_n232), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n346), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n350), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT5), .ZN(new_n357));
  OAI211_X1 g156(.A(KEYINPUT4), .B(new_n231), .C1(new_n316), .C2(new_n320), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n350), .B1(new_n346), .B2(new_n341), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n345), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n358), .A2(new_n345), .A3(KEYINPUT78), .A4(new_n359), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n357), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n339), .B1(new_n353), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n364), .ZN(new_n366));
  INV_X1    g165(.A(new_n339), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n352), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(KEYINPUT6), .B(new_n339), .C1(new_n353), .C2(new_n364), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT79), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n352), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT6), .A4(new_n339), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n377), .B(KEYINPUT72), .Z(new_n378));
  NAND2_X1  g177(.A1(new_n227), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n227), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n317), .B(new_n379), .C1(new_n381), .C2(new_n378), .ZN(new_n382));
  INV_X1    g181(.A(new_n379), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n378), .B1(new_n227), .B2(new_n318), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n298), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT30), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n393), .B1(new_n386), .B2(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n387), .A2(new_n393), .A3(new_n391), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n334), .B1(new_n376), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT84), .B1(new_n278), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n376), .A2(new_n397), .ZN(new_n400));
  INV_X1    g199(.A(new_n334), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n402), .A2(new_n403), .A3(new_n277), .A4(new_n273), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n348), .A2(new_n349), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT39), .B1(new_n355), .B2(new_n350), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n406), .B(KEYINPUT85), .Z(new_n407));
  NOR2_X1   g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(KEYINPUT40), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n350), .B1(new_n342), .B2(new_n347), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n367), .B1(new_n411), .B2(KEYINPUT39), .ZN(new_n412));
  OR3_X1    g211(.A1(new_n408), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n397), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n410), .B1(new_n408), .B2(new_n412), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n413), .A2(new_n365), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT37), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n391), .B1(new_n387), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT38), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n298), .B(new_n379), .C1(new_n381), .C2(new_n378), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n317), .B1(new_n383), .B2(new_n384), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT37), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n386), .A2(KEYINPUT37), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n392), .B(new_n423), .C1(new_n425), .C2(new_n419), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n416), .B(new_n334), .C1(new_n376), .C2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n399), .A2(new_n404), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n270), .A2(new_n260), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT71), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n272), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n268), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n334), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT35), .B1(new_n433), .B2(new_n400), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n274), .A2(new_n276), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(new_n401), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n400), .A2(KEYINPUT87), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT35), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n376), .A2(new_n439), .A3(new_n397), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n436), .A2(new_n437), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n428), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(G1gat), .ZN(new_n444));
  INV_X1    g243(.A(G15gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n323), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n447));
  NAND2_X1  g246(.A1(G15gat), .A2(G22gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n444), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G8gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n446), .A2(new_n448), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT90), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n444), .A2(KEYINPUT16), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n449), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n453), .B1(new_n452), .B2(new_n457), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT21), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT9), .ZN(new_n463));
  INV_X1    g262(.A(G64gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G57gat), .ZN(new_n465));
  INV_X1    g264(.A(G57gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(G64gat), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g267(.A1(G71gat), .A2(G78gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(G71gat), .A2(G78gat), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT92), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n469), .A2(new_n470), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT92), .ZN(new_n474));
  XNOR2_X1  g273(.A(G57gat), .B(G64gat), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n463), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT93), .ZN(new_n478));
  INV_X1    g277(.A(new_n469), .ZN(new_n479));
  INV_X1    g278(.A(G71gat), .ZN(new_n480));
  INV_X1    g279(.A(G78gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT9), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n475), .A2(new_n478), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n478), .B2(new_n475), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n461), .B1(new_n462), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(G231gat), .A2(G233gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n462), .ZN(new_n491));
  XOR2_X1   g290(.A(G127gat), .B(G155gat), .Z(new_n492));
  XOR2_X1   g291(.A(new_n491), .B(new_n492), .Z(new_n493));
  XNOR2_X1  g292(.A(new_n490), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G183gat), .B(G211gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n495), .B(new_n496), .Z(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n493), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n490), .B(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n497), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G230gat), .A2(G233gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT99), .ZN(new_n507));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT8), .ZN(new_n509));
  NAND2_X1  g308(.A1(G85gat), .A2(G92gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n514));
  AND4_X1   g313(.A1(new_n509), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT97), .ZN(new_n516));
  AND2_X1   g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G99gat), .ZN(new_n520));
  INV_X1    g319(.A(G106gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(KEYINPUT97), .A3(new_n508), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n515), .A2(new_n524), .A3(KEYINPUT98), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT98), .B1(new_n515), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n507), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT98), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n519), .A2(new_n523), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n509), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n524), .A3(KEYINPUT98), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(KEYINPUT99), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n530), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n527), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n485), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT10), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT101), .B1(new_n515), .B2(new_n524), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT101), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n530), .A2(new_n539), .A3(new_n519), .A4(new_n523), .ZN(new_n540));
  AND4_X1   g339(.A1(new_n477), .A2(new_n538), .A3(new_n484), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n531), .A2(new_n532), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n536), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n527), .A2(new_n533), .A3(new_n534), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n545), .A2(KEYINPUT10), .A3(new_n477), .A4(new_n484), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n506), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n505), .B1(new_n536), .B2(new_n543), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G120gat), .B(G148gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(G176gat), .B(G204gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n549), .A2(new_n553), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G197gat), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT11), .B(G169gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT12), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(G29gat), .A2(G36gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT14), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n567), .A2(new_n568), .B1(G29gat), .B2(G36gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(G43gat), .B(G50gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT15), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT88), .B1(new_n570), .B2(KEYINPUT15), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT88), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT15), .ZN(new_n575));
  INV_X1    g374(.A(G43gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n576), .A2(G50gat), .ZN(new_n577));
  INV_X1    g376(.A(G50gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(G43gat), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n574), .B(new_n575), .C1(new_n577), .C2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n573), .A2(new_n569), .A3(new_n580), .A4(new_n571), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n572), .B1(new_n581), .B2(KEYINPUT89), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n569), .A2(new_n571), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT89), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n580), .A4(new_n573), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n455), .A2(new_n456), .A3(new_n449), .ZN(new_n587));
  AOI21_X1  g386(.A(G1gat), .B1(new_n455), .B2(new_n449), .ZN(new_n588));
  OAI21_X1  g387(.A(G8gat), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n458), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(new_n585), .A3(KEYINPUT17), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n461), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT17), .B1(new_n582), .B2(new_n585), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n564), .B(new_n591), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT18), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n564), .B(KEYINPUT13), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n591), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n586), .A2(new_n590), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(new_n595), .B2(new_n596), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n563), .B1(new_n598), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n597), .A2(KEYINPUT91), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT91), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n595), .A2(new_n607), .A3(new_n596), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n603), .B(new_n562), .C1(new_n595), .C2(new_n596), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n557), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT17), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n586), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(new_n592), .A3(new_n535), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n545), .A2(new_n586), .ZN(new_n616));
  NAND3_X1  g415(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G162gat), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT96), .B(G134gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT100), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n620), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n620), .A2(new_n621), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n627), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n504), .A2(new_n612), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n443), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n376), .A2(KEYINPUT102), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n370), .A2(new_n375), .A3(new_n372), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g438(.A1(new_n633), .A2(new_n414), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT42), .B1(new_n640), .B2(new_n453), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT16), .B(G8gat), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  MUX2_X1   g442(.A(KEYINPUT42), .B(new_n641), .S(new_n643), .Z(G1325gat));
  INV_X1    g443(.A(new_n435), .ZN(new_n645));
  AOI21_X1  g444(.A(G15gat), .B1(new_n633), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n278), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n445), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n633), .B2(new_n648), .ZN(G1326gat));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n401), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT43), .B(G22gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  NOR2_X1   g451(.A1(new_n503), .A2(new_n612), .ZN(new_n653));
  INV_X1    g452(.A(new_n637), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(G29gat), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n443), .A2(new_n631), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT45), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n443), .A2(KEYINPUT44), .A3(new_n631), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n278), .A2(new_n398), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n434), .A2(new_n441), .B1(new_n660), .B2(new_n427), .ZN(new_n661));
  MUX2_X1   g460(.A(new_n626), .B(new_n630), .S(new_n628), .Z(new_n662));
  OAI21_X1  g461(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n498), .A2(new_n502), .A3(KEYINPUT103), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT103), .B1(new_n498), .B2(new_n502), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n664), .A2(new_n665), .A3(new_n612), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n658), .A2(new_n663), .A3(new_n637), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(G29gat), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n657), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT104), .ZN(G1328gat));
  AND3_X1   g469(.A1(new_n443), .A2(new_n631), .A3(new_n653), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n397), .A2(G36gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT46), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n658), .A2(new_n663), .A3(new_n414), .A4(new_n666), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G36gat), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n671), .A2(new_n677), .A3(new_n672), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT105), .ZN(G1329gat));
  NAND2_X1  g479(.A1(new_n671), .A2(new_n645), .ZN(new_n681));
  AOI22_X1  g480(.A1(new_n681), .A2(new_n576), .B1(KEYINPUT106), .B2(KEYINPUT47), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n658), .A2(new_n663), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n683), .A2(G43gat), .A3(new_n278), .A4(new_n666), .ZN(new_n684));
  OR2_X1    g483(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n682), .B2(new_n684), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(G1330gat));
  NAND4_X1  g487(.A1(new_n658), .A2(new_n663), .A3(new_n401), .A4(new_n666), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G50gat), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(KEYINPUT48), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n334), .A2(G50gat), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n671), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(KEYINPUT48), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1331gat));
  NAND2_X1  g496(.A1(new_n660), .A2(new_n427), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n442), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n611), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n503), .A2(new_n700), .A3(new_n662), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n557), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n699), .A2(KEYINPUT108), .A3(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n654), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(new_n466), .ZN(G1332gat));
  AND2_X1   g508(.A1(new_n705), .A2(new_n706), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT111), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n397), .B(KEYINPUT109), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT49), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(new_n464), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT110), .Z(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n710), .A2(new_n711), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT111), .B1(new_n707), .B2(new_n716), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n718), .A2(new_n714), .A3(new_n719), .A4(new_n464), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1333gat));
  NAND3_X1  g522(.A1(new_n710), .A2(new_n480), .A3(new_n645), .ZN(new_n724));
  OAI21_X1  g523(.A(G71gat), .B1(new_n707), .B2(new_n647), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n724), .B2(new_n725), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(G1334gat));
  NOR2_X1   g528(.A1(new_n707), .A2(new_n334), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(new_n481), .ZN(G1335gat));
  NOR3_X1   g530(.A1(new_n503), .A2(new_n611), .A3(new_n557), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n683), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n654), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n503), .A2(new_n611), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n699), .A2(new_n631), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n699), .A2(KEYINPUT51), .A3(new_n631), .A4(new_n735), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n557), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(new_n336), .A3(new_n637), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n734), .A2(new_n741), .ZN(G1336gat));
  NOR2_X1   g541(.A1(new_n712), .A2(G92gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n740), .A2(KEYINPUT113), .A3(new_n743), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n658), .A2(new_n663), .A3(new_n713), .A4(new_n732), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G92gat), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n658), .A2(new_n663), .A3(new_n414), .A4(new_n732), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G92gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n744), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT52), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n755), .ZN(G1337gat));
  OAI21_X1  g555(.A(G99gat), .B1(new_n733), .B2(new_n647), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n520), .A3(new_n645), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1338gat));
  NAND4_X1  g558(.A1(new_n658), .A2(new_n663), .A3(new_n401), .A4(new_n732), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(G106gat), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n334), .A2(G106gat), .A3(new_n557), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT115), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n738), .B2(new_n739), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n765));
  OR3_X1    g564(.A1(new_n761), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n760), .A2(KEYINPUT114), .A3(G106gat), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT114), .B1(new_n760), .B2(G106gat), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n767), .A2(new_n768), .A3(new_n764), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(G1339gat));
  INV_X1    g570(.A(new_n557), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n701), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n664), .A2(new_n665), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n544), .A2(new_n506), .A3(new_n546), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n776), .A2(new_n547), .A3(new_n777), .ZN(new_n778));
  AOI221_X4 g577(.A(KEYINPUT10), .B1(new_n541), .B2(new_n542), .C1(new_n535), .C2(new_n485), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n535), .A2(new_n537), .A3(new_n485), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n777), .B(new_n505), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n552), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n775), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n505), .B1(new_n779), .B2(new_n780), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n544), .A2(new_n546), .A3(new_n506), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(KEYINPUT54), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n553), .B1(new_n547), .B2(new_n777), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n788), .A3(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n554), .ZN(new_n790));
  INV_X1    g589(.A(new_n610), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n606), .A3(new_n608), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n614), .A2(new_n461), .A3(new_n592), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n564), .B1(new_n793), .B2(new_n591), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n601), .A2(new_n602), .A3(new_n600), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n561), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  NOR4_X1   g596(.A1(new_n662), .A2(new_n784), .A3(new_n790), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n611), .A3(new_n554), .A4(new_n789), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n792), .B(new_n796), .C1(new_n555), .C2(new_n556), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n631), .B1(new_n801), .B2(KEYINPUT117), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n798), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n774), .B1(new_n805), .B2(KEYINPUT118), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807));
  AOI211_X1 g606(.A(new_n807), .B(new_n798), .C1(new_n802), .C2(new_n804), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n773), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(new_n637), .ZN(new_n810));
  INV_X1    g609(.A(new_n433), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(new_n712), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n700), .A2(G113gat), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(KEYINPUT119), .Z(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n809), .A2(new_n436), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n637), .A2(new_n712), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(G113gat), .B1(new_n820), .B2(new_n700), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n816), .A2(new_n821), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n813), .A2(new_n823), .A3(new_n772), .ZN(new_n824));
  OAI21_X1  g623(.A(G120gat), .B1(new_n820), .B2(new_n557), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1341gat));
  AOI21_X1  g625(.A(G127gat), .B1(new_n813), .B2(new_n503), .ZN(new_n827));
  INV_X1    g626(.A(G127gat), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n774), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n827), .B1(new_n819), .B2(new_n829), .ZN(G1342gat));
  INV_X1    g629(.A(G134gat), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n662), .A2(new_n414), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n812), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n820), .B2(new_n662), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(G1343gat));
  NOR2_X1   g636(.A1(new_n278), .A2(new_n334), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n810), .A2(new_n712), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n700), .A2(G141gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n701), .A2(new_n772), .ZN(new_n842));
  XOR2_X1   g641(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n778), .B2(new_n782), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n844), .A2(new_n611), .A3(new_n554), .A4(new_n789), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n845), .A2(new_n846), .A3(new_n800), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n845), .B2(new_n800), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n662), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n798), .ZN(new_n852));
  OAI211_X1 g651(.A(KEYINPUT123), .B(new_n662), .C1(new_n847), .C2(new_n848), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n842), .B1(new_n854), .B2(new_n504), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n334), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n809), .A2(new_n857), .A3(new_n401), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n637), .A2(new_n277), .A3(new_n273), .A4(new_n712), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT120), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G141gat), .B1(new_n861), .B2(new_n700), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n841), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n841), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(KEYINPUT124), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n856), .A2(new_n858), .A3(new_n860), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n611), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n865), .B1(new_n870), .B2(G141gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n864), .B1(new_n871), .B2(new_n863), .ZN(G1344gat));
  INV_X1    g671(.A(G148gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n839), .A2(new_n873), .A3(new_n772), .ZN(new_n874));
  AOI211_X1 g673(.A(KEYINPUT59), .B(new_n873), .C1(new_n869), .C2(new_n772), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n809), .A2(new_n401), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT57), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n503), .B1(new_n849), .B2(new_n852), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n857), .B(new_n401), .C1(new_n842), .C2(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n878), .A2(new_n772), .A3(new_n860), .A4(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n876), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n874), .B1(new_n875), .B2(new_n882), .ZN(G1345gat));
  AOI21_X1  g682(.A(G155gat), .B1(new_n839), .B2(new_n503), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n774), .A2(new_n280), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n869), .B2(new_n885), .ZN(G1346gat));
  NAND4_X1  g685(.A1(new_n810), .A2(new_n281), .A3(new_n832), .A4(new_n838), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n662), .B1(new_n866), .B2(new_n868), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n281), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT125), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n891), .B(new_n887), .C1(new_n888), .C2(new_n281), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1347gat));
  AND2_X1   g692(.A1(new_n809), .A2(new_n654), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n894), .A2(new_n811), .A3(new_n713), .ZN(new_n895));
  INV_X1    g694(.A(G169gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(new_n896), .A3(new_n611), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n637), .A2(new_n397), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n817), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n700), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n897), .A2(new_n902), .ZN(G1348gat));
  AOI21_X1  g702(.A(G176gat), .B1(new_n895), .B2(new_n772), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n772), .A2(G176gat), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n900), .B2(new_n905), .ZN(G1349gat));
  NAND3_X1  g705(.A1(new_n895), .A2(new_n209), .A3(new_n503), .ZN(new_n907));
  OAI21_X1  g706(.A(G183gat), .B1(new_n901), .B2(new_n774), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g709(.A(new_n210), .B1(new_n900), .B2(new_n631), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT61), .Z(new_n912));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n210), .A3(new_n631), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1351gat));
  NOR3_X1   g713(.A1(new_n278), .A2(new_n334), .A3(new_n712), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n894), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT126), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n894), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(G197gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n921), .A3(new_n611), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n899), .A2(new_n278), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n878), .A2(new_n880), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G197gat), .B1(new_n924), .B2(new_n700), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n922), .A2(new_n925), .ZN(G1352gat));
  NOR3_X1   g725(.A1(new_n916), .A2(G204gat), .A3(new_n557), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT62), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n878), .A2(new_n772), .A3(new_n880), .ZN(new_n929));
  INV_X1    g728(.A(new_n923), .ZN(new_n930));
  OAI21_X1  g729(.A(G204gat), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(G1353gat));
  INV_X1    g731(.A(G211gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n920), .A2(new_n933), .A3(new_n503), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n924), .A2(new_n504), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  AOI21_X1  g738(.A(new_n662), .B1(new_n917), .B2(new_n919), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n631), .A2(G218gat), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n940), .A2(G218gat), .B1(new_n924), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT127), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944));
  OAI221_X1 g743(.A(new_n944), .B1(new_n924), .B2(new_n941), .C1(new_n940), .C2(G218gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1355gat));
endmodule


