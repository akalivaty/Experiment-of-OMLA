//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n212), .B1(new_n214), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT64), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n228), .B(new_n232), .Z(G358));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XNOR2_X1  g0034(.A(G107), .B(G116), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G50), .B(G68), .Z(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  NOR2_X1   g0040(.A1(G20), .A2(G33), .ZN(new_n241));
  AOI22_X1  g0041(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G33), .ZN(new_n243));
  OAI21_X1  g0043(.A(KEYINPUT65), .B1(new_n243), .B2(G20), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT65), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(new_n207), .A3(G33), .ZN(new_n246));
  AND2_X1   g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n242), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n202), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n251), .A3(new_n250), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n206), .A2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n253), .B(new_n256), .C1(new_n257), .C2(new_n259), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n260), .A2(KEYINPUT9), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(KEYINPUT9), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G222), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G77), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(G223), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n267), .B1(new_n268), .B2(new_n265), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G226), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(new_n213), .B2(new_n272), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n279), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n275), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n261), .A2(new_n262), .B1(G200), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT70), .ZN(new_n289));
  INV_X1    g0089(.A(new_n286), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(G190), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n286), .A2(KEYINPUT70), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT10), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n291), .A2(new_n293), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(new_n287), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n260), .B1(new_n290), .B2(G169), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT66), .B(G179), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n286), .A2(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT16), .ZN(new_n306));
  INV_X1    g0106(.A(G68), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n263), .A2(new_n207), .A3(new_n264), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT7), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n264), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G58), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(new_n307), .ZN(new_n314));
  OAI21_X1  g0114(.A(G20), .B1(new_n314), .B2(new_n201), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n241), .A2(G159), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n306), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT7), .B1(new_n321), .B2(new_n207), .ZN(new_n322));
  NOR4_X1   g0122(.A1(new_n319), .A2(new_n320), .A3(new_n309), .A4(G20), .ZN(new_n323));
  OAI21_X1  g0123(.A(G68), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n317), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n318), .A2(new_n326), .A3(new_n252), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n270), .A2(new_n266), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n278), .A2(G1698), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n328), .B(new_n329), .C1(new_n319), .C2(new_n320), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G87), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n274), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n284), .A2(new_n273), .A3(G274), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n273), .A2(G232), .A3(new_n276), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(new_n336), .A3(new_n292), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n273), .B1(new_n330), .B2(new_n331), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(new_n335), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT75), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n248), .A2(new_n255), .ZN(new_n344));
  INV_X1    g0144(.A(new_n248), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n258), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n343), .B(new_n344), .C1(new_n346), .C2(new_n257), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n257), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(new_n345), .A3(new_n258), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n343), .B1(new_n350), .B2(new_n344), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n327), .A2(new_n342), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT17), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n355));
  NAND4_X1  g0155(.A1(new_n327), .A2(new_n352), .A3(new_n342), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT18), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n344), .B1(new_n346), .B2(new_n257), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT75), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n347), .ZN(new_n362));
  INV_X1    g0162(.A(new_n252), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n324), .A2(new_n325), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(new_n306), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n362), .B1(new_n365), .B2(new_n326), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n333), .B2(new_n336), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n339), .A2(new_n340), .A3(new_n301), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g0170(.A(KEYINPUT77), .B(new_n359), .C1(new_n366), .C2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT77), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n370), .B1(new_n327), .B2(new_n352), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n373), .B2(KEYINPUT18), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT76), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n327), .A2(new_n352), .ZN(new_n377));
  INV_X1    g0177(.A(new_n370), .ZN(new_n378));
  AND4_X1   g0178(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT18), .A4(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n373), .B2(KEYINPUT18), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n358), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G238), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n334), .B1(new_n384), .B2(new_n277), .ZN(new_n385));
  OAI211_X1 g0185(.A(G232), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT71), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT71), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n265), .A2(new_n388), .A3(G232), .A4(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G97), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n265), .A2(G226), .A3(new_n266), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n387), .A2(new_n389), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n385), .B1(new_n392), .B2(new_n274), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI211_X1 g0195(.A(KEYINPUT13), .B(new_n385), .C1(new_n392), .C2(new_n274), .ZN(new_n396));
  OAI21_X1  g0196(.A(G169), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT14), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(G169), .C1(new_n395), .C2(new_n396), .ZN(new_n400));
  INV_X1    g0200(.A(new_n396), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT72), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n393), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT13), .B1(new_n393), .B2(new_n402), .ZN(new_n404));
  OAI211_X1 g0204(.A(G179), .B(new_n401), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n398), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n247), .A2(new_n268), .ZN(new_n407));
  INV_X1    g0207(.A(new_n241), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n408), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n252), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT11), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT68), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n363), .A2(new_n412), .A3(new_n254), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n257), .A2(KEYINPUT68), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(G68), .A4(new_n258), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT73), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT74), .B1(new_n254), .B2(G68), .ZN(new_n417));
  XOR2_X1   g0217(.A(new_n417), .B(KEYINPUT12), .Z(new_n418));
  AND3_X1   g0218(.A1(new_n411), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n406), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(G190), .B(new_n401), .C1(new_n403), .C2(new_n404), .ZN(new_n422));
  OAI21_X1  g0222(.A(G200), .B1(new_n395), .B2(new_n396), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G244), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n334), .B1(new_n426), .B2(new_n277), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT67), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n334), .B(KEYINPUT67), .C1(new_n426), .C2(new_n277), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n265), .A2(G232), .A3(new_n266), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n321), .A2(G107), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(new_n269), .C2(new_n384), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n274), .ZN(new_n435));
  AOI21_X1  g0235(.A(G169), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT69), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n429), .A3(new_n430), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n436), .A2(new_n437), .B1(new_n302), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n431), .A2(KEYINPUT69), .A3(new_n301), .A4(new_n435), .ZN(new_n440));
  XOR2_X1   g0240(.A(KEYINPUT15), .B(G87), .Z(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(new_n247), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n248), .A2(new_n408), .B1(new_n207), .B2(new_n268), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n252), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n413), .A2(new_n414), .A3(G77), .A4(new_n258), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n446), .C1(G77), .C2(new_n254), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n431), .A2(G190), .A3(new_n435), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n447), .B1(G200), .B2(new_n438), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n439), .A2(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g0252(.A1(new_n305), .A2(new_n383), .A3(new_n425), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  INV_X1    g0255(.A(G97), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n455), .B(new_n207), .C1(G33), .C2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G116), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G20), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n252), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT20), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n457), .A2(KEYINPUT20), .A3(new_n252), .A4(new_n459), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT83), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(new_n254), .B2(G116), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n255), .A2(KEYINPUT83), .A3(new_n458), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n462), .A2(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n458), .B1(new_n206), .B2(G33), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n413), .A2(new_n414), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(G264), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n472));
  OAI211_X1 g0272(.A(G257), .B(new_n266), .C1(new_n319), .C2(new_n320), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n263), .A2(G303), .A3(new_n264), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n475), .A2(new_n274), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT5), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT80), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(G41), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n282), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n206), .A2(G45), .ZN(new_n482));
  OAI211_X1 g0282(.A(G270), .B(new_n273), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n482), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n281), .A2(new_n484), .A3(new_n480), .A4(new_n479), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT82), .B1(new_n476), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n483), .A2(new_n485), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT82), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n475), .A2(new_n274), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(new_n491), .A3(G200), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n487), .A2(new_n491), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n471), .B(new_n492), .C1(new_n493), .C2(new_n292), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n367), .B1(new_n467), .B2(new_n469), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n495), .A2(new_n487), .A3(new_n491), .A4(KEYINPUT21), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n488), .A2(G179), .A3(new_n490), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n470), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n495), .A2(new_n487), .A3(new_n491), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT84), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT21), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(new_n501), .B2(new_n503), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n494), .B(new_n500), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n207), .B2(G107), .ZN(new_n508));
  INV_X1    g0308(.A(G107), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(KEYINPUT23), .A3(G20), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G116), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(G20), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n207), .B(G87), .C1(new_n319), .C2(new_n320), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT85), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n265), .A2(KEYINPUT85), .A3(new_n207), .A4(G87), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT22), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT86), .B1(new_n514), .B2(KEYINPUT22), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n513), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  XOR2_X1   g0321(.A(KEYINPUT87), .B(KEYINPUT24), .Z(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT86), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n516), .A2(new_n517), .A3(new_n524), .A4(KEYINPUT22), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n523), .B1(new_n521), .B2(new_n525), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n252), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n349), .B1(G1), .B2(new_n243), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT25), .B1(new_n255), .B2(new_n509), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n255), .A2(KEYINPUT25), .A3(new_n509), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n531), .A2(G107), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n265), .A2(G257), .A3(G1698), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G294), .ZN(new_n537));
  OAI211_X1 g0337(.A(G250), .B(new_n266), .C1(new_n319), .C2(new_n320), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n274), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n479), .A2(new_n480), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n274), .B1(new_n541), .B2(new_n484), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G264), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n543), .A3(new_n485), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n338), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(G190), .B2(new_n544), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n529), .A2(new_n535), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  AND2_X1   g0348(.A1(G97), .A2(G107), .ZN(new_n549));
  NOR2_X1   g0349(.A1(G97), .A2(G107), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n509), .A2(KEYINPUT6), .A3(G97), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n553), .A2(new_n207), .B1(new_n268), .B2(new_n408), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n509), .B1(new_n310), .B2(new_n311), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n252), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n255), .A2(new_n456), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n531), .A2(G97), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(G250), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n560));
  OAI211_X1 g0360(.A(G244), .B(new_n266), .C1(new_n319), .C2(new_n320), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT4), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n455), .B(new_n560), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  XOR2_X1   g0363(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n564));
  AND2_X1   g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n274), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(G257), .B(new_n273), .C1(new_n481), .C2(new_n482), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n567), .A2(new_n485), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n367), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n566), .A2(new_n568), .A3(new_n301), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n559), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(G200), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n557), .B1(new_n530), .B2(new_n456), .ZN(new_n574));
  OAI21_X1  g0374(.A(G107), .B1(new_n322), .B2(new_n323), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n551), .A2(new_n552), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(G20), .B1(G77), .B2(new_n241), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n574), .B1(new_n252), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n566), .A2(new_n568), .A3(G190), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n573), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n572), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n265), .A2(new_n207), .A3(G68), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n456), .B1(new_n244), .B2(new_n246), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n207), .B1(new_n390), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n550), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT81), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n586), .B2(new_n588), .ZN(new_n591));
  OAI221_X1 g0391(.A(new_n583), .B1(new_n584), .B2(KEYINPUT19), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n252), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n442), .A2(new_n255), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n531), .A2(G87), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(G244), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n597));
  OAI211_X1 g0397(.A(G238), .B(new_n266), .C1(new_n319), .C2(new_n320), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(new_n512), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n274), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n281), .A2(new_n484), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n273), .A2(G250), .A3(new_n482), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n603), .A3(new_n292), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n602), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n599), .B2(new_n274), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n604), .B1(new_n606), .B2(G200), .ZN(new_n607));
  AOI21_X1  g0407(.A(G169), .B1(new_n600), .B2(new_n603), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n301), .B2(new_n606), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n531), .A2(new_n441), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n593), .A2(new_n594), .A3(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n596), .A2(new_n607), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n547), .A2(new_n582), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n544), .A2(G169), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT88), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n274), .A2(new_n539), .B1(new_n542), .B2(G264), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(G179), .A3(new_n485), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n544), .A2(KEYINPUT88), .A3(G169), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n521), .A2(new_n525), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n522), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n363), .B1(new_n622), .B2(new_n526), .ZN(new_n623));
  INV_X1    g0423(.A(new_n535), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NOR4_X1   g0426(.A1(new_n454), .A2(new_n506), .A3(new_n613), .A4(new_n626), .ZN(G372));
  NOR2_X1   g0427(.A1(new_n300), .A2(new_n303), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n377), .A2(new_n378), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n359), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n377), .A2(KEYINPUT18), .A3(new_n378), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n437), .B1(new_n438), .B2(new_n367), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n438), .A2(new_n302), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n440), .B(new_n447), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n420), .A2(new_n406), .B1(new_n424), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(KEYINPUT89), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n357), .B1(new_n637), .B2(KEYINPUT89), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n632), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n628), .B1(new_n640), .B2(new_n299), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n625), .B(new_n500), .C1(new_n505), .C2(new_n504), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n609), .A2(new_n611), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n607), .A2(new_n593), .A3(new_n594), .A4(new_n595), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n572), .A2(new_n643), .A3(new_n581), .A4(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n623), .A2(new_n624), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(new_n546), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n643), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n643), .A2(new_n644), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(new_n572), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n559), .A2(new_n570), .A3(new_n571), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n612), .A2(KEYINPUT26), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n649), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n648), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n453), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n641), .A2(new_n657), .ZN(G369));
  OAI21_X1  g0458(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n659));
  INV_X1    g0459(.A(G13), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n660), .A2(G1), .A3(G20), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT90), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G213), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n471), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n659), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n506), .B2(new_n669), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n547), .B1(new_n646), .B2(new_n668), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n625), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n626), .A2(new_n668), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n674), .A2(new_n659), .A3(new_n625), .A4(new_n668), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n675), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT91), .ZN(G399));
  INV_X1    g0483(.A(new_n210), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G1), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n550), .A2(new_n587), .A3(new_n458), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT92), .Z(new_n689));
  OAI22_X1  g0489(.A1(new_n687), .A2(new_n689), .B1(new_n215), .B2(new_n686), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  INV_X1    g0491(.A(new_n668), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n648), .B2(new_n655), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(KEYINPUT29), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT29), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n649), .B1(new_n642), .B2(new_n647), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT26), .B1(new_n612), .B2(new_n653), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n654), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n612), .A2(KEYINPUT94), .A3(KEYINPUT26), .A4(new_n653), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n696), .B1(new_n703), .B2(new_n668), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n695), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT31), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n617), .A2(new_n606), .A3(new_n566), .A4(new_n568), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT30), .B1(new_n707), .B2(new_n497), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n606), .A2(new_n543), .A3(new_n540), .ZN(new_n709));
  INV_X1    g0509(.A(new_n569), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n709), .A2(new_n498), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n606), .A2(new_n302), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n713), .A2(new_n544), .A3(new_n569), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n708), .A2(new_n712), .B1(new_n714), .B2(new_n493), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT93), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n692), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n708), .A2(new_n712), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n714), .A2(new_n493), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n718), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n706), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n506), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n647), .A3(new_n625), .A4(new_n668), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(G330), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n705), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n691), .B1(new_n730), .B2(G1), .ZN(G364));
  NOR2_X1   g0531(.A1(new_n660), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n206), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n685), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n213), .B1(new_n207), .B2(G169), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT96), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(KEYINPUT96), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n207), .B1(new_n742), .B2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G97), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n207), .A2(new_n292), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n338), .A2(G179), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n745), .B(new_n265), .C1(new_n587), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n207), .A2(G190), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n742), .ZN(new_n751));
  INV_X1    g0551(.A(G159), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT32), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n750), .A2(new_n747), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT99), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G107), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n301), .A2(new_n207), .A3(new_n338), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n292), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n754), .B(new_n757), .C1(new_n307), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n301), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n750), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n749), .B(new_n760), .C1(G77), .C2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT98), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n758), .A2(new_n765), .A3(G190), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(new_n758), .B2(G190), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n761), .A2(KEYINPUT97), .A3(new_n746), .ZN(new_n769));
  AOI21_X1  g0569(.A(KEYINPUT97), .B1(new_n761), .B2(new_n746), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n764), .B1(new_n202), .B2(new_n768), .C1(new_n313), .C2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n756), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n773), .A2(new_n774), .B1(new_n775), .B2(new_n762), .ZN(new_n776));
  INV_X1    g0576(.A(new_n759), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G329), .ZN(new_n780));
  INV_X1    g0580(.A(G294), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n751), .B1(new_n743), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n321), .B1(new_n748), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT101), .ZN(new_n785));
  NOR4_X1   g0585(.A1(new_n776), .A2(new_n779), .A3(new_n782), .A4(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT100), .B(G326), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n786), .B1(new_n787), .B2(new_n771), .C1(new_n768), .C2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n741), .B1(new_n772), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n740), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n684), .A2(new_n265), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(G45), .B2(new_n215), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n239), .A2(new_n283), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n684), .A2(new_n321), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G355), .B1(new_n458), .B2(new_n684), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n798), .B1(KEYINPUT95), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(KEYINPUT95), .B2(new_n801), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n736), .B(new_n790), .C1(new_n794), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n793), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n671), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n672), .A2(new_n735), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(G330), .B2(new_n671), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  NAND2_X1  g0610(.A1(new_n741), .A2(new_n792), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n735), .B1(new_n811), .B2(G77), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n777), .A2(G150), .B1(new_n763), .B2(G159), .ZN(new_n813));
  INV_X1    g0613(.A(G143), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n813), .B1(new_n771), .B2(new_n814), .C1(new_n768), .C2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT34), .Z(new_n817));
  AND3_X1   g0617(.A1(new_n750), .A2(G132), .A3(new_n742), .ZN(new_n818));
  INV_X1    g0618(.A(new_n748), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n321), .B(new_n818), .C1(G50), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n756), .A2(G68), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(new_n313), .C2(new_n743), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n756), .A2(G87), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n775), .B2(new_n751), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT102), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n265), .B1(new_n819), .B2(G107), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n826), .B(new_n745), .C1(new_n458), .C2(new_n762), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G283), .B2(new_n777), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n828), .B1(new_n781), .B2(new_n771), .C1(new_n783), .C2(new_n768), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n817), .A2(new_n822), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n830), .A2(new_n740), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT103), .B1(new_n635), .B2(new_n668), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT103), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n439), .A2(new_n448), .A3(new_n833), .A4(new_n692), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n692), .A2(new_n447), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n832), .A2(new_n834), .B1(new_n451), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n812), .B(new_n831), .C1(new_n791), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n728), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n694), .A2(new_n836), .ZN(new_n839));
  INV_X1    g0639(.A(new_n836), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n693), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n838), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT104), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n736), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n842), .A2(KEYINPUT104), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n837), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G384));
  NOR2_X1   g0649(.A1(new_n732), .A2(new_n206), .ZN(new_n850));
  INV_X1    g0650(.A(G330), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n722), .A2(KEYINPUT93), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n715), .A2(new_n716), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n852), .A2(KEYINPUT31), .A3(new_n853), .A4(new_n692), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n726), .A2(new_n721), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n420), .A2(new_n692), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n421), .A2(new_n424), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n422), .A2(new_n419), .A3(new_n423), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n420), .B(new_n692), .C1(new_n858), .C2(new_n406), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n836), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n855), .A2(new_n860), .A3(KEYINPUT40), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n357), .A2(KEYINPUT108), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT108), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n354), .A2(new_n863), .A3(new_n356), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n632), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n377), .A2(new_n667), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n629), .A2(new_n866), .A3(new_n353), .ZN(new_n869));
  XOR2_X1   g0669(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n869), .B(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n327), .A2(new_n344), .A3(new_n350), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n667), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n631), .A2(KEYINPUT76), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n373), .A2(new_n376), .A3(KEYINPUT18), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(new_n371), .A3(new_n374), .A4(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n875), .B1(new_n878), .B2(new_n357), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n629), .A2(new_n866), .A3(new_n353), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n874), .A2(new_n378), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n875), .A2(new_n882), .A3(new_n353), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n881), .A2(new_n870), .B1(new_n883), .B2(KEYINPUT37), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n879), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT110), .B1(new_n873), .B2(new_n885), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n357), .A2(KEYINPUT108), .B1(new_n630), .B2(new_n631), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n866), .B1(new_n887), .B2(new_n864), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n869), .B(new_n870), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n880), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n883), .A2(KEYINPUT37), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n871), .B2(new_n869), .ZN(new_n892));
  OAI211_X1 g0692(.A(KEYINPUT38), .B(new_n892), .C1(new_n382), .C2(new_n875), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT110), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n890), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n861), .A2(new_n886), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n880), .B1(new_n879), .B2(new_n884), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n855), .A2(new_n860), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n902), .B(KEYINPUT111), .Z(new_n903));
  INV_X1    g0703(.A(new_n855), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n454), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n851), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n453), .B1(new_n695), .B2(new_n704), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n641), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT109), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n632), .A2(new_n667), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n857), .A2(new_n859), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n635), .A2(new_n692), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n913), .B1(new_n841), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n893), .A2(new_n898), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n873), .B2(new_n885), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n406), .A2(new_n420), .A3(new_n668), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT107), .Z(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n893), .A2(new_n898), .A3(KEYINPUT39), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n918), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n910), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n850), .B1(new_n907), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n927), .B2(new_n907), .ZN(new_n929));
  OAI21_X1  g0729(.A(G77), .B1(new_n313), .B2(new_n307), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n930), .A2(new_n215), .B1(G50), .B2(new_n307), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(G1), .A3(new_n660), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT105), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n458), .B(new_n214), .C1(new_n576), .C2(KEYINPUT35), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(KEYINPUT35), .B2(new_n576), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT36), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n936), .B2(new_n935), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n929), .A2(new_n938), .ZN(G367));
  OAI21_X1  g0739(.A(new_n582), .B1(new_n579), .B2(new_n668), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n653), .A2(new_n692), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n680), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n572), .B1(new_n940), .B2(new_n625), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n943), .A2(KEYINPUT42), .B1(new_n668), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(KEYINPUT42), .B2(new_n943), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n596), .A2(new_n668), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n649), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n651), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT112), .Z(new_n951));
  AOI22_X1  g0751(.A1(new_n951), .A2(KEYINPUT113), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n678), .A2(new_n942), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n946), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n953), .B1(new_n946), .B2(new_n952), .ZN(new_n956));
  OR4_X1    g0756(.A1(KEYINPUT113), .A2(new_n955), .A3(new_n951), .A4(new_n956), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n955), .A2(new_n956), .B1(KEYINPUT113), .B2(new_n951), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n685), .B(KEYINPUT41), .Z(new_n959));
  NAND2_X1  g0759(.A1(new_n681), .A2(new_n942), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT44), .Z(new_n961));
  NOR2_X1   g0761(.A1(new_n681), .A2(new_n942), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n679), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n659), .A2(new_n668), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n676), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n680), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(new_n672), .Z(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(new_n729), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n961), .A2(new_n678), .A3(new_n963), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n965), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n959), .B1(new_n972), .B2(new_n730), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n957), .B(new_n958), .C1(new_n973), .C2(new_n734), .ZN(new_n974));
  INV_X1    g0774(.A(new_n795), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n232), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n794), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n684), .B2(new_n441), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n736), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n768), .ZN(new_n980));
  INV_X1    g0780(.A(new_n771), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n980), .A2(G143), .B1(new_n981), .B2(G150), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n743), .A2(new_n307), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n265), .B1(new_n755), .B2(new_n268), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(new_n777), .C2(G159), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n748), .A2(new_n313), .B1(new_n751), .B2(new_n815), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT115), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n762), .A2(new_n202), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n987), .B2(new_n986), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n982), .A2(new_n985), .A3(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT114), .B(G311), .Z(new_n991));
  NAND2_X1  g0791(.A1(new_n980), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(G317), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n321), .B1(new_n751), .B2(new_n993), .C1(new_n456), .C2(new_n755), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n762), .A2(new_n774), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G294), .C2(new_n777), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n748), .A2(new_n458), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT46), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G107), .B2(new_n744), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n981), .A2(G303), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n992), .A2(new_n996), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n990), .A2(KEYINPUT47), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n740), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT47), .B1(new_n990), .B2(new_n1001), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n979), .B1(new_n949), .B2(new_n805), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n974), .A2(new_n1005), .ZN(G387));
  AOI21_X1  g0806(.A(new_n975), .B1(new_n228), .B2(G45), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n689), .B2(new_n799), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT50), .B1(new_n248), .B2(G50), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1009), .B(new_n283), .C1(new_n307), .C2(new_n268), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n248), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1010), .A2(new_n689), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n509), .B2(new_n684), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n735), .B1(new_n1014), .B2(new_n977), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT116), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n773), .A2(new_n456), .B1(new_n307), .B2(new_n762), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n442), .A2(new_n743), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(KEYINPUT117), .B(G150), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n265), .B1(new_n751), .B2(new_n1019), .C1(new_n268), .C2(new_n748), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n759), .A2(new_n248), .ZN(new_n1021));
  NOR4_X1   g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n202), .B2(new_n771), .C1(new_n752), .C2(new_n768), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n755), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n265), .B1(new_n1024), .B2(G116), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n748), .A2(new_n781), .B1(new_n743), .B2(new_n774), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n777), .A2(new_n991), .B1(new_n763), .B2(G303), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n771), .B2(new_n993), .C1(new_n768), .C2(new_n787), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT48), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT49), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1025), .B1(new_n751), .B2(new_n788), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1023), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1016), .B1(new_n740), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n676), .A2(new_n793), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n970), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n685), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n969), .A2(new_n729), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1038), .B1(new_n733), .B2(new_n969), .C1(new_n1040), .C2(new_n1041), .ZN(G393));
  INV_X1    g0842(.A(new_n971), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n678), .B1(new_n961), .B2(new_n963), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1043), .A2(new_n733), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n942), .A2(new_n793), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n794), .B1(new_n456), .B2(new_n210), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n975), .A2(new_n236), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n735), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n321), .B1(new_n751), .B2(new_n787), .C1(new_n774), .C2(new_n748), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n757), .B1(new_n781), .B2(new_n762), .C1(new_n783), .C2(new_n759), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(G116), .C2(new_n744), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n768), .A2(new_n993), .B1(new_n771), .B2(new_n775), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT52), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(G150), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n768), .A2(new_n1056), .B1(new_n771), .B2(new_n752), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT51), .Z(new_n1058));
  OAI221_X1 g0858(.A(new_n823), .B1(new_n202), .B2(new_n759), .C1(new_n248), .C2(new_n762), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n743), .A2(new_n268), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n265), .B1(new_n751), .B2(new_n814), .C1(new_n307), .C2(new_n748), .ZN(new_n1061));
  OR3_X1    g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1055), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1049), .B1(new_n1063), .B2(new_n740), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1045), .B1(new_n1046), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1039), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1066), .A2(new_n685), .A3(new_n972), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1067), .ZN(G390));
  XNOR2_X1  g0868(.A(KEYINPUT54), .B(G143), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n759), .A2(new_n815), .B1(new_n762), .B2(new_n1069), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n748), .A2(new_n1019), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1071), .A2(KEYINPUT53), .B1(G159), .B2(new_n744), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(KEYINPUT53), .B2(new_n1071), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1070), .B(new_n1073), .C1(new_n980), .C2(G128), .ZN(new_n1074));
  INV_X1    g0874(.A(G125), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n265), .B1(new_n751), .B2(new_n1075), .C1(new_n202), .C2(new_n755), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT120), .Z(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G132), .B2(new_n981), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n821), .B1(new_n456), .B2(new_n762), .C1(new_n509), .C2(new_n759), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n321), .B1(new_n751), .B2(new_n781), .C1(new_n587), .C2(new_n748), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1079), .A2(new_n1060), .A3(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n980), .A2(G283), .B1(new_n981), .B2(G116), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1074), .A2(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n735), .B1(new_n345), .B2(new_n811), .C1(new_n1083), .C2(new_n741), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n920), .A2(new_n924), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n791), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n886), .A2(new_n895), .A3(new_n922), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n692), .B(new_n836), .C1(new_n697), .C2(new_n702), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n912), .B1(new_n1088), .B2(new_n914), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n914), .B1(new_n693), .B2(new_n840), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n922), .B1(new_n1090), .B2(new_n913), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1087), .A2(new_n1089), .B1(new_n1091), .B2(new_n1085), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT118), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n838), .A2(new_n840), .A3(new_n912), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1089), .A2(new_n922), .A3(new_n886), .A4(new_n895), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1091), .A2(new_n1085), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT118), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n855), .A2(G330), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n860), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1092), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1095), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1086), .B1(new_n1104), .B2(new_n734), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n913), .B1(new_n728), .B2(new_n836), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1090), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT119), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1100), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n855), .A2(KEYINPUT119), .A3(G330), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n840), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1113), .A2(new_n913), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1088), .A2(new_n914), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1094), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1109), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1101), .A2(new_n453), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n908), .A2(new_n641), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n685), .B1(new_n1104), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1093), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(new_n860), .A3(new_n1101), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1123), .B1(new_n1127), .B2(new_n1095), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1105), .B1(new_n1122), .B2(new_n1128), .ZN(G378));
  NAND3_X1  g0929(.A1(new_n896), .A2(new_n901), .A3(G330), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n305), .A2(new_n260), .A3(new_n667), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n667), .A2(new_n260), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n299), .A2(new_n304), .A3(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1130), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n918), .A2(new_n925), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n917), .A2(new_n855), .A3(new_n860), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n851), .B1(new_n1140), .B2(new_n897), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n896), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1138), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT122), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1138), .A2(KEYINPUT122), .A3(new_n1139), .A4(new_n1143), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1139), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1148), .A2(KEYINPUT123), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT123), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1150), .B(new_n1139), .C1(new_n1138), .C2(new_n1143), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1146), .B(new_n1147), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1152));
  AND4_X1   g0952(.A1(new_n1093), .A2(new_n1096), .A3(new_n1097), .A4(new_n1094), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1120), .B1(new_n1154), .B2(new_n1123), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT57), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1119), .B1(new_n1104), .B2(new_n1121), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1141), .A2(new_n1142), .A3(new_n896), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1142), .B1(new_n1141), .B2(new_n896), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n926), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1144), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT57), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n685), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1156), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1142), .A2(new_n791), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n735), .B1(new_n811), .B2(G50), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(G33), .A2(G41), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G50), .B(new_n1167), .C1(new_n321), .C2(new_n282), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n759), .A2(new_n456), .B1(new_n762), .B2(new_n442), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n282), .B(new_n321), .C1(new_n748), .C2(new_n268), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n755), .A2(new_n313), .B1(new_n751), .B2(new_n774), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1169), .A2(new_n983), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n509), .B2(new_n771), .C1(new_n458), .C2(new_n768), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1168), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n748), .A2(new_n1069), .B1(new_n743), .B2(new_n1056), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n762), .A2(new_n815), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(G132), .C2(new_n777), .ZN(new_n1178));
  INV_X1    g0978(.A(G128), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1178), .B1(new_n1075), .B2(new_n768), .C1(new_n1179), .C2(new_n771), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  INV_X1    g0981(.A(G124), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1167), .B1(new_n751), .B2(new_n1182), .C1(new_n752), .C2(new_n755), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT121), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1175), .B1(new_n1174), .B2(new_n1173), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1166), .B1(new_n1187), .B2(new_n740), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1165), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1152), .B2(new_n734), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1164), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT124), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT124), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1164), .A2(new_n1194), .A3(new_n1191), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(G375));
  INV_X1    g0997(.A(new_n959), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1119), .B(new_n1109), .C1(new_n1114), .C2(new_n1116), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1123), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n733), .B(KEYINPUT125), .Z(new_n1201));
  NAND2_X1  g1001(.A1(new_n913), .A2(new_n791), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n735), .B1(new_n811), .B2(G68), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n773), .A2(new_n268), .B1(new_n458), .B2(new_n759), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n321), .B1(new_n751), .B2(new_n783), .C1(new_n456), .C2(new_n748), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n762), .A2(new_n509), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1204), .A2(new_n1018), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n774), .B2(new_n771), .C1(new_n781), .C2(new_n768), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n980), .A2(G132), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n981), .A2(G137), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n265), .B1(new_n755), .B2(new_n313), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n748), .A2(new_n752), .B1(new_n751), .B2(new_n1179), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(G50), .C2(new_n744), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1069), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n777), .A2(new_n1214), .B1(new_n763), .B2(G150), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1209), .A2(new_n1210), .A3(new_n1213), .A4(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1208), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1203), .B1(new_n1217), .B2(new_n740), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1117), .A2(new_n1201), .B1(new_n1202), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1200), .A2(new_n1219), .ZN(G381));
  INV_X1    g1020(.A(G378), .ZN(new_n1221));
  OR3_X1    g1021(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(G387), .A2(new_n1222), .A3(G381), .A4(G390), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1196), .A2(new_n1221), .A3(new_n1223), .ZN(G407));
  AOI21_X1  g1024(.A(G378), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(G407), .B(G213), .C1(new_n1226), .C2(G343), .ZN(G409));
  INV_X1    g1027(.A(KEYINPUT126), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1190), .B1(new_n1161), .B2(new_n1201), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1160), .A2(new_n1150), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1148), .A2(KEYINPUT123), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n959), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1230), .B1(new_n1235), .B2(new_n1155), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1228), .B1(new_n1236), .B2(G378), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G378), .B(new_n1191), .C1(new_n1156), .C2(new_n1163), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1152), .A2(new_n1155), .A3(new_n1198), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1229), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(KEYINPUT126), .A3(new_n1221), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1237), .A2(new_n1238), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(G343), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(G213), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT60), .ZN(new_n1245));
  OAI211_X1 g1045(.A(KEYINPUT127), .B(new_n1199), .C1(new_n1121), .C2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT127), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1245), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1199), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n686), .B1(new_n1249), .B2(KEYINPUT60), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1246), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1252), .A2(G384), .A3(new_n1219), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G384), .B1(new_n1252), .B2(new_n1219), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1242), .A2(new_n1244), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT62), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1243), .A2(G213), .A3(G2897), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1252), .A2(new_n1219), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n848), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1252), .A2(G384), .A3(new_n1219), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1259), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1261), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1258), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1242), .A2(new_n1269), .A3(new_n1244), .A4(new_n1255), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1257), .A2(new_n1267), .A3(new_n1268), .A4(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G393), .B(new_n809), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n974), .A2(G390), .A3(new_n1005), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G390), .B1(new_n974), .B2(new_n1005), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(G390), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G387), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n974), .A2(G390), .A3(new_n1005), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1272), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1271), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1256), .B2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT61), .B1(new_n1258), .B2(new_n1266), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1284), .B(new_n1285), .C1(new_n1283), .C2(new_n1256), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1282), .A2(new_n1286), .ZN(G405));
  AOI21_X1  g1087(.A(new_n1221), .B1(new_n1164), .B2(new_n1191), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1225), .A2(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1276), .A2(new_n1255), .A3(new_n1280), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1255), .B1(new_n1276), .B2(new_n1280), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1289), .B(new_n1292), .ZN(G402));
endmodule


