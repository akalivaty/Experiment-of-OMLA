//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927;
  OAI21_X1  g000(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g002(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n203), .A2(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT64), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT25), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n208), .B(new_n209), .C1(new_n210), .C2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(KEYINPUT65), .A3(new_n214), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n213), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n215), .B1(KEYINPUT65), .B2(new_n214), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT25), .B1(new_n221), .B2(new_n207), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT27), .B(G183gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(new_n212), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT28), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NOR3_X1   g025(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT26), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(new_n205), .B2(new_n206), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n215), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n217), .A2(new_n222), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G134gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G127gat), .ZN(new_n233));
  INV_X1    g032(.A(G127gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G134gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G120gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n238));
  INV_X1    g037(.A(G120gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G113gat), .ZN(new_n240));
  INV_X1    g039(.A(G113gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G120gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G127gat), .B(G134gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n238), .A2(new_n246), .A3(KEYINPUT67), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n230), .A2(new_n222), .ZN(new_n253));
  INV_X1    g052(.A(new_n251), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n217), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G227gat), .ZN(new_n257));
  INV_X1    g056(.A(G233gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT33), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n259), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n252), .B2(new_n255), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT68), .B1(new_n265), .B2(KEYINPUT33), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n260), .A2(KEYINPUT32), .ZN(new_n267));
  XNOR2_X1  g066(.A(G15gat), .B(G43gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(G71gat), .ZN(new_n269));
  INV_X1    g068(.A(G99gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n263), .A2(new_n266), .A3(new_n267), .A4(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(KEYINPUT33), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n260), .A2(KEYINPUT32), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n252), .A2(new_n255), .A3(new_n264), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT34), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT69), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n277), .A2(KEYINPUT69), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(new_n279), .B2(new_n276), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n275), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT3), .ZN(new_n284));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285));
  INV_X1    g084(.A(G211gat), .ZN(new_n286));
  INV_X1    g085(.A(G218gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n285), .B1(KEYINPUT22), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n284), .B1(new_n291), .B2(KEYINPUT29), .ZN(new_n292));
  XNOR2_X1  g091(.A(G141gat), .B(G148gat), .ZN(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(G162gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(G155gat), .ZN(new_n297));
  OAI22_X1  g096(.A1(new_n293), .A2(KEYINPUT2), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G148gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G141gat), .ZN(new_n300));
  INV_X1    g099(.A(G141gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G148gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G155gat), .B(G162gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT2), .B1(new_n305), .B2(new_n296), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n298), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n298), .A2(new_n307), .A3(new_n284), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n298), .A2(new_n307), .A3(KEYINPUT73), .A4(new_n284), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT29), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n291), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G228gat), .A2(G233gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(G22gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT79), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n319), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT31), .B(G50gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G78gat), .B(G106gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n283), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330));
  INV_X1    g129(.A(G64gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G92gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n231), .A2(KEYINPUT70), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT70), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n253), .A2(new_n337), .A3(new_n217), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(KEYINPUT29), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n231), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n315), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n336), .A2(new_n338), .A3(new_n342), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n253), .A2(new_n217), .A3(new_n340), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n315), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n335), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n339), .A2(new_n340), .B1(new_n231), .B2(new_n342), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n347), .B(new_n334), .C1(new_n350), .C2(new_n315), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT30), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n347), .B1(new_n350), .B2(new_n315), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n335), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n243), .A2(new_n245), .B1(new_n233), .B2(new_n235), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n238), .A2(new_n246), .A3(KEYINPUT72), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n312), .A2(new_n313), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n308), .A2(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(new_n251), .B2(new_n308), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n308), .A2(new_n247), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n364), .B(new_n366), .C1(new_n365), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OR3_X1    g169(.A1(new_n368), .A2(KEYINPUT5), .A3(new_n370), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n362), .A2(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n372));
  INV_X1    g171(.A(new_n308), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n249), .A2(new_n373), .A3(KEYINPUT4), .A4(new_n250), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n374), .A2(new_n369), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n238), .A2(new_n246), .A3(KEYINPUT72), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT72), .B1(new_n238), .B2(new_n246), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n308), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n369), .B1(new_n379), .B2(new_n367), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n376), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n308), .A2(new_n247), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n360), .A2(new_n361), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(new_n308), .ZN(new_n385));
  OAI211_X1 g184(.A(KEYINPUT74), .B(KEYINPUT5), .C1(new_n385), .C2(new_n369), .ZN(new_n386));
  AOI221_X4 g185(.A(KEYINPUT75), .B1(new_n372), .B2(new_n375), .C1(new_n382), .C2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT75), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(new_n386), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n375), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n371), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(G1gat), .B(G29gat), .Z(new_n393));
  XNOR2_X1  g192(.A(G57gat), .B(G85gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  AND2_X1   g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT6), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n392), .A2(new_n397), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n401));
  INV_X1    g200(.A(new_n397), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n402), .B(new_n371), .C1(new_n387), .C2(new_n391), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT35), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n329), .A2(new_n356), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n329), .A2(KEYINPUT80), .A3(new_n356), .A4(new_n405), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT77), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n403), .A2(new_n410), .A3(new_n401), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n400), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n403), .B2(new_n401), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n399), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n356), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT78), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(KEYINPUT78), .A3(new_n356), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n329), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n408), .A2(new_n409), .B1(new_n419), .B2(KEYINPUT35), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n282), .B(KEYINPUT36), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n352), .A2(new_n355), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT39), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n385), .A2(new_n369), .ZN(new_n424));
  AOI211_X1 g223(.A(new_n423), .B(new_n424), .C1(new_n368), .C2(new_n370), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n368), .A2(new_n423), .A3(new_n370), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n425), .A2(new_n426), .A3(new_n397), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n427), .A2(KEYINPUT40), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n398), .B1(KEYINPUT40), .B2(new_n427), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n422), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n335), .B1(new_n353), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT38), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n345), .A2(new_n346), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n291), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n341), .A2(new_n343), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n435), .B(KEYINPUT37), .C1(new_n436), .C2(new_n291), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n403), .A2(new_n401), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n438), .B(new_n399), .C1(new_n398), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n291), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(KEYINPUT37), .A3(new_n347), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n349), .B1(new_n443), .B2(new_n433), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n430), .B(new_n327), .C1(new_n440), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n421), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n417), .A2(new_n418), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(new_n328), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n420), .A2(new_n448), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n331), .A2(G57gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n331), .A2(G57gat), .ZN(new_n451));
  INV_X1    g250(.A(G71gat), .ZN(new_n452));
  INV_X1    g251(.A(G78gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI22_X1  g253(.A1(new_n450), .A2(new_n451), .B1(new_n454), .B2(KEYINPUT9), .ZN(new_n455));
  XNOR2_X1  g254(.A(G71gat), .B(G78gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT21), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n461));
  XOR2_X1   g260(.A(new_n460), .B(new_n461), .Z(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  XOR2_X1   g262(.A(G15gat), .B(G22gat), .Z(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G1gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466));
  INV_X1    g265(.A(G1gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(KEYINPUT16), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(KEYINPUT85), .A3(G8gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(KEYINPUT85), .A2(G8gat), .ZN(new_n471));
  OR2_X1    g270(.A1(KEYINPUT85), .A2(G8gat), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n465), .A2(new_n468), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n458), .B2(new_n459), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(G183gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT88), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n475), .B(new_n211), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AND4_X1   g279(.A1(G231gat), .A2(new_n477), .A3(new_n480), .A4(G233gat), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n477), .A2(new_n480), .B1(G231gat), .B2(G233gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(G127gat), .B(G155gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(new_n286), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n484), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n477), .A2(new_n480), .ZN(new_n487));
  NAND2_X1  g286(.A1(G231gat), .A2(G233gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n477), .A2(new_n480), .A3(G231gat), .A4(G233gat), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n463), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n484), .B1(new_n481), .B2(new_n482), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n489), .A2(new_n490), .A3(new_n486), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n462), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G190gat), .B(G218gat), .Z(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(KEYINPUT91), .ZN(new_n498));
  INV_X1    g297(.A(G43gat), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n499), .A2(G50gat), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT15), .B1(new_n499), .B2(G50gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n499), .A2(G50gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT83), .B(G50gat), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(G43gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT15), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(G29gat), .A2(G36gat), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n508), .B(KEYINPUT14), .Z(new_n509));
  XOR2_X1   g308(.A(KEYINPUT82), .B(G36gat), .Z(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(KEYINPUT84), .A3(G29gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(G29gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT84), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n507), .A2(new_n509), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(new_n512), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n502), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT17), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n520));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521));
  INV_X1    g320(.A(G85gat), .ZN(new_n522));
  AOI22_X1  g321(.A1(KEYINPUT8), .A2(new_n521), .B1(new_n522), .B2(new_n333), .ZN(new_n523));
  NAND2_X1  g322(.A1(KEYINPUT89), .A2(KEYINPUT7), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(new_n522), .B2(new_n333), .ZN(new_n525));
  NAND4_X1  g324(.A1(KEYINPUT89), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G99gat), .B(G106gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n520), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n525), .A2(new_n526), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n531), .A2(KEYINPUT90), .A3(new_n528), .A4(new_n523), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n527), .A2(new_n529), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n498), .B1(new_n519), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n533), .A3(new_n534), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G134gat), .B(G162gat), .Z(new_n540));
  OR2_X1    g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n497), .A2(KEYINPUT91), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT41), .ZN(new_n544));
  INV_X1    g343(.A(G232gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n545), .B2(new_n258), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n543), .B(new_n546), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n541), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n547), .B1(new_n541), .B2(new_n542), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n496), .A2(new_n550), .A3(KEYINPUT92), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT92), .B1(new_n496), .B2(new_n550), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n449), .A2(new_n553), .ZN(new_n554));
  AOI211_X1 g353(.A(new_n500), .B(new_n501), .C1(new_n509), .C2(new_n512), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n514), .A2(new_n509), .A3(new_n511), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(new_n507), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT87), .B1(new_n557), .B2(new_n474), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT87), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n518), .A2(new_n559), .A3(new_n470), .A4(new_n473), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n518), .A2(KEYINPUT17), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n563), .B1(new_n515), .B2(new_n517), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n474), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT86), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n561), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n557), .A2(new_n474), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n561), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n567), .B(KEYINPUT13), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n561), .A2(new_n565), .A3(KEYINPUT18), .A4(new_n568), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G113gat), .B(G141gat), .Z(new_n578));
  XNOR2_X1  g377(.A(G169gat), .B(G197gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT81), .B(KEYINPUT11), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT12), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n571), .A2(new_n575), .A3(new_n576), .A4(new_n583), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n535), .A2(new_n458), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT10), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n531), .A2(new_n591), .A3(new_n523), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n527), .A2(KEYINPUT93), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n593), .A3(new_n529), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n533), .A2(new_n457), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n589), .A2(new_n590), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n533), .A2(new_n457), .A3(KEYINPUT10), .A4(new_n534), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G230gat), .A2(G233gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT94), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n589), .A2(new_n595), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G176gat), .B(G204gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT95), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G120gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G148gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n604), .B(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n588), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n554), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n414), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n414), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(new_n467), .ZN(G1324gat));
  OAI21_X1  g417(.A(G8gat), .B1(new_n611), .B2(new_n356), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT97), .ZN(new_n620));
  NOR2_X1   g419(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n611), .A2(new_n356), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT42), .ZN(new_n623));
  NAND2_X1  g422(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n623), .B1(new_n622), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n620), .B1(new_n625), .B2(new_n626), .ZN(G1325gat));
  INV_X1    g426(.A(G15gat), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n611), .A2(new_n628), .A3(new_n421), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n554), .A2(new_n610), .A3(new_n282), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n628), .B2(new_n630), .ZN(G1326gat));
  XNOR2_X1  g430(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n611), .A2(new_n327), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n611), .B2(new_n327), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT43), .B(G22gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(G1327gat));
  INV_X1    g436(.A(new_n550), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n492), .A2(new_n495), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n610), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n449), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n642), .A2(G29gat), .A3(new_n616), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT45), .Z(new_n644));
  OAI211_X1 g443(.A(KEYINPUT44), .B(new_n638), .C1(new_n420), .C2(new_n448), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n420), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n414), .A2(KEYINPUT78), .A3(new_n356), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT78), .B1(new_n414), .B2(new_n356), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n328), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT100), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n653), .B(new_n328), .C1(new_n649), .C2(new_n650), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n446), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n648), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI211_X1 g456(.A(KEYINPUT101), .B(new_n446), .C1(new_n652), .C2(new_n654), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n647), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n638), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n646), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n641), .ZN(new_n663));
  OAI21_X1  g462(.A(G29gat), .B1(new_n663), .B2(new_n616), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n644), .A2(new_n664), .ZN(G1328gat));
  OAI21_X1  g464(.A(new_n510), .B1(new_n663), .B2(new_n356), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n642), .A2(new_n510), .A3(new_n356), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT46), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(G1329gat));
  NAND2_X1  g468(.A1(KEYINPUT102), .A2(KEYINPUT47), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n499), .B1(new_n642), .B2(new_n283), .ZN(new_n671));
  INV_X1    g470(.A(new_n421), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(G43gat), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n670), .B(new_n671), .C1(new_n663), .C2(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(KEYINPUT102), .A2(KEYINPUT47), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1330gat));
  INV_X1    g475(.A(KEYINPUT48), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n653), .B1(new_n447), .B2(new_n328), .ZN(new_n678));
  INV_X1    g477(.A(new_n654), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n656), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT101), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n655), .A2(new_n648), .A3(new_n656), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n420), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n661), .B1(new_n683), .B2(new_n550), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n327), .A2(new_n504), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n684), .A2(new_n641), .A3(new_n645), .A4(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n504), .B1(new_n642), .B2(new_n327), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n677), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n659), .B2(new_n638), .ZN(new_n692));
  INV_X1    g491(.A(new_n685), .ZN(new_n693));
  NOR4_X1   g492(.A1(new_n692), .A2(new_n640), .A3(new_n646), .A4(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n688), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT103), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(KEYINPUT48), .A3(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n691), .A2(new_n698), .ZN(G1331gat));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n587), .ZN(new_n700));
  INV_X1    g499(.A(new_n609), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n551), .A2(new_n552), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n615), .B(KEYINPUT104), .Z(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g506(.A1(new_n703), .A2(new_n356), .ZN(new_n708));
  NOR2_X1   g507(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n709));
  AND2_X1   g508(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n708), .B2(new_n709), .ZN(G1333gat));
  NAND4_X1  g511(.A1(new_n700), .A2(G71gat), .A3(new_n672), .A4(new_n702), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n282), .B(KEYINPUT105), .Z(new_n714));
  NAND4_X1  g513(.A1(new_n659), .A2(new_n588), .A3(new_n702), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n452), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT107), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n719));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n713), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n719), .B1(new_n718), .B2(new_n721), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(G1334gat));
  NOR2_X1   g523(.A1(new_n703), .A2(new_n327), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(new_n453), .ZN(G1335gat));
  NOR2_X1   g525(.A1(new_n496), .A2(new_n587), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n659), .A2(new_n638), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n609), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n522), .B1(new_n731), .B2(new_n616), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n662), .A2(new_n609), .A3(new_n727), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(G85gat), .A3(new_n615), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n732), .A2(new_n734), .ZN(G1336gat));
  NAND4_X1  g534(.A1(new_n662), .A2(new_n609), .A3(new_n422), .A4(new_n727), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G92gat), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n356), .A2(G92gat), .A3(new_n701), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n730), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n728), .A2(new_n742), .A3(KEYINPUT51), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT51), .B1(new_n728), .B2(new_n742), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n738), .B(KEYINPUT108), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n745), .A2(new_n746), .B1(new_n736), .B2(G92gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n741), .B1(new_n747), .B2(new_n740), .ZN(G1337gat));
  AND2_X1   g547(.A1(new_n733), .A2(G99gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n609), .A3(new_n282), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n749), .A2(new_n672), .B1(new_n270), .B2(new_n750), .ZN(G1338gat));
  INV_X1    g550(.A(KEYINPUT53), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n327), .A2(G106gat), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n731), .B2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n662), .A2(new_n609), .A3(new_n328), .A4(new_n727), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(G106gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n609), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n745), .A2(new_n759), .B1(new_n756), .B2(G106gat), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n755), .A2(new_n757), .B1(new_n760), .B2(new_n752), .ZN(G1339gat));
  INV_X1    g560(.A(KEYINPUT92), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n639), .B2(new_n638), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n496), .A2(new_n550), .A3(KEYINPUT92), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n763), .A2(new_n588), .A3(new_n701), .A4(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n553), .A2(KEYINPUT110), .A3(new_n588), .A4(new_n701), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT111), .B1(new_n598), .B2(new_n601), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n602), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n596), .A2(new_n773), .A3(new_n600), .A4(new_n597), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n774), .A2(KEYINPUT54), .B1(new_n598), .B2(new_n601), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n608), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n604), .A2(new_n608), .ZN(new_n779));
  OAI211_X1 g578(.A(KEYINPUT55), .B(new_n608), .C1(new_n772), .C2(new_n775), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n573), .A2(new_n574), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n568), .B1(new_n561), .B2(new_n565), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n582), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n586), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n638), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n587), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n609), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n786), .B1(new_n789), .B2(new_n638), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n639), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n769), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n792), .A2(new_n329), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n793), .A2(KEYINPUT112), .A3(new_n705), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT112), .B1(new_n793), .B2(new_n705), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n794), .A2(new_n795), .A3(new_n422), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n241), .A3(new_n587), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n615), .A3(new_n356), .ZN(new_n798));
  OAI21_X1  g597(.A(G113gat), .B1(new_n798), .B2(new_n588), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1340gat));
  NAND3_X1  g599(.A1(new_n796), .A2(new_n239), .A3(new_n609), .ZN(new_n801));
  OAI21_X1  g600(.A(G120gat), .B1(new_n798), .B2(new_n701), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(G1341gat));
  NOR3_X1   g602(.A1(new_n798), .A2(new_n234), .A3(new_n639), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n796), .A2(new_n496), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n234), .ZN(G1342gat));
  NAND3_X1  g605(.A1(new_n796), .A2(new_n232), .A3(new_n638), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n807), .A2(KEYINPUT56), .ZN(new_n808));
  OAI21_X1  g607(.A(G134gat), .B1(new_n798), .B2(new_n550), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(KEYINPUT56), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(G1343gat));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n787), .A2(KEYINPUT113), .A3(new_n788), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT113), .B1(new_n787), .B2(new_n788), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n550), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT114), .B(new_n550), .C1(new_n813), .C2(new_n814), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n786), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n639), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n769), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(KEYINPUT57), .A3(new_n328), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n792), .A2(new_n328), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n821), .A2(KEYINPUT115), .A3(KEYINPUT57), .A4(new_n328), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n824), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n421), .A2(new_n356), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n616), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n587), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n812), .B1(new_n832), .B2(G141gat), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n327), .B1(new_n769), .B2(new_n791), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n834), .A2(new_n356), .A3(new_n421), .A4(new_n705), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(G141gat), .A3(new_n588), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n832), .B2(G141gat), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n833), .A2(new_n837), .A3(KEYINPUT58), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839));
  AOI221_X4 g638(.A(new_n836), .B1(new_n812), .B2(new_n839), .C1(new_n832), .C2(G141gat), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n838), .A2(new_n840), .ZN(G1344gat));
  NAND3_X1  g640(.A1(new_n829), .A2(new_n609), .A3(new_n831), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(G148gat), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n825), .A2(KEYINPUT57), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT119), .B1(new_n830), .B2(new_n616), .ZN(new_n848));
  INV_X1    g647(.A(new_n765), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n496), .B1(new_n815), .B2(new_n786), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n826), .B(new_n328), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n701), .B1(new_n831), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n847), .A2(new_n848), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G148gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n854), .A2(new_n855), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT59), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n842), .A2(KEYINPUT118), .A3(new_n843), .A4(G148gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n846), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n835), .A2(G148gat), .A3(new_n701), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT117), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(G1345gat));
  NAND4_X1  g663(.A1(new_n829), .A2(G155gat), .A3(new_n496), .A4(new_n831), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n294), .B1(new_n835), .B2(new_n639), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(G1346gat));
  NOR2_X1   g666(.A1(new_n835), .A2(new_n550), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n829), .A2(new_n638), .A3(new_n831), .ZN(new_n869));
  XNOR2_X1  g668(.A(KEYINPUT71), .B(G162gat), .ZN(new_n870));
  MUX2_X1   g669(.A(new_n868), .B(new_n869), .S(new_n870), .Z(G1347gat));
  NOR2_X1   g670(.A1(new_n615), .A2(new_n356), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n793), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n205), .A3(new_n587), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n705), .A2(new_n356), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n327), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n792), .A2(new_n714), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n877), .A2(new_n878), .A3(new_n588), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n875), .B1(new_n205), .B2(new_n879), .ZN(G1348gat));
  OAI21_X1  g679(.A(new_n206), .B1(new_n873), .B2(new_n701), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT121), .Z(new_n882));
  NOR2_X1   g681(.A1(new_n877), .A2(new_n878), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n701), .A2(new_n206), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(G1349gat));
  AOI21_X1  g684(.A(new_n211), .B1(new_n883), .B2(new_n496), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n496), .A2(new_n223), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n874), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g688(.A(new_n212), .B1(new_n883), .B2(new_n638), .ZN(new_n890));
  XNOR2_X1  g689(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n890), .B(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n212), .A3(new_n638), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1351gat));
  AND2_X1   g693(.A1(new_n847), .A2(new_n851), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n421), .A3(new_n876), .ZN(new_n896));
  OR3_X1    g695(.A1(new_n896), .A2(KEYINPUT124), .A3(new_n588), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT124), .B1(new_n896), .B2(new_n588), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(G197gat), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n834), .A2(new_n421), .A3(new_n872), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n900), .B(KEYINPUT123), .Z(new_n901));
  INV_X1    g700(.A(G197gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n902), .A3(new_n587), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n899), .A2(new_n903), .ZN(G1352gat));
  AND2_X1   g703(.A1(new_n895), .A2(new_n876), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n905), .A2(new_n906), .A3(new_n609), .A4(new_n421), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT127), .B1(new_n896), .B2(new_n701), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(G204gat), .A3(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n900), .A2(G204gat), .A3(new_n701), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(KEYINPUT125), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(KEYINPUT125), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT126), .B1(new_n913), .B2(KEYINPUT62), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(KEYINPUT62), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n911), .A2(new_n912), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n909), .A2(new_n914), .A3(new_n915), .A4(new_n918), .ZN(G1353gat));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n286), .A3(new_n496), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n421), .A3(new_n496), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n922));
  OAI211_X1 g721(.A(KEYINPUT63), .B(G211gat), .C1(new_n896), .C2(new_n639), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n920), .B1(new_n922), .B2(new_n924), .ZN(G1354gat));
  OAI21_X1  g724(.A(G218gat), .B1(new_n896), .B2(new_n550), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n901), .A2(new_n287), .A3(new_n638), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1355gat));
endmodule


