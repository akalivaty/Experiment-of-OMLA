//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G227), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT81), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(KEYINPUT3), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT82), .A2(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT82), .A2(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT83), .B1(new_n197), .B2(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT83), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(new_n192), .A3(G107), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT85), .B(KEYINPUT4), .Z(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(G101), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  OR2_X1    g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n208), .B2(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n206), .A2(KEYINPUT64), .A3(G143), .ZN(new_n216));
  INV_X1    g030(.A(new_n211), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n209), .A4(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n205), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n196), .A2(new_n201), .A3(new_n221), .A4(new_n202), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(G104), .B2(new_n197), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT82), .A2(G107), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT82), .A2(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n225), .B1(new_n228), .B2(new_n193), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n221), .B1(new_n229), .B2(new_n201), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT84), .B1(new_n223), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n232));
  AOI21_X1  g046(.A(G101), .B1(new_n198), .B2(new_n200), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n203), .A2(G101), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT84), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n220), .B1(new_n231), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(G104), .B1(new_n194), .B2(new_n195), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n192), .A2(G107), .ZN(new_n240));
  OAI21_X1  g054(.A(G101), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n222), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT1), .ZN(new_n245));
  AND4_X1   g059(.A1(new_n215), .A2(new_n216), .A3(new_n245), .A4(new_n209), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT1), .B1(new_n208), .B2(G146), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n247), .A2(G128), .B1(new_n207), .B2(new_n209), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT10), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n243), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n215), .A2(new_n216), .A3(new_n209), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n247), .A2(G128), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n215), .A2(new_n216), .A3(new_n245), .A4(new_n209), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n222), .A3(new_n241), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n250), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n238), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(G137), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(G137), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT11), .A3(G134), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G131), .ZN(new_n269));
  INV_X1    g083(.A(G131), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n264), .A2(new_n267), .A3(new_n270), .A4(new_n265), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n191), .B1(new_n261), .B2(new_n273), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n257), .A2(new_n222), .A3(new_n241), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n254), .A2(new_n210), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n256), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n222), .B2(new_n241), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n272), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT12), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n242), .A2(new_n249), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n258), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT12), .A3(new_n272), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT87), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT12), .B1(new_n283), .B2(new_n272), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n280), .B(new_n273), .C1(new_n282), .C2(new_n258), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT87), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n274), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT88), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT86), .B1(new_n238), .B2(new_n260), .ZN(new_n293));
  INV_X1    g107(.A(new_n220), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n236), .B1(new_n234), .B2(new_n235), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n243), .A2(new_n251), .B1(new_n258), .B2(new_n250), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(new_n300), .A3(new_n272), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n261), .A2(new_n273), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n191), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n288), .B1(new_n286), .B2(new_n287), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n281), .A2(KEYINPUT87), .A3(new_n284), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT88), .A3(new_n274), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n292), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G469), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n281), .A2(new_n284), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n302), .A2(new_n314), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n315), .A2(new_n191), .B1(new_n301), .B2(new_n274), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n313), .B1(new_n316), .B2(G469), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT9), .B(G234), .ZN(new_n319));
  OAI21_X1  g133(.A(G221), .B1(new_n319), .B2(G902), .ZN(new_n320));
  XOR2_X1   g134(.A(G128), .B(G143), .Z(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(G134), .ZN(new_n322));
  INV_X1    g136(.A(G122), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G116), .ZN(new_n324));
  INV_X1    g138(.A(G116), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G122), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n228), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(KEYINPUT14), .A3(G122), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n326), .ZN(new_n329));
  OAI211_X1 g143(.A(G107), .B(new_n328), .C1(new_n329), .C2(KEYINPUT14), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n322), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  OR3_X1    g145(.A1(new_n321), .A2(KEYINPUT99), .A3(G134), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n329), .B1(new_n227), .B2(new_n226), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n327), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT99), .B1(new_n321), .B2(G134), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT13), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n208), .A3(G128), .ZN(new_n337));
  OAI211_X1 g151(.A(G134), .B(new_n337), .C1(new_n321), .C2(new_n336), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n332), .A2(new_n334), .A3(new_n335), .A4(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G217), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n319), .A2(new_n340), .A3(G953), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n331), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(new_n331), .B2(new_n339), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n311), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G478), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(KEYINPUT15), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n344), .B(new_n346), .Z(new_n347));
  INV_X1    g161(.A(G125), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n348), .A2(KEYINPUT16), .A3(G140), .ZN(new_n349));
  XNOR2_X1  g163(.A(G125), .B(G140), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(new_n350), .B2(KEYINPUT16), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G146), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n351), .A2(G146), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G237), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n187), .A3(G214), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n208), .ZN(new_n358));
  NOR2_X1   g172(.A1(G237), .A2(G953), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(G143), .A3(G214), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT17), .A3(G131), .ZN(new_n362));
  AND4_X1   g176(.A1(G143), .A2(new_n356), .A3(new_n187), .A4(G214), .ZN(new_n363));
  AOI21_X1  g177(.A(G143), .B1(new_n359), .B2(G214), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n270), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(G131), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n355), .B(new_n362), .C1(KEYINPUT17), .C2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G140), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G125), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n348), .A2(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT75), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n350), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n376), .A3(new_n206), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(G146), .ZN(new_n378));
  NAND2_X1  g192(.A1(KEYINPUT18), .A2(G131), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n377), .A2(new_n378), .B1(new_n365), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT97), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT96), .B1(new_n363), .B2(new_n364), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT96), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n358), .A2(new_n383), .A3(new_n360), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n379), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n381), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI211_X1 g201(.A(KEYINPUT97), .B(new_n379), .C1(new_n382), .C2(new_n384), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n380), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G113), .B(G122), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n192), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n369), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n369), .B2(new_n389), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n311), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G475), .ZN(new_n396));
  NOR2_X1   g210(.A1(G475), .A2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n377), .A2(new_n378), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n365), .A2(new_n379), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT96), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n383), .B1(new_n358), .B2(new_n360), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n386), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT97), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n385), .A2(new_n381), .A3(new_n386), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n401), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n366), .A2(new_n367), .B1(G146), .B2(new_n351), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n373), .A2(KEYINPUT19), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n374), .A2(new_n376), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n206), .B(new_n409), .C1(new_n410), .C2(KEYINPUT19), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT98), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n391), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT98), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n389), .A2(new_n416), .A3(new_n412), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  AOI211_X1 g232(.A(KEYINPUT20), .B(new_n398), .C1(new_n418), .C2(new_n392), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n415), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n416), .B1(new_n389), .B2(new_n412), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n392), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n420), .B1(new_n423), .B2(new_n397), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n347), .B(new_n396), .C1(new_n419), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(G234), .A2(G237), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n426), .A2(G952), .A3(new_n187), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n426), .A2(G902), .A3(G953), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(G898), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n318), .A2(new_n320), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G122), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n433), .B(KEYINPUT89), .Z(new_n434));
  INV_X1    g248(.A(G119), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G116), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n325), .A2(G119), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT2), .B(G113), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT66), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT66), .ZN(new_n442));
  INV_X1    g256(.A(G113), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT2), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT2), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G113), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G116), .B(G119), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n442), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n440), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n205), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n231), .B2(new_n237), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT66), .B1(new_n438), .B2(new_n439), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n447), .A2(new_n448), .A3(new_n442), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT5), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n435), .A3(G116), .ZN(new_n457));
  OAI211_X1 g271(.A(G113), .B(new_n457), .C1(new_n438), .C2(new_n456), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n455), .A2(new_n222), .A3(new_n241), .A4(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n434), .B1(new_n452), .B2(new_n460), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n230), .A2(new_n204), .B1(new_n455), .B2(new_n440), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n295), .B2(new_n296), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n459), .A3(new_n433), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n464), .A3(KEYINPUT6), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n213), .A2(new_n218), .ZN(new_n466));
  AOI21_X1  g280(.A(G125), .B1(new_n254), .B2(new_n210), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n466), .A2(G125), .B1(new_n467), .B2(new_n256), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n187), .A2(G224), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n463), .A2(new_n459), .ZN(new_n472));
  INV_X1    g286(.A(new_n434), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n473), .A2(KEYINPUT6), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n471), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  AOI211_X1 g290(.A(KEYINPUT90), .B(new_n474), .C1(new_n463), .C2(new_n459), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n465), .B(new_n470), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n433), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n452), .A2(new_n460), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT92), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n469), .B1(KEYINPUT91), .B2(KEYINPUT7), .ZN(new_n482));
  AND2_X1   g296(.A1(KEYINPUT91), .A2(KEYINPUT7), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n481), .B1(new_n468), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n484), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n276), .A2(new_n348), .A3(new_n256), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n348), .B1(new_n213), .B2(new_n218), .ZN(new_n489));
  OAI211_X1 g303(.A(KEYINPUT92), .B(new_n486), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n433), .B(KEYINPUT8), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n455), .A2(new_n458), .B1(new_n222), .B2(new_n241), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n492), .B1(new_n460), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT93), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n469), .A2(KEYINPUT7), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n495), .B1(new_n497), .B2(new_n489), .ZN(new_n498));
  INV_X1    g312(.A(new_n489), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n499), .A2(KEYINPUT93), .A3(new_n487), .A4(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n491), .A2(new_n494), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(KEYINPUT94), .B(new_n311), .C1(new_n480), .C2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n455), .A2(new_n458), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n242), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n459), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n507), .A2(new_n492), .B1(new_n498), .B2(new_n500), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n464), .A2(new_n491), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT94), .B1(new_n509), .B2(new_n311), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n478), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G210), .B1(G237), .B2(G902), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n478), .B(new_n512), .C1(new_n504), .C2(new_n510), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(KEYINPUT95), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G214), .B1(G237), .B2(G902), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n311), .B1(new_n480), .B2(new_n502), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT94), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n503), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n512), .B1(new_n521), .B2(new_n478), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT95), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n516), .A2(new_n517), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n432), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n340), .B1(G234), .B2(new_n311), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n352), .A2(new_n377), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT73), .B1(new_n435), .B2(G128), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT73), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n244), .A3(G119), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n435), .A2(G128), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT24), .B(G110), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT74), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT23), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n435), .B2(G128), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n244), .A2(KEYINPUT23), .A3(G119), .ZN(new_n539));
  INV_X1    g353(.A(G110), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n532), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n536), .B1(new_n535), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n528), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n533), .A2(new_n534), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n532), .A3(new_n539), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G110), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n545), .B(new_n547), .C1(new_n353), .C2(new_n354), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT77), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT22), .B(G137), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n544), .A2(new_n548), .A3(new_n549), .A4(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n544), .A2(new_n548), .A3(new_n552), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT77), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n552), .B(KEYINPUT76), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n544), .B2(new_n548), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n553), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n558), .A2(KEYINPUT25), .A3(new_n311), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT25), .B1(new_n558), .B2(new_n311), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n527), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT79), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n527), .A2(G902), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n563), .B(KEYINPUT78), .Z(new_n564));
  AND3_X1   g378(.A1(new_n558), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n562), .B1(new_n558), .B2(new_n564), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT80), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n561), .A2(new_n567), .A3(KEYINPUT80), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(G472), .A2(G902), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n359), .A2(G210), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT27), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT26), .B(G101), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n577), .B(KEYINPUT68), .Z(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT28), .ZN(new_n580));
  INV_X1    g394(.A(new_n450), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n266), .A2(G134), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n263), .A2(G137), .ZN(new_n583));
  OAI21_X1  g397(.A(G131), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n584), .B(new_n271), .C1(new_n246), .C2(new_n248), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n585), .A2(KEYINPUT65), .B1(new_n219), .B2(new_n272), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n271), .A2(new_n584), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT65), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n277), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n581), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT69), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n219), .A2(new_n272), .B1(new_n587), .B2(new_n277), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT67), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n455), .A2(new_n593), .A3(new_n440), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n455), .B2(new_n440), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n590), .A2(new_n591), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n271), .A2(new_n584), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT65), .B1(new_n249), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n219), .A2(new_n272), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n589), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n450), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT69), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n580), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n450), .A2(KEYINPUT67), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n455), .A2(new_n593), .A3(new_n440), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n592), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n580), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(KEYINPUT70), .B(new_n579), .C1(new_n604), .C2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT30), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n601), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n592), .A2(KEYINPUT30), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n450), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n607), .A3(new_n577), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT31), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n614), .A2(KEYINPUT31), .A3(new_n607), .A4(new_n577), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n610), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n601), .A2(new_n591), .A3(new_n450), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n607), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n591), .B1(new_n601), .B2(new_n450), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT28), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n578), .B1(new_n624), .B2(new_n608), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(KEYINPUT70), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n573), .B1(new_n620), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT32), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT70), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n603), .A2(new_n607), .A3(new_n621), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n609), .B1(new_n630), .B2(KEYINPUT28), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n629), .B1(new_n631), .B2(new_n578), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n619), .A3(new_n610), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT32), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n634), .A3(new_n573), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n605), .A2(new_n606), .ZN(new_n637));
  INV_X1    g451(.A(new_n592), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n580), .B1(new_n639), .B2(new_n607), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n609), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n577), .A2(KEYINPUT29), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT71), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n607), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n592), .B1(new_n605), .B2(new_n606), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT28), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n646), .A2(KEYINPUT71), .A3(new_n608), .A4(new_n642), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n311), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT72), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n631), .A2(new_n578), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n614), .A2(new_n607), .ZN(new_n651));
  INV_X1    g465(.A(new_n577), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT29), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n646), .A2(new_n608), .A3(new_n642), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT71), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT72), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n658), .A3(new_n311), .A4(new_n647), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n649), .A2(new_n654), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(G472), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n572), .B1(new_n636), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n526), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G101), .ZN(G3));
  NAND2_X1  g478(.A1(new_n633), .A2(new_n311), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n665), .A2(G472), .B1(new_n573), .B2(new_n633), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n561), .A2(KEYINPUT80), .A3(new_n567), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT80), .B1(new_n561), .B2(new_n567), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n320), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n312), .B2(new_n317), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n515), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n517), .B1(new_n674), .B2(new_n522), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n396), .B1(new_n419), .B2(new_n424), .ZN(new_n676));
  INV_X1    g490(.A(new_n430), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n331), .A2(new_n339), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT33), .ZN(new_n681));
  OR3_X1    g495(.A1(new_n681), .A2(new_n342), .A3(new_n343), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n681), .B1(new_n342), .B2(new_n343), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n345), .A2(G902), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n344), .A2(new_n686), .A3(new_n345), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n686), .B1(new_n344), .B2(new_n345), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n676), .A2(new_n677), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT102), .B1(new_n675), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n690), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  INV_X1    g507(.A(new_n517), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n514), .B2(new_n515), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n673), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT34), .B(G104), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G6));
  NOR3_X1   g514(.A1(new_n676), .A2(new_n430), .A3(new_n347), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n675), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n673), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT35), .B(G107), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G9));
  AOI22_X1  g520(.A1(new_n625), .A2(KEYINPUT70), .B1(new_n617), .B2(new_n618), .ZN(new_n707));
  AOI21_X1  g521(.A(G902), .B1(new_n707), .B2(new_n632), .ZN(new_n708));
  INV_X1    g522(.A(G472), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n627), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n544), .A2(new_n548), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT103), .ZN(new_n712));
  INV_X1    g526(.A(new_n556), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n712), .A2(KEYINPUT36), .A3(new_n713), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n713), .A2(KEYINPUT36), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n564), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n561), .A2(new_n717), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n432), .A2(new_n525), .A3(new_n710), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT37), .B(G110), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G12));
  INV_X1    g535(.A(new_n573), .ZN(new_n722));
  AOI211_X1 g536(.A(KEYINPUT32), .B(new_n722), .C1(new_n707), .C2(new_n632), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n634), .B1(new_n633), .B2(new_n573), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n661), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n675), .A2(new_n718), .ZN(new_n726));
  INV_X1    g540(.A(G900), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n427), .B1(new_n428), .B2(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n676), .A2(new_n347), .A3(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n725), .A2(new_n726), .A3(new_n671), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G128), .ZN(G30));
  NOR2_X1   g545(.A1(new_n644), .A2(new_n645), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n615), .B1(new_n732), .B2(new_n578), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n733), .A2(new_n311), .ZN(new_n734));
  OAI22_X1  g548(.A1(new_n723), .A2(new_n724), .B1(new_n709), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT104), .ZN(new_n736));
  INV_X1    g550(.A(new_n347), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n676), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n738), .A2(new_n739), .A3(new_n517), .A4(new_n718), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n676), .A2(new_n737), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n561), .A2(new_n717), .A3(new_n517), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT105), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n728), .B(KEYINPUT39), .Z(new_n745));
  NAND2_X1  g559(.A1(new_n671), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n744), .B1(KEYINPUT40), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n516), .A2(new_n524), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n748), .B(KEYINPUT38), .Z(new_n749));
  OR2_X1    g563(.A1(new_n746), .A2(KEYINPUT40), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n736), .A2(new_n747), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G143), .ZN(G45));
  INV_X1    g566(.A(new_n718), .ZN(new_n753));
  INV_X1    g567(.A(new_n728), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n676), .A2(new_n689), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n671), .A2(new_n695), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT106), .A3(new_n725), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n671), .A2(new_n695), .A3(new_n753), .A4(new_n756), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n628), .A2(new_n635), .B1(G472), .B2(new_n660), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT107), .B(G146), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G48));
  INV_X1    g579(.A(new_n662), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n307), .A2(KEYINPUT88), .A3(new_n274), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT88), .B1(new_n307), .B2(new_n274), .ZN(new_n769));
  INV_X1    g583(.A(new_n191), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n301), .B2(new_n302), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n767), .B1(new_n772), .B2(G902), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n309), .A2(KEYINPUT108), .A3(new_n311), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(G469), .A3(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n312), .A2(new_n320), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n766), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n697), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT41), .B(G113), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(G15));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n703), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G116), .ZN(G18));
  NAND2_X1  g597(.A1(new_n725), .A2(new_n431), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n775), .A2(new_n776), .A3(new_n695), .A4(new_n753), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G119), .ZN(G21));
  NOR2_X1   g601(.A1(new_n741), .A2(new_n430), .ZN(new_n788));
  AND4_X1   g602(.A1(new_n695), .A2(new_n775), .A3(new_n776), .A4(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n579), .B1(new_n640), .B2(new_n609), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n722), .B1(new_n619), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n665), .B2(G472), .ZN(new_n792));
  INV_X1    g606(.A(new_n568), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G122), .ZN(G24));
  INV_X1    g610(.A(KEYINPUT109), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n755), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n676), .A2(KEYINPUT109), .A3(new_n689), .A4(new_n754), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n792), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n785), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n348), .ZN(G27));
  AND2_X1   g616(.A1(new_n798), .A2(new_n799), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n694), .B1(new_n516), .B2(new_n524), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(KEYINPUT42), .A3(new_n671), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n725), .A2(new_n806), .A3(new_n793), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT110), .B1(new_n761), .B2(new_n568), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n725), .A2(new_n669), .A3(new_n671), .A4(new_n804), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT42), .B1(new_n810), .B2(new_n803), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n270), .ZN(G33));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n729), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G134), .ZN(G36));
  OAI211_X1 g629(.A(new_n689), .B(new_n396), .C1(new_n424), .C2(new_n419), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT43), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT111), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n816), .B(new_n817), .C1(new_n818), .C2(new_n676), .ZN(new_n819));
  INV_X1    g633(.A(new_n676), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n820), .B(new_n689), .C1(KEYINPUT111), .C2(KEYINPUT43), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n819), .A2(new_n821), .A3(KEYINPUT112), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n666), .A2(new_n718), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n824), .A2(KEYINPUT44), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT113), .ZN(new_n828));
  INV_X1    g642(.A(new_n804), .ZN(new_n829));
  INV_X1    g643(.A(new_n313), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n316), .A2(KEYINPUT45), .ZN(new_n831));
  OAI21_X1  g645(.A(G469), .B1(new_n316), .B2(KEYINPUT45), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT46), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(KEYINPUT46), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n312), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n320), .A3(new_n745), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT44), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n829), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n828), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G137), .ZN(G39));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n320), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT47), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n837), .A2(KEYINPUT47), .A3(new_n320), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n761), .A2(new_n572), .A3(new_n756), .A4(new_n804), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(new_n370), .ZN(G42));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n775), .A2(new_n312), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n670), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n427), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n819), .B2(new_n821), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n794), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n829), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n852), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n749), .A2(new_n858), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n775), .A2(new_n694), .A3(new_n776), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT118), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT50), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n777), .A2(new_n829), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n669), .A3(new_n427), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n736), .ZN(new_n870));
  INV_X1    g684(.A(new_n689), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n820), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n868), .A2(new_n857), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n792), .A2(new_n753), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n870), .A2(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n861), .B1(new_n867), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n865), .A2(new_n866), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT50), .B1(new_n862), .B2(new_n864), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n876), .B(new_n861), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n860), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT120), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n884), .B(new_n860), .C1(new_n877), .C2(new_n881), .ZN(new_n885));
  INV_X1    g699(.A(new_n807), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n806), .B1(new_n725), .B2(new_n793), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n874), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g702(.A(KEYINPUT121), .B(KEYINPUT48), .Z(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n777), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n695), .ZN(new_n892));
  OAI211_X1 g706(.A(G952), .B(new_n187), .C1(new_n892), .C2(new_n858), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n820), .A2(new_n871), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n870), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n888), .A2(new_n889), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n854), .B(KEYINPUT117), .Z(new_n898));
  INV_X1    g712(.A(new_n848), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n859), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n867), .A2(new_n876), .A3(new_n900), .ZN(new_n901));
  AOI211_X1 g715(.A(new_n890), .B(new_n897), .C1(new_n901), .C2(new_n852), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n883), .A2(new_n885), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT106), .B1(new_n757), .B2(new_n725), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n760), .A2(new_n761), .A3(new_n759), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT116), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n675), .A2(new_n741), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n753), .A2(new_n728), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n735), .A2(new_n909), .A3(new_n910), .A4(new_n671), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n911), .B(new_n730), .C1(new_n785), .C2(new_n800), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n907), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n671), .A2(new_n695), .A3(new_n753), .A4(new_n729), .ZN(new_n914));
  OAI22_X1  g728(.A1(new_n785), .A2(new_n800), .B1(new_n914), .B2(new_n761), .ZN(new_n915));
  INV_X1    g729(.A(new_n911), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT116), .B1(new_n917), .B2(new_n763), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n904), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  OR3_X1    g733(.A1(new_n425), .A2(KEYINPUT115), .A3(new_n728), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT115), .B1(new_n425), .B2(new_n728), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n800), .B1(new_n761), .B2(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n804), .A2(new_n671), .A3(new_n753), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n729), .A2(new_n810), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n809), .B2(new_n811), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT114), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n672), .A2(new_n525), .A3(new_n702), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n719), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n526), .A2(new_n666), .A3(new_n753), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n669), .A2(new_n671), .ZN(new_n931));
  INV_X1    g745(.A(new_n525), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n931), .A2(new_n932), .A3(new_n666), .A4(new_n701), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n930), .A2(new_n933), .A3(KEYINPUT114), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  AOI22_X1  g749(.A1(new_n789), .A2(new_n794), .B1(new_n526), .B2(new_n662), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n673), .A2(new_n932), .A3(new_n692), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n891), .B(new_n662), .C1(new_n697), .C2(new_n703), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n936), .A2(new_n786), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n926), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT52), .B1(new_n907), .B2(new_n912), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n919), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT53), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n908), .B1(new_n907), .B2(new_n912), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n917), .A2(KEYINPUT116), .A3(new_n763), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT52), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n919), .A2(new_n940), .A3(KEYINPUT53), .A4(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT54), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n919), .A2(new_n940), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n943), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT54), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n919), .A2(new_n940), .A3(KEYINPUT53), .A4(new_n941), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n903), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(G952), .A2(G953), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n853), .B(KEYINPUT49), .Z(new_n959));
  NAND3_X1  g773(.A1(new_n793), .A2(new_n517), .A3(new_n320), .ZN(new_n960));
  OR4_X1    g774(.A1(new_n749), .A2(new_n959), .A3(new_n816), .A4(new_n960), .ZN(new_n961));
  OAI22_X1  g775(.A1(new_n957), .A2(new_n958), .B1(new_n736), .B2(new_n961), .ZN(G75));
  AOI21_X1  g776(.A(new_n311), .B1(new_n952), .B2(new_n954), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(G210), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT56), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n465), .B1(new_n476), .B2(new_n477), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(new_n470), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT55), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n964), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n964), .B2(new_n965), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n187), .A2(G952), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(G51));
  INV_X1    g786(.A(KEYINPUT122), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n831), .A2(new_n832), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n963), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n973), .B1(new_n963), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n313), .B(KEYINPUT57), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n953), .B1(new_n952), .B2(new_n954), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n309), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n971), .B1(new_n977), .B2(new_n982), .ZN(G54));
  INV_X1    g797(.A(new_n971), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n952), .A2(new_n954), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(G902), .ZN(new_n986));
  INV_X1    g800(.A(new_n423), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT58), .ZN(new_n988));
  INV_X1    g802(.A(G475), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n984), .B1(new_n986), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n423), .B1(new_n963), .B2(new_n990), .ZN(new_n995));
  OAI21_X1  g809(.A(KEYINPUT123), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n987), .B1(new_n986), .B2(new_n991), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT123), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n971), .B1(new_n963), .B2(new_n992), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n996), .A2(new_n1000), .ZN(G60));
  NAND2_X1  g815(.A1(new_n682), .A2(new_n683), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT124), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G478), .A2(G902), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT59), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n1003), .B(new_n1005), .C1(new_n979), .C2(new_n980), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n984), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1003), .B1(new_n956), .B2(new_n1005), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n1008), .ZN(G63));
  INV_X1    g823(.A(KEYINPUT61), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G217), .A2(G902), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT60), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n952), .B2(new_n954), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n714), .A2(new_n716), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n984), .B1(new_n1013), .B2(new_n558), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1010), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OR2_X1    g832(.A1(new_n1013), .A2(new_n558), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1019), .A2(KEYINPUT61), .A3(new_n984), .A4(new_n1015), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1018), .A2(new_n1020), .ZN(G66));
  INV_X1    g835(.A(G224), .ZN(new_n1022));
  OAI21_X1  g836(.A(G953), .B1(new_n429), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(KEYINPUT125), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n935), .A2(new_n939), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1025), .A2(G953), .ZN(new_n1026));
  MUX2_X1   g840(.A(new_n1024), .B(KEYINPUT125), .S(new_n1026), .Z(new_n1027));
  OAI21_X1  g841(.A(new_n966), .B1(G898), .B2(new_n187), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(G69));
  AOI21_X1  g843(.A(new_n850), .B1(new_n828), .B2(new_n841), .ZN(new_n1030));
  INV_X1    g844(.A(new_n915), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n763), .A2(new_n1031), .A3(new_n814), .ZN(new_n1032));
  INV_X1    g846(.A(new_n909), .ZN(new_n1033));
  AOI211_X1 g847(.A(new_n1033), .B(new_n838), .C1(new_n807), .C2(new_n808), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n812), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1030), .A2(new_n1035), .A3(new_n187), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n612), .A2(new_n613), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n409), .B1(new_n410), .B2(KEYINPUT19), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n1036), .B(new_n1039), .C1(new_n727), .C2(new_n187), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n751), .A2(new_n763), .A3(new_n1031), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT62), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g857(.A1(new_n751), .A2(KEYINPUT62), .A3(new_n763), .A4(new_n1031), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g859(.A(new_n894), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1046), .B1(new_n347), .B2(new_n676), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  OR4_X1    g862(.A1(new_n766), .A2(new_n1048), .A3(new_n746), .A4(new_n829), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1045), .A2(new_n1030), .A3(new_n1049), .ZN(new_n1050));
  AND2_X1   g864(.A1(new_n1050), .A2(new_n187), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1040), .B1(new_n1051), .B2(new_n1039), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1053));
  XNOR2_X1  g867(.A(new_n1052), .B(new_n1053), .ZN(G72));
  NAND2_X1  g868(.A1(new_n651), .A2(new_n577), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n1045), .A2(new_n1025), .A3(new_n1030), .A4(new_n1049), .ZN(new_n1056));
  NAND2_X1  g870(.A1(G472), .A2(G902), .ZN(new_n1057));
  XOR2_X1   g871(.A(new_n1057), .B(KEYINPUT63), .Z(new_n1058));
  AOI21_X1  g872(.A(new_n1055), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n614), .A2(new_n607), .A3(new_n652), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1030), .A2(new_n1035), .A3(new_n1025), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n1060), .B1(new_n1061), .B2(new_n1058), .ZN(new_n1062));
  NOR3_X1   g876(.A1(new_n1059), .A2(new_n971), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g877(.A(KEYINPUT126), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1055), .A2(new_n1060), .A3(new_n1058), .ZN(new_n1065));
  INV_X1    g879(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n1064), .B1(new_n949), .B2(new_n1066), .ZN(new_n1067));
  AOI211_X1 g881(.A(KEYINPUT126), .B(new_n1065), .C1(new_n944), .C2(new_n948), .ZN(new_n1068));
  OAI21_X1  g882(.A(new_n1063), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g883(.A(KEYINPUT127), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g885(.A(new_n1063), .B(KEYINPUT127), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1072));
  NAND2_X1  g886(.A1(new_n1071), .A2(new_n1072), .ZN(G57));
endmodule


