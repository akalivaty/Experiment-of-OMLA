

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(G543), .A2(G651), .ZN(n654) );
  INV_X1 U553 ( .A(n733), .ZN(n710) );
  NOR2_X2 U554 ( .A1(n529), .A2(n528), .ZN(G160) );
  INV_X1 U555 ( .A(KEYINPUT97), .ZN(n728) );
  XNOR2_X1 U556 ( .A(n520), .B(n519), .ZN(n521) );
  NAND2_X1 U557 ( .A1(n733), .A2(G1341), .ZN(n516) );
  NAND2_X1 U558 ( .A1(G8), .A2(n730), .ZN(n517) );
  AND2_X1 U559 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U560 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U561 ( .A1(n740), .A2(G8), .ZN(n743) );
  NOR2_X1 U562 ( .A1(n727), .A2(n726), .ZN(n729) );
  NOR2_X1 U563 ( .A1(G164), .A2(G1384), .ZN(n794) );
  INV_X1 U564 ( .A(KEYINPUT13), .ZN(n573) );
  XNOR2_X1 U565 ( .A(n574), .B(n573), .ZN(n575) );
  INV_X1 U566 ( .A(KEYINPUT64), .ZN(n519) );
  NOR2_X1 U567 ( .A1(n627), .A2(n541), .ZN(n649) );
  NOR2_X1 U568 ( .A1(n627), .A2(G651), .ZN(n650) );
  AND2_X1 U569 ( .A1(G101), .A2(G2104), .ZN(n518) );
  INV_X1 U570 ( .A(G2105), .ZN(n533) );
  NAND2_X1 U571 ( .A1(n518), .A2(n533), .ZN(n520) );
  XNOR2_X1 U572 ( .A(n521), .B(KEYINPUT23), .ZN(n523) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n879) );
  NAND2_X1 U574 ( .A1(G113), .A2(n879), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n523), .A2(n522), .ZN(n529) );
  XNOR2_X1 U576 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n525) );
  NOR2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  XNOR2_X2 U578 ( .A(n525), .B(n524), .ZN(n884) );
  NAND2_X1 U579 ( .A1(G137), .A2(n884), .ZN(n527) );
  NOR2_X4 U580 ( .A1(G2104), .A2(n533), .ZN(n880) );
  NAND2_X1 U581 ( .A1(G125), .A2(n880), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U583 ( .A1(n880), .A2(G126), .ZN(n530) );
  XNOR2_X1 U584 ( .A(n530), .B(KEYINPUT84), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G138), .A2(n884), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n537) );
  AND2_X1 U587 ( .A1(n533), .A2(G2104), .ZN(n883) );
  NAND2_X1 U588 ( .A1(G102), .A2(n883), .ZN(n535) );
  NAND2_X1 U589 ( .A1(G114), .A2(n879), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U591 ( .A1(n537), .A2(n536), .ZN(G164) );
  INV_X1 U592 ( .A(G651), .ZN(n541) );
  NOR2_X1 U593 ( .A1(G543), .A2(n541), .ZN(n538) );
  XOR2_X2 U594 ( .A(KEYINPUT1), .B(n538), .Z(n653) );
  NAND2_X1 U595 ( .A1(G60), .A2(n653), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G85), .A2(n654), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n545) );
  XOR2_X1 U598 ( .A(KEYINPUT0), .B(G543), .Z(n627) );
  NAND2_X1 U599 ( .A1(G72), .A2(n649), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G47), .A2(n650), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U602 ( .A1(n545), .A2(n544), .ZN(G290) );
  XOR2_X1 U603 ( .A(KEYINPUT104), .B(G2446), .Z(n547) );
  XNOR2_X1 U604 ( .A(KEYINPUT105), .B(G2451), .ZN(n546) );
  XNOR2_X1 U605 ( .A(n547), .B(n546), .ZN(n551) );
  XOR2_X1 U606 ( .A(KEYINPUT106), .B(G2435), .Z(n549) );
  XNOR2_X1 U607 ( .A(G2438), .B(G2454), .ZN(n548) );
  XNOR2_X1 U608 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U609 ( .A(n551), .B(n550), .Z(n553) );
  XNOR2_X1 U610 ( .A(G2443), .B(G2427), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n553), .B(n552), .ZN(n556) );
  XNOR2_X1 U612 ( .A(G1348), .B(G2430), .ZN(n554) );
  INV_X1 U613 ( .A(G1341), .ZN(n970) );
  XNOR2_X1 U614 ( .A(n554), .B(n970), .ZN(n555) );
  XOR2_X1 U615 ( .A(n556), .B(n555), .Z(n557) );
  AND2_X1 U616 ( .A1(G14), .A2(n557), .ZN(G401) );
  NAND2_X1 U617 ( .A1(G65), .A2(n653), .ZN(n559) );
  NAND2_X1 U618 ( .A1(G53), .A2(n650), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G91), .A2(n654), .ZN(n561) );
  NAND2_X1 U621 ( .A1(G78), .A2(n649), .ZN(n560) );
  NAND2_X1 U622 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n703) );
  INV_X1 U624 ( .A(n703), .ZN(G299) );
  INV_X1 U625 ( .A(G132), .ZN(G219) );
  NAND2_X1 U626 ( .A1(G94), .A2(G452), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT66), .B(n564), .Z(G173) );
  XOR2_X1 U628 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n566) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n566), .B(n565), .ZN(G223) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n568) );
  INV_X1 U632 ( .A(G223), .ZN(n828) );
  NAND2_X1 U633 ( .A1(G567), .A2(n828), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G234) );
  NAND2_X1 U635 ( .A1(G56), .A2(n653), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n569), .Z(n576) );
  NAND2_X1 U637 ( .A1(G68), .A2(n649), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n654), .A2(G81), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n570), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n574) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n650), .A2(G43), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n961) );
  INV_X1 U644 ( .A(n961), .ZN(n689) );
  NAND2_X1 U645 ( .A1(n689), .A2(G860), .ZN(G153) );
  NAND2_X1 U646 ( .A1(G90), .A2(n654), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G77), .A2(n649), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U649 ( .A(KEYINPUT9), .B(n581), .ZN(n585) );
  NAND2_X1 U650 ( .A1(G64), .A2(n653), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G52), .A2(n650), .ZN(n582) );
  AND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n585), .A2(n584), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U655 ( .A1(G66), .A2(n653), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G92), .A2(n654), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G79), .A2(n649), .ZN(n589) );
  NAND2_X1 U659 ( .A1(G54), .A2(n650), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U662 ( .A(KEYINPUT15), .B(n592), .Z(n897) );
  INV_X1 U663 ( .A(n897), .ZN(n945) );
  INV_X1 U664 ( .A(G868), .ZN(n667) );
  NAND2_X1 U665 ( .A1(n945), .A2(n667), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U667 ( .A1(n654), .A2(G89), .ZN(n595) );
  XNOR2_X1 U668 ( .A(n595), .B(KEYINPUT4), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G76), .A2(n649), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT5), .ZN(n603) );
  NAND2_X1 U672 ( .A1(G63), .A2(n653), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G51), .A2(n650), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U675 ( .A(KEYINPUT6), .B(n601), .Z(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n604), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U678 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U679 ( .A1(G286), .A2(n667), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(G297) );
  INV_X1 U682 ( .A(G559), .ZN(n607) );
  NOR2_X1 U683 ( .A1(G860), .A2(n607), .ZN(n608) );
  XNOR2_X1 U684 ( .A(KEYINPUT71), .B(n608), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n609), .A2(n897), .ZN(n610) );
  XNOR2_X1 U686 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n961), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G868), .A2(n897), .ZN(n611) );
  NOR2_X1 U689 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U690 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G123), .A2(n880), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT18), .ZN(n617) );
  NAND2_X1 U693 ( .A1(G111), .A2(n879), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n615), .B(KEYINPUT72), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G99), .A2(n883), .ZN(n619) );
  NAND2_X1 U697 ( .A1(G135), .A2(n884), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n918) );
  XNOR2_X1 U700 ( .A(n918), .B(G2096), .ZN(n623) );
  INV_X1 U701 ( .A(G2100), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U703 ( .A1(G49), .A2(n650), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n653), .A2(n626), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G87), .A2(n627), .ZN(n628) );
  XOR2_X1 U708 ( .A(KEYINPUT75), .B(n628), .Z(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U710 ( .A1(G88), .A2(n654), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G75), .A2(n649), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U713 ( .A(KEYINPUT78), .B(n633), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G62), .A2(n653), .ZN(n634) );
  XNOR2_X1 U715 ( .A(KEYINPUT77), .B(n634), .ZN(n635) );
  NOR2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n650), .A2(G50), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U719 ( .A(KEYINPUT79), .B(n639), .ZN(G166) );
  NAND2_X1 U720 ( .A1(n654), .A2(G86), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n653), .A2(G61), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U723 ( .A(KEYINPUT76), .B(n642), .ZN(n645) );
  NAND2_X1 U724 ( .A1(G73), .A2(n649), .ZN(n643) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U726 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n650), .A2(G48), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(G305) );
  NAND2_X1 U729 ( .A1(G559), .A2(n897), .ZN(n648) );
  XNOR2_X1 U730 ( .A(n648), .B(n961), .ZN(n908) );
  XNOR2_X1 U731 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n661) );
  NAND2_X1 U732 ( .A1(G80), .A2(n649), .ZN(n652) );
  NAND2_X1 U733 ( .A1(G55), .A2(n650), .ZN(n651) );
  NAND2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n658) );
  NAND2_X1 U735 ( .A1(G67), .A2(n653), .ZN(n656) );
  NAND2_X1 U736 ( .A1(G93), .A2(n654), .ZN(n655) );
  NAND2_X1 U737 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U738 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n659), .B(KEYINPUT74), .ZN(n909) );
  XOR2_X1 U740 ( .A(G288), .B(n909), .Z(n660) );
  XNOR2_X1 U741 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U742 ( .A(G290), .B(n662), .ZN(n664) );
  XNOR2_X1 U743 ( .A(G166), .B(n703), .ZN(n663) );
  XNOR2_X1 U744 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U745 ( .A(n665), .B(G305), .ZN(n896) );
  XNOR2_X1 U746 ( .A(n908), .B(n896), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n666), .A2(G868), .ZN(n669) );
  NAND2_X1 U748 ( .A1(n667), .A2(n909), .ZN(n668) );
  NAND2_X1 U749 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U750 ( .A(KEYINPUT81), .B(n670), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U755 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U756 ( .A(KEYINPUT67), .B(G57), .ZN(G237) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U758 ( .A(KEYINPUT68), .B(G82), .Z(G220) );
  NAND2_X1 U759 ( .A1(G108), .A2(G120), .ZN(n675) );
  NOR2_X1 U760 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U761 ( .A1(G69), .A2(n676), .ZN(n912) );
  NAND2_X1 U762 ( .A1(n912), .A2(G567), .ZN(n682) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U765 ( .A1(G218), .A2(n678), .ZN(n679) );
  XNOR2_X1 U766 ( .A(KEYINPUT82), .B(n679), .ZN(n680) );
  NAND2_X1 U767 ( .A1(n680), .A2(G96), .ZN(n913) );
  NAND2_X1 U768 ( .A1(n913), .A2(G2106), .ZN(n681) );
  NAND2_X1 U769 ( .A1(n682), .A2(n681), .ZN(n832) );
  NAND2_X1 U770 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U771 ( .A1(n832), .A2(n683), .ZN(n684) );
  XOR2_X1 U772 ( .A(KEYINPUT83), .B(n684), .Z(n831) );
  NAND2_X1 U773 ( .A1(n831), .A2(G36), .ZN(G176) );
  INV_X1 U774 ( .A(G166), .ZN(G303) );
  INV_X1 U775 ( .A(G301), .ZN(G171) );
  NAND2_X1 U776 ( .A1(G160), .A2(G40), .ZN(n793) );
  INV_X1 U777 ( .A(n793), .ZN(n685) );
  NAND2_X1 U778 ( .A1(n794), .A2(n685), .ZN(n733) );
  NAND2_X1 U779 ( .A1(G8), .A2(n733), .ZN(n773) );
  NOR2_X1 U780 ( .A1(G1966), .A2(n773), .ZN(n727) );
  NOR2_X1 U781 ( .A1(n710), .A2(G1348), .ZN(n687) );
  NOR2_X1 U782 ( .A1(G2067), .A2(n733), .ZN(n686) );
  NOR2_X1 U783 ( .A1(n687), .A2(n686), .ZN(n693) );
  XOR2_X1 U784 ( .A(G1996), .B(KEYINPUT93), .Z(n1002) );
  NAND2_X1 U785 ( .A1(n710), .A2(n1002), .ZN(n688) );
  XNOR2_X1 U786 ( .A(n688), .B(KEYINPUT26), .ZN(n691) );
  AND2_X1 U787 ( .A1(n516), .A2(n689), .ZN(n690) );
  NAND2_X1 U788 ( .A1(n695), .A2(n897), .ZN(n692) );
  NAND2_X1 U789 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U790 ( .A(n694), .B(KEYINPUT94), .ZN(n697) );
  OR2_X1 U791 ( .A1(n695), .A2(n897), .ZN(n696) );
  NAND2_X1 U792 ( .A1(n697), .A2(n696), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n710), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U794 ( .A(n698), .B(KEYINPUT27), .ZN(n700) );
  XNOR2_X1 U795 ( .A(G1956), .B(KEYINPUT91), .ZN(n971) );
  NOR2_X1 U796 ( .A1(n971), .A2(n710), .ZN(n699) );
  NOR2_X1 U797 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n701) );
  NAND2_X1 U799 ( .A1(n702), .A2(n701), .ZN(n708) );
  NOR2_X1 U800 ( .A1(n704), .A2(n703), .ZN(n706) );
  XOR2_X1 U801 ( .A(KEYINPUT28), .B(KEYINPUT92), .Z(n705) );
  XNOR2_X1 U802 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U804 ( .A(n709), .B(KEYINPUT29), .ZN(n714) );
  OR2_X1 U805 ( .A1(n710), .A2(G1961), .ZN(n712) );
  XNOR2_X1 U806 ( .A(G2078), .B(KEYINPUT25), .ZN(n998) );
  NAND2_X1 U807 ( .A1(n710), .A2(n998), .ZN(n711) );
  NAND2_X1 U808 ( .A1(n712), .A2(n711), .ZN(n716) );
  AND2_X1 U809 ( .A1(G171), .A2(n716), .ZN(n713) );
  XNOR2_X1 U810 ( .A(n715), .B(KEYINPUT95), .ZN(n725) );
  NOR2_X1 U811 ( .A1(G171), .A2(n716), .ZN(n721) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n733), .ZN(n730) );
  NOR2_X1 U813 ( .A1(n730), .A2(n727), .ZN(n717) );
  NAND2_X1 U814 ( .A1(G8), .A2(n717), .ZN(n718) );
  XNOR2_X1 U815 ( .A(KEYINPUT30), .B(n718), .ZN(n719) );
  NOR2_X1 U816 ( .A1(G168), .A2(n719), .ZN(n720) );
  NOR2_X1 U817 ( .A1(n721), .A2(n720), .ZN(n723) );
  XOR2_X1 U818 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n722) );
  XNOR2_X1 U819 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U820 ( .A1(n725), .A2(n724), .ZN(n732) );
  INV_X1 U821 ( .A(n732), .ZN(n726) );
  XNOR2_X1 U822 ( .A(n729), .B(n728), .ZN(n731) );
  NAND2_X1 U823 ( .A1(n731), .A2(n517), .ZN(n747) );
  NAND2_X1 U824 ( .A1(G286), .A2(n732), .ZN(n739) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n773), .ZN(n735) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U827 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U828 ( .A1(n736), .A2(G303), .ZN(n737) );
  XNOR2_X1 U829 ( .A(n737), .B(KEYINPUT98), .ZN(n738) );
  NAND2_X1 U830 ( .A1(n739), .A2(n738), .ZN(n740) );
  INV_X1 U831 ( .A(n743), .ZN(n742) );
  INV_X1 U832 ( .A(KEYINPUT32), .ZN(n741) );
  NAND2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n745) );
  NAND2_X1 U834 ( .A1(KEYINPUT32), .A2(n743), .ZN(n744) );
  NAND2_X1 U835 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n764) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U839 ( .A1(n756), .A2(n748), .ZN(n955) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n752) );
  AND2_X1 U841 ( .A1(n955), .A2(n752), .ZN(n749) );
  NAND2_X1 U842 ( .A1(n764), .A2(n749), .ZN(n754) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n951) );
  INV_X1 U844 ( .A(n773), .ZN(n750) );
  NAND2_X1 U845 ( .A1(n951), .A2(n750), .ZN(n751) );
  NAND2_X1 U846 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U847 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U848 ( .A(n755), .B(KEYINPUT99), .ZN(n761) );
  XNOR2_X1 U849 ( .A(G1981), .B(G305), .ZN(n943) );
  NAND2_X1 U850 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  NOR2_X1 U851 ( .A1(n757), .A2(n773), .ZN(n758) );
  XNOR2_X1 U852 ( .A(KEYINPUT100), .B(n758), .ZN(n759) );
  NOR2_X1 U853 ( .A1(n943), .A2(n759), .ZN(n760) );
  NAND2_X1 U854 ( .A1(n761), .A2(n760), .ZN(n768) );
  NOR2_X1 U855 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U856 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U857 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U858 ( .A1(n773), .A2(n765), .ZN(n766) );
  XOR2_X1 U859 ( .A(KEYINPUT101), .B(n766), .Z(n767) );
  NAND2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U861 ( .A(n769), .B(KEYINPUT102), .ZN(n775) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n770) );
  XOR2_X1 U863 ( .A(n770), .B(KEYINPUT24), .Z(n771) );
  XNOR2_X1 U864 ( .A(KEYINPUT90), .B(n771), .ZN(n772) );
  NOR2_X1 U865 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n810) );
  NAND2_X1 U867 ( .A1(G107), .A2(n879), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G119), .A2(n880), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U870 ( .A(KEYINPUT88), .B(n778), .Z(n782) );
  NAND2_X1 U871 ( .A1(G95), .A2(n883), .ZN(n780) );
  NAND2_X1 U872 ( .A1(G131), .A2(n884), .ZN(n779) );
  AND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n890) );
  AND2_X1 U875 ( .A1(n890), .A2(G1991), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G117), .A2(n879), .ZN(n784) );
  NAND2_X1 U877 ( .A1(G129), .A2(n880), .ZN(n783) );
  NAND2_X1 U878 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U879 ( .A1(G105), .A2(n883), .ZN(n785) );
  XNOR2_X1 U880 ( .A(n785), .B(KEYINPUT89), .ZN(n786) );
  XNOR2_X1 U881 ( .A(n786), .B(KEYINPUT38), .ZN(n787) );
  NOR2_X1 U882 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U883 ( .A1(n884), .A2(G141), .ZN(n789) );
  NAND2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n870) );
  AND2_X1 U885 ( .A1(G1996), .A2(n870), .ZN(n791) );
  NOR2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n926) );
  NOR2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n823) );
  INV_X1 U888 ( .A(n823), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n926), .A2(n795), .ZN(n815) );
  INV_X1 U890 ( .A(n815), .ZN(n808) );
  NAND2_X1 U891 ( .A1(n883), .A2(G104), .ZN(n796) );
  XOR2_X1 U892 ( .A(KEYINPUT85), .B(n796), .Z(n798) );
  NAND2_X1 U893 ( .A1(n884), .A2(G140), .ZN(n797) );
  NAND2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U895 ( .A(KEYINPUT34), .B(n799), .ZN(n805) );
  NAND2_X1 U896 ( .A1(G116), .A2(n879), .ZN(n801) );
  NAND2_X1 U897 ( .A1(G128), .A2(n880), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U899 ( .A(KEYINPUT86), .B(n802), .Z(n803) );
  XNOR2_X1 U900 ( .A(KEYINPUT35), .B(n803), .ZN(n804) );
  NOR2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U902 ( .A(KEYINPUT36), .B(n806), .Z(n861) );
  XOR2_X1 U903 ( .A(KEYINPUT37), .B(G2067), .Z(n820) );
  NAND2_X1 U904 ( .A1(n861), .A2(n820), .ZN(n807) );
  XNOR2_X1 U905 ( .A(KEYINPUT87), .B(n807), .ZN(n937) );
  NAND2_X1 U906 ( .A1(n823), .A2(n937), .ZN(n818) );
  NAND2_X1 U907 ( .A1(n808), .A2(n818), .ZN(n809) );
  NOR2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n812) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n957) );
  NAND2_X1 U910 ( .A1(n957), .A2(n823), .ZN(n811) );
  NAND2_X1 U911 ( .A1(n812), .A2(n811), .ZN(n826) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n870), .ZN(n928) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U914 ( .A1(G1991), .A2(n890), .ZN(n919) );
  NOR2_X1 U915 ( .A1(n813), .A2(n919), .ZN(n814) );
  NOR2_X1 U916 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U917 ( .A1(n928), .A2(n816), .ZN(n817) );
  XNOR2_X1 U918 ( .A(KEYINPUT39), .B(n817), .ZN(n819) );
  NAND2_X1 U919 ( .A1(n819), .A2(n818), .ZN(n821) );
  OR2_X1 U920 ( .A1(n861), .A2(n820), .ZN(n920) );
  NAND2_X1 U921 ( .A1(n821), .A2(n920), .ZN(n822) );
  NAND2_X1 U922 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U923 ( .A(KEYINPUT103), .B(n824), .Z(n825) );
  NAND2_X1 U924 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U925 ( .A(KEYINPUT40), .B(n827), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U928 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U930 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U931 ( .A(n832), .ZN(G319) );
  XOR2_X1 U932 ( .A(KEYINPUT42), .B(G2072), .Z(n834) );
  XNOR2_X1 U933 ( .A(G2084), .B(G2078), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U935 ( .A(n835), .B(G2100), .Z(n837) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2090), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U938 ( .A(G2096), .B(KEYINPUT43), .Z(n839) );
  XNOR2_X1 U939 ( .A(KEYINPUT107), .B(G2678), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n841), .B(n840), .Z(G227) );
  XOR2_X1 U942 ( .A(KEYINPUT109), .B(G1981), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U945 ( .A(n844), .B(KEYINPUT41), .Z(n846) );
  XNOR2_X1 U946 ( .A(G1976), .B(G1971), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U948 ( .A(G1986), .B(G1956), .Z(n848) );
  XNOR2_X1 U949 ( .A(G1966), .B(G1961), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U951 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U952 ( .A(KEYINPUT108), .B(G2474), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G100), .A2(n883), .ZN(n854) );
  NAND2_X1 U955 ( .A1(G112), .A2(n879), .ZN(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n860) );
  NAND2_X1 U957 ( .A1(G136), .A2(n884), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n855), .B(KEYINPUT110), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G124), .A2(n880), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n856), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U962 ( .A1(n860), .A2(n859), .ZN(G162) );
  XNOR2_X1 U963 ( .A(n861), .B(G162), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G103), .A2(n883), .ZN(n863) );
  NAND2_X1 U965 ( .A1(G139), .A2(n884), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G115), .A2(n879), .ZN(n865) );
  NAND2_X1 U968 ( .A1(G127), .A2(n880), .ZN(n864) );
  NAND2_X1 U969 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n914) );
  XNOR2_X1 U972 ( .A(n869), .B(n914), .ZN(n873) );
  XOR2_X1 U973 ( .A(n870), .B(G164), .Z(n871) );
  XNOR2_X1 U974 ( .A(n871), .B(G160), .ZN(n872) );
  XOR2_X1 U975 ( .A(n873), .B(n872), .Z(n878) );
  XOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n875) );
  XNOR2_X1 U977 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U979 ( .A(KEYINPUT111), .B(n876), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n878), .B(n877), .ZN(n894) );
  NAND2_X1 U981 ( .A1(G118), .A2(n879), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G130), .A2(n880), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G106), .A2(n883), .ZN(n886) );
  NAND2_X1 U985 ( .A1(G142), .A2(n884), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U987 ( .A(n887), .B(KEYINPUT45), .Z(n888) );
  NOR2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n918), .B(n892), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U992 ( .A1(G37), .A2(n895), .ZN(G395) );
  XOR2_X1 U993 ( .A(KEYINPUT114), .B(n896), .Z(n899) );
  XNOR2_X1 U994 ( .A(n897), .B(G286), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n901) );
  XOR2_X1 U996 ( .A(n961), .B(G171), .Z(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U998 ( .A1(G37), .A2(n902), .ZN(G397) );
  NOR2_X1 U999 ( .A1(G227), .A2(G229), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(KEYINPUT49), .B(n903), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(G401), .A2(n904), .ZN(n905) );
  AND2_X1 U1002 ( .A1(G319), .A2(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(G225) );
  XNOR2_X1 U1005 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  NOR2_X1 U1007 ( .A1(G860), .A2(n908), .ZN(n911) );
  XOR2_X1 U1008 ( .A(n909), .B(KEYINPUT73), .Z(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(G145) );
  INV_X1 U1010 ( .A(G120), .ZN(G236) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  INV_X1 U1012 ( .A(G96), .ZN(G221) );
  INV_X1 U1013 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(G325) );
  INV_X1 U1015 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1016 ( .A(G2072), .B(n914), .Z(n916) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n915) );
  NOR2_X1 U1018 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1019 ( .A(KEYINPUT50), .B(n917), .ZN(n935) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n924) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n922) );
  XNOR2_X1 U1023 ( .A(KEYINPUT116), .B(n922), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n933) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1028 ( .A(KEYINPUT51), .B(n929), .Z(n931) );
  XNOR2_X1 U1029 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(n931), .B(n930), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(n938), .ZN(n940) );
  INV_X1 U1035 ( .A(KEYINPUT55), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n941), .A2(G29), .ZN(n1024) );
  XNOR2_X1 U1038 ( .A(G16), .B(KEYINPUT56), .ZN(n967) );
  XOR2_X1 U1039 ( .A(G1966), .B(G168), .Z(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1041 ( .A(KEYINPUT57), .B(n944), .Z(n965) );
  XNOR2_X1 U1042 ( .A(G1348), .B(KEYINPUT122), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n946), .B(n945), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G1961), .B(G301), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n960) );
  XNOR2_X1 U1046 ( .A(G1956), .B(KEYINPUT123), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(n949), .B(G299), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n953) );
  AND2_X1 U1049 ( .A1(G303), .A2(G1971), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(n958), .B(KEYINPUT124), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(G1341), .B(n961), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n996) );
  INV_X1 U1059 ( .A(G16), .ZN(n994) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G21), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(G5), .B(G1961), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n982) );
  XNOR2_X1 U1063 ( .A(n970), .B(G19), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(n971), .B(G20), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n979) );
  XOR2_X1 U1066 ( .A(G1981), .B(G6), .Z(n977) );
  XOR2_X1 U1067 ( .A(KEYINPUT59), .B(G4), .Z(n974) );
  XNOR2_X1 U1068 ( .A(KEYINPUT125), .B(n974), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(n975), .B(G1348), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n980), .B(KEYINPUT60), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n990) );
  XNOR2_X1 U1074 ( .A(G1976), .B(G23), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G22), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1077 ( .A(G1986), .B(KEYINPUT126), .Z(n985) );
  XNOR2_X1 U1078 ( .A(G24), .B(n985), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT58), .B(n988), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1082 ( .A(n991), .B(KEYINPUT61), .Z(n992) );
  XNOR2_X1 U1083 ( .A(KEYINPUT127), .B(n992), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n1022) );
  XOR2_X1 U1086 ( .A(G25), .B(G1991), .Z(n997) );
  NAND2_X1 U1087 ( .A1(n997), .A2(G28), .ZN(n1001) );
  XOR2_X1 U1088 ( .A(G27), .B(n998), .Z(n999) );
  XNOR2_X1 U1089 ( .A(KEYINPUT120), .B(n999), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1009) );
  XNOR2_X1 U1091 ( .A(n1002), .B(G32), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(G2067), .B(G26), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G2072), .B(G33), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT119), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(n1010), .B(KEYINPUT53), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(G2084), .B(G34), .Z(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT54), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G35), .B(G2090), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(KEYINPUT55), .B(n1016), .ZN(n1018) );
  INV_X1 U1105 ( .A(G29), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(G11), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(KEYINPUT121), .B(n1020), .Z(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

