//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G217), .A3(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G128), .B(G143), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT95), .ZN(new_n194));
  INV_X1    g008(.A(G122), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G116), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT95), .A3(G122), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n197), .A2(G122), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT97), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT97), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n199), .A2(new_n205), .A3(new_n200), .A4(new_n202), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT98), .ZN(new_n208));
  INV_X1    g022(.A(new_n199), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT14), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n208), .B(new_n202), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n210), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n210), .B1(new_n196), .B2(new_n198), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT98), .B1(new_n213), .B2(new_n201), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  AOI211_X1 g029(.A(new_n193), .B(new_n207), .C1(new_n215), .C2(G107), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT13), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  OAI22_X1  g032(.A1(KEYINPUT96), .A2(new_n217), .B1(new_n218), .B2(G128), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n217), .A2(KEYINPUT96), .ZN(new_n220));
  OAI21_X1  g034(.A(G134), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g035(.A(new_n221), .B(new_n190), .Z(new_n222));
  OAI21_X1  g036(.A(G107), .B1(new_n209), .B2(new_n201), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n203), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n189), .B1(new_n216), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n207), .B1(new_n215), .B2(G107), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n192), .ZN(new_n229));
  INV_X1    g043(.A(new_n189), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT99), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G902), .ZN(new_n234));
  OAI211_X1 g048(.A(KEYINPUT99), .B(new_n189), .C1(new_n216), .C2(new_n226), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT100), .ZN(new_n237));
  INV_X1    g051(.A(G478), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(KEYINPUT15), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT100), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n233), .A2(new_n240), .A3(new_n234), .A4(new_n235), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  OR2_X1    g056(.A1(new_n236), .A2(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(G237), .A2(G953), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(G143), .A3(G214), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(G143), .B1(new_n245), .B2(G214), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT17), .B(G131), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT93), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(G214), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n218), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n246), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT93), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT17), .A4(G131), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G140), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G125), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT77), .B1(new_n258), .B2(KEYINPUT16), .ZN(new_n259));
  OR3_X1    g073(.A1(new_n258), .A2(KEYINPUT77), .A3(KEYINPUT16), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n257), .A2(KEYINPUT76), .A3(G125), .ZN(new_n261));
  XNOR2_X1  g075(.A(G125), .B(G140), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(KEYINPUT76), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT16), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n259), .B(new_n260), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n261), .ZN(new_n268));
  INV_X1    g082(.A(G125), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G140), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n258), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT76), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT16), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n274), .A2(G146), .A3(new_n259), .A4(new_n260), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n256), .A2(new_n267), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT94), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n253), .B(G131), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n278), .A2(KEYINPUT17), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT94), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n256), .A2(new_n267), .A3(new_n275), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G113), .B(G122), .ZN(new_n283));
  INV_X1    g097(.A(G104), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n262), .A2(new_n266), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n273), .B2(new_n266), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT92), .ZN(new_n288));
  INV_X1    g102(.A(new_n253), .ZN(new_n289));
  AND4_X1   g103(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT18), .A4(G131), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n289), .A2(new_n288), .B1(KEYINPUT18), .B2(G131), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n282), .A2(new_n285), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n263), .A2(KEYINPUT19), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n294), .B1(KEYINPUT19), .B2(new_n271), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n275), .B(new_n278), .C1(new_n295), .C2(G146), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n285), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G475), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n234), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT20), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n293), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n285), .B1(new_n282), .B2(new_n292), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n234), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G475), .ZN(new_n308));
  AOI21_X1  g122(.A(G475), .B1(new_n293), .B2(new_n299), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT20), .A3(new_n234), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n304), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n244), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G952), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(G953), .ZN(new_n314));
  NAND2_X1  g128(.A1(G234), .A2(G237), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT21), .B(G898), .Z(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(G902), .A3(G953), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n317), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G210), .B1(G237), .B2(G902), .ZN(new_n323));
  XOR2_X1   g137(.A(new_n323), .B(KEYINPUT91), .Z(new_n324));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n200), .A4(G104), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n284), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n328));
  OAI22_X1  g142(.A1(new_n284), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G101), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n331), .A2(KEYINPUT4), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT2), .A2(G113), .ZN(new_n333));
  NAND2_X1  g147(.A1(KEYINPUT2), .A2(G113), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n333), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G119), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G116), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n197), .A2(G119), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n338), .B(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n332), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n330), .A2(new_n346), .A3(G101), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT4), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n330), .B2(G101), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n350));
  INV_X1    g164(.A(G101), .ZN(new_n351));
  AND4_X1   g165(.A1(new_n351), .A2(new_n327), .A3(new_n328), .A4(new_n329), .ZN(new_n352));
  NOR4_X1   g166(.A1(new_n348), .A2(new_n349), .A3(new_n350), .A4(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n347), .A2(KEYINPUT4), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(KEYINPUT80), .B2(new_n331), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT81), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n345), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT87), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT5), .ZN(new_n359));
  OR3_X1    g173(.A1(new_n197), .A2(KEYINPUT5), .A3(G119), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G113), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT86), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n338), .A2(new_n342), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT86), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n359), .A2(new_n360), .A3(new_n364), .A4(G113), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n327), .A2(new_n328), .A3(new_n329), .A4(new_n351), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n200), .A2(G104), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n284), .A2(G107), .ZN(new_n369));
  OAI21_X1  g183(.A(G101), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n358), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n361), .A2(KEYINPUT86), .B1(new_n338), .B2(new_n342), .ZN(new_n373));
  INV_X1    g187(.A(new_n371), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT87), .A4(new_n365), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(G110), .B(G122), .Z(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n357), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n371), .A3(new_n365), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n377), .B(KEYINPUT8), .Z(new_n381));
  NAND2_X1  g195(.A1(new_n363), .A2(new_n361), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n382), .B(KEYINPUT88), .Z(new_n383));
  OAI211_X1 g197(.A(new_n380), .B(new_n381), .C1(new_n383), .C2(new_n371), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n188), .A2(G224), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT7), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT65), .B1(new_n218), .B2(G146), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT65), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n266), .A3(G143), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT1), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n218), .A2(G146), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n392), .A2(new_n393), .A3(G128), .A4(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n218), .A2(G146), .ZN(new_n396));
  OAI21_X1  g210(.A(G128), .B1(new_n396), .B2(new_n393), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n266), .A2(G143), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n269), .ZN(new_n402));
  OR2_X1    g216(.A1(KEYINPUT0), .A2(G128), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT0), .A2(G128), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n266), .A2(G143), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n403), .B(new_n404), .C1(new_n405), .C2(new_n396), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT64), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n392), .A2(KEYINPUT0), .A3(G128), .A4(new_n394), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n399), .A2(KEYINPUT64), .A3(new_n403), .A4(new_n404), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n408), .A2(new_n409), .A3(G125), .A4(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n388), .B1(new_n402), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT89), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n402), .A2(new_n388), .A3(new_n411), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n379), .A2(new_n384), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT90), .A3(new_n234), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n331), .A2(KEYINPUT80), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(KEYINPUT4), .A3(new_n347), .A4(new_n367), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n350), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT81), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n344), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n372), .A2(new_n375), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n377), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n379), .A3(KEYINPUT6), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n402), .A2(new_n411), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n426), .B(new_n385), .Z(new_n427));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n428), .B(new_n377), .C1(new_n422), .C2(new_n423), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n417), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT90), .B1(new_n416), .B2(new_n234), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n324), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n416), .A2(new_n234), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(new_n323), .A3(new_n430), .A4(new_n417), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n322), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G214), .B1(G237), .B2(G902), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT85), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n312), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n332), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n353), .B2(new_n356), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT11), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n191), .B2(G137), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT66), .B(new_n446), .C1(new_n191), .C2(G137), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G137), .ZN(new_n453));
  INV_X1    g267(.A(G137), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(KEYINPUT67), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT11), .B(G134), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G131), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n454), .A2(G134), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n451), .A2(new_n456), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n454), .A2(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n452), .A2(G137), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n446), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n458), .B1(new_n464), .B2(G134), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n457), .B1(new_n465), .B2(new_n451), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n374), .A2(new_n401), .A3(KEYINPUT10), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n392), .A2(new_n394), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n397), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n371), .B1(new_n470), .B2(new_n395), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n472));
  OAI21_X1  g286(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n445), .A2(new_n467), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT83), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n445), .A2(new_n477), .A3(new_n467), .A4(new_n474), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n467), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n443), .B1(new_n420), .B2(new_n421), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n480), .B1(new_n481), .B2(new_n473), .ZN(new_n482));
  XNOR2_X1  g296(.A(G110), .B(G140), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n188), .A2(G227), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n483), .B(new_n484), .Z(new_n485));
  NAND3_X1  g299(.A1(new_n479), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n471), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n401), .B2(new_n374), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n488), .A2(KEYINPUT12), .A3(new_n480), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT12), .B1(new_n488), .B2(new_n480), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n476), .B2(new_n478), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n486), .B(G469), .C1(new_n492), .C2(new_n485), .ZN(new_n493));
  NAND2_X1  g307(.A1(G469), .A2(G902), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n420), .A2(new_n421), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n473), .B1(new_n496), .B2(new_n444), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n477), .B1(new_n497), .B2(new_n467), .ZN(new_n498));
  NOR4_X1   g312(.A1(new_n481), .A2(KEYINPUT83), .A3(new_n480), .A4(new_n473), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n485), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT84), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n491), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n479), .A2(KEYINPUT84), .A3(new_n485), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n485), .B1(new_n479), .B2(new_n482), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G469), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n495), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n187), .ZN(new_n511));
  OAI21_X1  g325(.A(G221), .B1(new_n511), .B2(G902), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n441), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(G101), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n245), .A2(G210), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT74), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n456), .A2(new_n459), .ZN(new_n521));
  INV_X1    g335(.A(new_n450), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n454), .A2(G134), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT66), .B1(new_n523), .B2(new_n446), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G131), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n520), .B1(new_n526), .B2(new_n460), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n462), .A2(new_n463), .A3(new_n191), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n523), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G131), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n401), .A2(new_n460), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n519), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n442), .B1(new_n461), .B2(new_n466), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n401), .A2(new_n460), .A3(new_n530), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(KEYINPUT74), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n343), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT28), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n527), .A2(new_n531), .A3(new_n343), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n536), .B1(new_n533), .B2(new_n534), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n518), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT70), .ZN(new_n546));
  INV_X1    g360(.A(new_n518), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n546), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n533), .A2(new_n536), .A3(new_n534), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(KEYINPUT70), .A3(new_n518), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(KEYINPUT68), .A2(KEYINPUT30), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT68), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n552), .B(new_n555), .C1(new_n527), .C2(new_n531), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n533), .A2(new_n553), .A3(new_n554), .A4(new_n534), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n343), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n545), .B1(new_n551), .B2(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n561));
  NAND3_X1  g375(.A1(new_n551), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT72), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n548), .A2(new_n550), .B1(new_n558), .B2(new_n343), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(KEYINPUT72), .A3(new_n561), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n544), .B(new_n560), .C1(new_n564), .C2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(G472), .A2(G902), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT75), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n544), .ZN(new_n571));
  INV_X1    g385(.A(new_n560), .ZN(new_n572));
  AND4_X1   g386(.A1(KEYINPUT72), .A2(new_n551), .A3(new_n559), .A4(new_n561), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT72), .B1(new_n565), .B2(new_n561), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n568), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT32), .B1(new_n575), .B2(new_n568), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n570), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT75), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT32), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n579), .B(new_n580), .C1(new_n575), .C2(new_n568), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n539), .A2(new_n518), .A3(new_n543), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n559), .A2(new_n549), .ZN(new_n584));
  AOI211_X1 g398(.A(KEYINPUT29), .B(new_n583), .C1(new_n547), .C2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT28), .B1(new_n541), .B2(new_n542), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n539), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n518), .A2(KEYINPUT29), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n234), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G472), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n578), .A2(new_n582), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n267), .A2(new_n275), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT23), .ZN(new_n593));
  INV_X1    g407(.A(G128), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(G119), .B2(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n339), .A2(KEYINPUT23), .A3(G128), .ZN(new_n596));
  OAI22_X1  g410(.A1(new_n595), .A2(new_n596), .B1(G119), .B2(new_n594), .ZN(new_n597));
  XNOR2_X1  g411(.A(G119), .B(G128), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT24), .B(G110), .Z(new_n599));
  AOI22_X1  g413(.A1(new_n597), .A2(G110), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n592), .A2(new_n600), .ZN(new_n601));
  OAI22_X1  g415(.A1(new_n597), .A2(G110), .B1(new_n598), .B2(new_n599), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n275), .A2(new_n286), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT22), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G137), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n604), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n234), .ZN(new_n609));
  AND2_X1   g423(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n610));
  NOR2_X1   g424(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n611));
  OR3_X1    g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G234), .ZN(new_n613));
  OAI21_X1  g427(.A(G217), .B1(new_n613), .B2(G902), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n609), .B2(new_n610), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(G902), .B1(new_n613), .B2(G217), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n608), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n514), .A2(new_n591), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT101), .B(G101), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G3));
  INV_X1    g437(.A(new_n439), .ZN(new_n624));
  INV_X1    g438(.A(new_n323), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n431), .B2(new_n432), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n624), .B1(new_n626), .B2(new_n437), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n237), .A2(new_n238), .A3(new_n241), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT102), .B(KEYINPUT33), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n233), .A2(new_n235), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n227), .A2(new_n231), .A3(KEYINPUT33), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(G478), .A3(new_n234), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n311), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n628), .A2(new_n636), .A3(new_n322), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n575), .A2(new_n568), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n560), .B1(new_n564), .B2(new_n566), .ZN(new_n639));
  AOI21_X1  g453(.A(G902), .B1(new_n639), .B2(new_n571), .ZN(new_n640));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n510), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n619), .A2(new_n513), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n637), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  AND3_X1   g461(.A1(new_n304), .A2(new_n308), .A3(new_n310), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n244), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n628), .A2(new_n322), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n643), .A3(new_n644), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  INV_X1    g467(.A(new_n607), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n604), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n617), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n616), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n642), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n514), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n660), .B(KEYINPUT37), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G110), .ZN(G12));
  NOR3_X1   g476(.A1(new_n510), .A2(new_n513), .A3(new_n658), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n320), .A2(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n316), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n648), .A2(new_n244), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(KEYINPUT103), .A3(new_n627), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(new_n628), .B2(new_n666), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n591), .A2(new_n663), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  NAND2_X1  g486(.A1(new_n505), .A2(new_n507), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n509), .A3(new_n234), .ZN(new_n674));
  INV_X1    g488(.A(new_n495), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n513), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n665), .B(KEYINPUT105), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT39), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT38), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n433), .A2(new_n437), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT104), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n682), .A2(KEYINPUT104), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n681), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n682), .A2(KEYINPUT104), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(KEYINPUT38), .A3(new_n683), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n565), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n547), .B1(new_n541), .B2(new_n542), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n641), .B1(new_n692), .B2(new_n234), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n578), .A2(new_n582), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n680), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n244), .A2(new_n311), .A3(new_n439), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n658), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n218), .ZN(G45));
  NAND3_X1  g515(.A1(new_n635), .A2(new_n311), .A3(new_n665), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n591), .A2(new_n663), .A3(new_n627), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  NAND2_X1  g519(.A1(KEYINPUT106), .A2(G469), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n508), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n706), .ZN(new_n708));
  AOI211_X1 g522(.A(G902), .B(new_n708), .C1(new_n505), .C2(new_n507), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n707), .A2(new_n709), .A3(new_n513), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n591), .A2(new_n620), .A3(new_n637), .A4(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT41), .B(G113), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT107), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n711), .B(new_n713), .ZN(G15));
  NAND4_X1  g528(.A1(new_n591), .A2(new_n620), .A3(new_n650), .A4(new_n710), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  AOI21_X1  g530(.A(KEYINPUT84), .B1(new_n479), .B2(new_n485), .ZN(new_n717));
  INV_X1    g531(.A(new_n485), .ZN(new_n718));
  AOI211_X1 g532(.A(new_n501), .B(new_n718), .C1(new_n476), .C2(new_n478), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n506), .B1(new_n720), .B2(new_n503), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n708), .B1(new_n721), .B2(G902), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n508), .A2(new_n706), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n512), .A2(new_n722), .A3(new_n627), .A4(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n658), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n648), .A2(new_n243), .A3(new_n242), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n322), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n724), .A2(new_n591), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NAND2_X1  g543(.A1(new_n575), .A2(new_n234), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT108), .B1(new_n730), .B2(G472), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n732), .B(new_n641), .C1(new_n575), .C2(new_n234), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n587), .A2(new_n547), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n569), .B1(new_n639), .B2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n731), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n322), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n626), .A2(new_n437), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n698), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n736), .A2(new_n710), .A3(new_n739), .A4(new_n620), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT109), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  XNOR2_X1  g556(.A(new_n702), .B(KEYINPUT110), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n724), .A2(new_n725), .A3(new_n736), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  NAND2_X1  g559(.A1(new_n638), .A2(new_n580), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n568), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n581), .B1(new_n748), .B2(new_n570), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n619), .B1(new_n749), .B2(new_n590), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n433), .A2(new_n439), .A3(new_n437), .ZN(new_n751));
  AOI211_X1 g565(.A(G469), .B(G902), .C1(new_n505), .C2(new_n507), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n512), .B(new_n751), .C1(new_n752), .C2(new_n495), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT111), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n676), .A2(new_n755), .A3(new_n751), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n750), .A2(new_n757), .A3(new_n743), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  INV_X1    g573(.A(new_n743), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n754), .B2(new_n756), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n746), .A2(new_n747), .A3(new_n590), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n762), .A2(new_n620), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n759), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n758), .A2(new_n759), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n457), .ZN(G33));
  NAND2_X1  g581(.A1(new_n591), .A2(new_n620), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n756), .B2(new_n754), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n667), .A2(KEYINPUT112), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n667), .A2(KEYINPUT112), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(new_n770), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n750), .A2(new_n757), .A3(new_n771), .A4(new_n772), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT113), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n479), .A2(new_n482), .A3(new_n485), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n485), .B1(new_n479), .B2(new_n503), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n486), .B(KEYINPUT45), .C1(new_n492), .C2(new_n485), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n782), .A3(G469), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(new_n494), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(KEYINPUT46), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n494), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n674), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(KEYINPUT114), .A3(new_n674), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n785), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n513), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n648), .A2(new_n635), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT43), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(new_n642), .A3(new_n725), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT44), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n792), .A2(new_n678), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n751), .B1(new_n797), .B2(KEYINPUT44), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n454), .ZN(G39));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n791), .B2(new_n513), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n785), .A2(new_n789), .A3(new_n790), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(KEYINPUT47), .A3(new_n512), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n591), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n751), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n808), .A2(new_n620), .A3(new_n702), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  NAND2_X1  g625(.A1(new_n313), .A2(new_n188), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n813));
  INV_X1    g627(.A(new_n806), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT47), .B1(new_n805), .B2(new_n512), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n804), .A2(KEYINPUT117), .A3(new_n806), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n722), .A2(new_n723), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n512), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n620), .A2(new_n795), .A3(new_n736), .A4(new_n317), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n823), .A2(new_n751), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n822), .B1(new_n821), .B2(new_n824), .ZN(new_n826));
  INV_X1    g640(.A(new_n695), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n818), .A2(new_n513), .A3(new_n808), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n620), .A3(new_n317), .A4(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n829), .A2(new_n311), .A3(new_n635), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n818), .A2(new_n513), .A3(new_n439), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n689), .B1(new_n831), .B2(KEYINPUT119), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n831), .A2(KEYINPUT119), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n823), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT50), .A4(new_n823), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n830), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n828), .A2(new_n317), .A3(new_n795), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n736), .A2(new_n725), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n825), .A2(new_n826), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT120), .B1(new_n845), .B2(KEYINPUT51), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n821), .A2(new_n824), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT118), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n847), .B(new_n848), .C1(new_n852), .C2(new_n844), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n829), .A2(new_n636), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n804), .A2(new_n806), .A3(new_n820), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n848), .B1(new_n856), .B2(new_n824), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n838), .A2(new_n857), .A3(new_n843), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n840), .A2(new_n763), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT48), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n823), .A2(new_n724), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n314), .A2(new_n858), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n744), .A2(new_n671), .A3(new_n704), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n725), .B1(new_n749), .B2(new_n694), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n698), .A2(new_n738), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n865), .A2(new_n676), .A3(new_n665), .A4(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT52), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n744), .A2(new_n671), .A3(new_n704), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n695), .A2(new_n676), .A3(new_n658), .A4(new_n665), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n866), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n776), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n758), .A2(new_n759), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n761), .A2(new_n765), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n728), .A2(new_n711), .A3(new_n715), .A4(new_n740), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n438), .A2(new_n440), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n649), .A2(new_n636), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n643), .A2(new_n644), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n621), .A2(new_n660), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n665), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT115), .B1(new_n726), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n312), .A2(new_n887), .A3(new_n665), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n751), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT116), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n886), .A2(new_n891), .A3(new_n888), .A4(new_n751), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n890), .A2(new_n591), .A3(new_n663), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n761), .A2(new_n842), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n878), .A2(new_n884), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n863), .B1(new_n875), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n728), .A2(new_n715), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n621), .A2(new_n660), .A3(new_n882), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n711), .A2(new_n740), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n893), .A4(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n894), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n900), .A2(new_n766), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n744), .A2(new_n671), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(KEYINPUT52), .A3(new_n704), .A4(new_n868), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n873), .B1(new_n870), .B2(new_n872), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n904), .A2(new_n905), .B1(new_n773), .B2(new_n775), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n906), .A3(KEYINPUT53), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n896), .A2(KEYINPUT54), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT54), .B1(new_n896), .B2(new_n907), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n855), .B(new_n862), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n812), .B1(new_n854), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n818), .B(KEYINPUT49), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n644), .A2(new_n648), .A3(new_n440), .A4(new_n635), .ZN(new_n914));
  OR4_X1    g728(.A1(new_n689), .A2(new_n913), .A3(new_n695), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n912), .A2(new_n915), .ZN(G75));
  NAND2_X1  g730(.A1(new_n425), .A2(new_n429), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n427), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT55), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n234), .B1(new_n896), .B2(new_n907), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(G210), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n188), .A2(G952), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n922), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n920), .B2(new_n324), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(G51));
  NAND2_X1  g741(.A1(new_n896), .A2(new_n907), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT54), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n494), .B(KEYINPUT57), .Z(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n908), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n721), .B(KEYINPUT121), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n783), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n920), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n924), .B1(new_n934), .B2(new_n936), .ZN(G54));
  NAND3_X1  g751(.A1(new_n920), .A2(KEYINPUT58), .A3(G475), .ZN(new_n938));
  INV_X1    g752(.A(new_n300), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(new_n924), .ZN(G60));
  XNOR2_X1  g756(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n238), .A2(new_n234), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n930), .A2(new_n908), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n632), .A2(new_n633), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n924), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT60), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n875), .A2(new_n895), .A3(new_n863), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT53), .B1(new_n902), .B2(new_n906), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n656), .B(new_n953), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n924), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n952), .B1(new_n896), .B2(new_n907), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n956), .B(new_n957), .C1(new_n608), .C2(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n959), .A2(KEYINPUT123), .A3(KEYINPUT61), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT61), .B1(new_n959), .B2(KEYINPUT123), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(G66));
  INV_X1    g776(.A(new_n884), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n188), .B1(new_n318), .B2(G224), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n963), .A2(new_n188), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n964), .B2(new_n965), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n917), .B1(G898), .B2(new_n188), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G69));
  NAND2_X1  g783(.A1(G900), .A2(G953), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n801), .B1(new_n807), .B2(new_n809), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n792), .A2(new_n678), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n972), .A2(new_n973), .A3(new_n867), .A4(new_n763), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n792), .A2(new_n678), .A3(new_n867), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT126), .B1(new_n975), .B2(new_n764), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n766), .A2(new_n870), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n971), .A2(new_n977), .A3(new_n776), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n970), .B1(new_n979), .B2(G953), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n295), .B(KEYINPUT125), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n558), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(G227), .A2(G900), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(G953), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n700), .A2(new_n870), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT62), .ZN(new_n987));
  INV_X1    g801(.A(new_n753), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n750), .A2(new_n678), .A3(new_n988), .A4(new_n881), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n971), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n188), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n983), .B(new_n985), .C1(new_n982), .C2(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n980), .A2(G953), .A3(new_n984), .A4(new_n982), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  OAI211_X1 g810(.A(KEYINPUT127), .B(new_n996), .C1(new_n979), .C2(new_n963), .ZN(new_n997));
  INV_X1    g811(.A(new_n584), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n810), .ZN(new_n1000));
  INV_X1    g814(.A(new_n776), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n1000), .A2(new_n1001), .A3(new_n801), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1002), .A2(new_n884), .A3(new_n978), .A4(new_n977), .ZN(new_n1003));
  AOI21_X1  g817(.A(KEYINPUT127), .B1(new_n1003), .B2(new_n996), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n999), .A2(new_n1004), .A3(new_n518), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n996), .B1(new_n990), .B2(new_n963), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n518), .A3(new_n584), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n690), .B1(new_n998), .B2(new_n518), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n928), .A2(new_n996), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1007), .A2(new_n957), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1005), .A2(new_n1010), .ZN(G57));
endmodule


