//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  AND2_X1   g001(.A1(KEYINPUT69), .A2(G237), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT69), .A2(G237), .ZN(new_n189));
  OAI211_X1 g003(.A(G214), .B(new_n187), .C1(new_n188), .C2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT69), .B(G237), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n193), .A2(G143), .A3(G214), .A4(new_n187), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G131), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT85), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n198), .A2(KEYINPUT85), .A3(new_n199), .A4(new_n200), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(G125), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n207), .B1(new_n211), .B2(new_n205), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI211_X1 g028(.A(G146), .B(new_n207), .C1(new_n211), .C2(new_n205), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n196), .B1(new_n192), .B2(new_n194), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n216), .B1(KEYINPUT17), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n203), .A2(new_n204), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n220));
  INV_X1    g034(.A(G131), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT82), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n192), .A2(new_n194), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n211), .B(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n223), .B1(new_n192), .B2(new_n194), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT83), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n195), .A2(new_n222), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT83), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n229), .A2(new_n230), .A3(new_n225), .A4(new_n224), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n219), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G113), .B(G122), .ZN(new_n234));
  INV_X1    g048(.A(G104), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n219), .A2(new_n236), .A3(new_n232), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G475), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT19), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT19), .B1(new_n208), .B2(new_n210), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n213), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n215), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(new_n198), .B2(new_n200), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n232), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT84), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(new_n237), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n248), .B1(new_n228), .B2(new_n231), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT84), .B1(new_n253), .B2(new_n236), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n252), .A2(new_n239), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT86), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT20), .ZN(new_n258));
  NOR2_X1   g072(.A1(G475), .A2(G902), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n257), .A2(new_n258), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n255), .A2(KEYINPUT86), .A3(new_n258), .A4(new_n259), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n243), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT87), .B1(new_n191), .B2(G128), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT87), .ZN(new_n266));
  INV_X1    g080(.A(G128), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT88), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n191), .A2(G128), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n269), .B2(new_n271), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n264), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n271), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT88), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(G134), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT89), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n274), .A2(new_n278), .A3(KEYINPUT89), .ZN(new_n282));
  INV_X1    g096(.A(G116), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G122), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT14), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT14), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n283), .A3(G122), .ZN(new_n287));
  INV_X1    g101(.A(G122), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G116), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT90), .A4(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT91), .ZN(new_n291));
  INV_X1    g105(.A(G107), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n288), .A2(KEYINPUT14), .A3(G116), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT90), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n290), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n290), .A2(new_n295), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n289), .A2(new_n284), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n297), .A2(KEYINPUT91), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n281), .A2(new_n282), .A3(new_n296), .A4(new_n299), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n271), .B(KEYINPUT13), .Z(new_n301));
  INV_X1    g115(.A(new_n269), .ZN(new_n302));
  OAI21_X1  g116(.A(G134), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n298), .B(new_n292), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n274), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT73), .B(G217), .Z(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT9), .B(G234), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n307), .A2(G953), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n305), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n299), .A2(new_n296), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(new_n279), .B2(new_n280), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n312), .B1(new_n314), .B2(new_n282), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n309), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT72), .B(G902), .ZN(new_n318));
  INV_X1    g132(.A(G478), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT15), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n317), .A2(KEYINPUT92), .A3(new_n318), .A4(new_n321), .ZN(new_n322));
  AOI211_X1 g136(.A(new_n312), .B(new_n310), .C1(new_n314), .C2(new_n282), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n309), .B1(new_n300), .B2(new_n305), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT92), .B(new_n318), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n320), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n187), .A2(G952), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n327), .B1(G234), .B2(G237), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT21), .B(G898), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n329), .B(KEYINPUT93), .Z(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI211_X1 g145(.A(new_n187), .B(new_n318), .C1(G234), .C2(G237), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n322), .A2(new_n326), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT94), .B1(new_n263), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n257), .A2(new_n258), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n255), .A2(new_n259), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n261), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n322), .A2(new_n326), .A3(new_n334), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT94), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .A4(new_n243), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT67), .ZN(new_n345));
  INV_X1    g159(.A(G137), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G134), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(G134), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT65), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT11), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n345), .A2(new_n347), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n264), .A2(G137), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT11), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(KEYINPUT65), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n349), .A2(KEYINPUT11), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT67), .B1(new_n346), .B2(G134), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n351), .A2(new_n356), .A3(new_n196), .A4(new_n357), .ZN(new_n358));
  OAI22_X1  g172(.A1(KEYINPUT65), .A2(new_n353), .B1(new_n264), .B2(G137), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n345), .A2(new_n264), .A3(G137), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n353), .A2(KEYINPUT65), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n348), .B1(new_n350), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G131), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT64), .B1(new_n191), .B2(G146), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT64), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n213), .A3(G143), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n191), .A2(G146), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n191), .A2(G146), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT1), .ZN(new_n372));
  OAI21_X1  g186(.A(G128), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n267), .A2(KEYINPUT1), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n366), .A2(new_n368), .A3(new_n369), .A4(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n292), .A3(G104), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n235), .A2(G107), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT77), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n235), .A2(G107), .ZN(new_n382));
  OAI211_X1 g196(.A(G101), .B(new_n379), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n292), .A2(KEYINPUT76), .A3(G104), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT3), .ZN(new_n385));
  INV_X1    g199(.A(G101), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n387), .A2(new_n292), .A3(KEYINPUT76), .A4(G104), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n385), .A2(new_n386), .A3(new_n388), .A4(new_n380), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n377), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n383), .A2(new_n389), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n213), .A2(G143), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n369), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n373), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n376), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n365), .B1(new_n391), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT12), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(KEYINPUT12), .B(new_n365), .C1(new_n391), .C2(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(KEYINPUT0), .A2(G128), .ZN(new_n403));
  OR2_X1    g217(.A1(KEYINPUT0), .A2(G128), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n213), .A2(G143), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n403), .B(new_n404), .C1(new_n371), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n403), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n366), .A2(new_n368), .A3(new_n407), .A4(new_n369), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n384), .A2(KEYINPUT3), .B1(new_n235), .B2(G107), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n386), .B1(new_n410), .B2(new_n388), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n385), .A2(new_n388), .A3(new_n380), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G101), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT4), .A3(new_n389), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT10), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(new_n395), .B2(new_n376), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n413), .A2(new_n416), .B1(new_n392), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n365), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n374), .A2(new_n376), .ZN(new_n421));
  AOI211_X1 g235(.A(KEYINPUT78), .B(KEYINPUT10), .C1(new_n392), .C2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT78), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n389), .A3(new_n383), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n424), .B2(new_n417), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n419), .B(new_n420), .C1(new_n422), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n402), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G110), .B(G140), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n187), .A2(G227), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n409), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n414), .A2(new_n412), .A3(G101), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n389), .A2(KEYINPUT4), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n431), .B(new_n432), .C1(new_n433), .C2(new_n411), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n392), .A2(new_n418), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n417), .B1(new_n377), .B2(new_n390), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT78), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n424), .A2(new_n423), .A3(new_n417), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n430), .B1(new_n440), .B2(new_n420), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n419), .B1(new_n422), .B2(new_n425), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n365), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n427), .A2(new_n430), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G469), .ZN(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  INV_X1    g260(.A(new_n430), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n402), .A2(new_n426), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n447), .B1(new_n443), .B2(new_n426), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n446), .B(new_n318), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n446), .A2(new_n241), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n445), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G214), .B1(G237), .B2(G902), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT2), .B(G113), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G119), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G116), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n283), .A2(G119), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT5), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n462), .B(G113), .C1(KEYINPUT5), .C2(new_n458), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n392), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(new_n459), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n455), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n467), .B(new_n432), .C1(new_n433), .C2(new_n411), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G122), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n464), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(KEYINPUT8), .ZN(new_n471));
  AND4_X1   g285(.A1(new_n461), .A2(new_n463), .A3(new_n389), .A4(new_n383), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n461), .A2(new_n463), .B1(new_n383), .B2(new_n389), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT80), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n395), .A2(new_n475), .A3(new_n209), .A4(new_n376), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n187), .A2(G224), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n478), .A2(KEYINPUT81), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(KEYINPUT81), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n395), .A2(new_n209), .A3(new_n376), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT80), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n209), .B1(new_n406), .B2(new_n408), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n476), .B(new_n481), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n470), .A2(new_n474), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n482), .B1(new_n484), .B2(KEYINPUT79), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n484), .A2(KEYINPUT79), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n488), .A2(KEYINPUT7), .A3(new_n477), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(G902), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n464), .A2(new_n468), .ZN(new_n492));
  INV_X1    g306(.A(new_n469), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT6), .A3(new_n470), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n488), .A2(new_n477), .A3(new_n489), .ZN(new_n496));
  INV_X1    g310(.A(new_n489), .ZN(new_n497));
  OAI211_X1 g311(.A(G224), .B(new_n187), .C1(new_n497), .C2(new_n487), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT6), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n492), .A2(new_n500), .A3(new_n493), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n491), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G210), .B1(G237), .B2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n491), .A2(new_n502), .A3(new_n504), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(G221), .B1(new_n308), .B2(G902), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n453), .A2(new_n454), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n344), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT95), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n307), .B1(G234), .B2(new_n318), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT25), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT74), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G137), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT23), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n457), .B2(G128), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n267), .A2(KEYINPUT23), .A3(G119), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(new_n523), .C1(G119), .C2(new_n267), .ZN(new_n524));
  XNOR2_X1  g338(.A(G119), .B(G128), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT24), .B(G110), .Z(new_n526));
  AOI22_X1  g340(.A1(new_n524), .A2(G110), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n216), .A2(new_n527), .ZN(new_n528));
  OAI22_X1  g342(.A1(new_n524), .A2(G110), .B1(new_n525), .B2(new_n526), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n529), .B(new_n215), .C1(G146), .C2(new_n211), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n528), .A2(KEYINPUT75), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT75), .B1(new_n528), .B2(new_n530), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n520), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n532), .A2(new_n520), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n318), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n516), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT25), .A4(new_n318), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n515), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n535), .A2(G902), .A3(new_n514), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT70), .ZN(new_n543));
  INV_X1    g357(.A(new_n189), .ZN(new_n544));
  NAND2_X1  g358(.A1(KEYINPUT69), .A2(G237), .ZN(new_n545));
  AOI21_X1  g359(.A(G953), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G210), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT27), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT27), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n549), .A3(G210), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT26), .B(G101), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n548), .B2(new_n550), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n543), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(KEYINPUT70), .A3(new_n552), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n359), .A2(new_n357), .A3(new_n360), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n221), .B1(new_n559), .B2(new_n356), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n361), .A2(new_n197), .A3(new_n363), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n431), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n467), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n348), .A2(KEYINPUT68), .ZN(new_n564));
  INV_X1    g378(.A(new_n347), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n348), .A2(KEYINPUT68), .ZN(new_n567));
  OAI21_X1  g381(.A(G131), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n396), .A2(new_n358), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n562), .A2(KEYINPUT28), .A3(new_n563), .A4(new_n569), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n396), .A2(new_n358), .A3(new_n568), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n409), .B1(new_n358), .B2(new_n364), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n467), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n562), .A2(new_n563), .A3(new_n569), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT28), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n558), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT30), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT30), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n562), .B2(new_n569), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n467), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n553), .A2(new_n554), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n575), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT31), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n575), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT30), .B1(new_n571), .B2(new_n572), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n562), .A2(new_n580), .A3(new_n569), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n587), .B1(new_n590), .B2(new_n467), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(KEYINPUT31), .A3(new_n583), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n578), .B1(new_n586), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(G472), .A2(G902), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT32), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n578), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT31), .B1(new_n591), .B2(new_n583), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n563), .B1(new_n588), .B2(new_n589), .ZN(new_n599));
  INV_X1    g413(.A(new_n583), .ZN(new_n600));
  NOR4_X1   g414(.A1(new_n599), .A2(new_n600), .A3(new_n587), .A4(new_n585), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n597), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT32), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n603), .A3(new_n594), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n596), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n574), .A2(new_n577), .A3(new_n558), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT29), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n591), .A2(new_n583), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n318), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT71), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n573), .A2(new_n575), .A3(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(KEYINPUT71), .B(new_n467), .C1(new_n571), .C2(new_n572), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n577), .B1(new_n614), .B2(new_n576), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n615), .A2(new_n607), .A3(new_n600), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n610), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n542), .B1(new_n605), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n344), .A2(new_n619), .A3(new_n511), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n513), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  NAND2_X1  g436(.A1(new_n602), .A2(new_n318), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n623), .A2(G472), .B1(new_n594), .B2(new_n602), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n453), .A2(new_n509), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n625), .A2(new_n542), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n324), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT98), .B1(new_n315), .B2(new_n309), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n629), .A2(new_n630), .A3(KEYINPUT33), .A4(new_n316), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n632));
  NAND2_X1  g446(.A1(new_n317), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n536), .A2(new_n319), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n317), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n319), .B1(new_n636), .B2(new_n536), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n263), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n491), .A2(new_n502), .A3(new_n504), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n504), .B1(new_n491), .B2(new_n502), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n454), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT96), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n508), .A2(KEYINPUT96), .A3(new_n454), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n333), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n627), .A2(new_n640), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT34), .B(G104), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  NOR2_X1   g465(.A1(new_n338), .A2(KEYINPUT20), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n258), .B1(new_n255), .B2(new_n259), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n243), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n322), .A2(new_n326), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n647), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n647), .A2(new_n656), .A3(KEYINPUT100), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n627), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT35), .B(G107), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT101), .B(KEYINPUT102), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NOR2_X1   g480(.A1(new_n520), .A2(KEYINPUT36), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n528), .A2(new_n530), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n669), .A2(new_n241), .A3(new_n515), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n539), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n625), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n513), .A2(new_n620), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NOR3_X1   g489(.A1(new_n593), .A2(KEYINPUT32), .A3(new_n595), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n603), .B1(new_n602), .B2(new_n594), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n617), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n645), .A2(new_n646), .ZN(new_n679));
  INV_X1    g493(.A(new_n509), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n440), .A2(new_n420), .ZN(new_n681));
  INV_X1    g495(.A(new_n426), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n430), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n441), .A2(new_n402), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n536), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n451), .B1(new_n685), .B2(new_n446), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n680), .B1(new_n686), .B2(new_n445), .ZN(new_n687));
  INV_X1    g501(.A(new_n671), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n678), .A2(new_n679), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n328), .B(KEYINPUT104), .Z(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT103), .B(G900), .Z(new_n692));
  AND2_X1   g506(.A1(new_n332), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n656), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT105), .B1(new_n689), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n626), .B1(new_n645), .B2(new_n646), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n654), .A2(new_n655), .A3(new_n694), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n671), .B1(new_n605), .B2(new_n617), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n698), .A2(new_n699), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  XOR2_X1   g518(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n508), .B(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n454), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n706), .A2(new_n707), .A3(new_n688), .ZN(new_n708));
  INV_X1    g522(.A(new_n584), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n614), .A2(new_n558), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n241), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G472), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n605), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n263), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n655), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n708), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n717), .A2(KEYINPUT107), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n694), .B(KEYINPUT39), .Z(new_n719));
  NAND2_X1  g533(.A1(new_n687), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n720), .B(KEYINPUT40), .Z(new_n721));
  NAND2_X1  g535(.A1(new_n717), .A2(KEYINPUT107), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n718), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G143), .ZN(G45));
  AND3_X1   g538(.A1(new_n263), .A2(new_n638), .A3(new_n695), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n689), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n213), .ZN(G48));
  NAND2_X1  g542(.A1(new_n443), .A2(new_n426), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n729), .A2(new_n430), .B1(new_n441), .B2(new_n402), .ZN(new_n730));
  OAI21_X1  g544(.A(G469), .B1(new_n730), .B2(new_n536), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n509), .A3(new_n450), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n640), .A2(new_n618), .A3(new_n647), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT109), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n736), .B(KEYINPUT108), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n734), .B(new_n737), .ZN(G15));
  NAND2_X1  g552(.A1(new_n618), .A2(new_n733), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n659), .B2(new_n660), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n283), .ZN(G18));
  INV_X1    g555(.A(new_n344), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n732), .B1(new_n645), .B2(new_n646), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n701), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n457), .ZN(G21));
  NAND2_X1  g560(.A1(new_n322), .A2(new_n326), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n679), .A2(new_n263), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n732), .A2(new_n333), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n586), .A2(new_n592), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n615), .A2(new_n557), .A3(new_n555), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n595), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(G472), .B1(new_n593), .B2(new_n536), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT110), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n623), .A2(new_n756), .A3(G472), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n753), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n541), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(KEYINPUT111), .A3(new_n541), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n750), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n288), .ZN(G24));
  NAND4_X1  g578(.A1(new_n725), .A2(new_n758), .A3(new_n688), .A4(new_n743), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT112), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n753), .B(new_n671), .C1(new_n755), .C2(new_n757), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n768), .A3(new_n725), .A4(new_n743), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  NAND2_X1  g585(.A1(KEYINPUT114), .A2(KEYINPUT42), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n445), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n444), .A2(KEYINPUT113), .A3(G469), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n686), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n506), .A2(new_n454), .A3(new_n507), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n680), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n618), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n772), .B1(new_n781), .B2(new_n726), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT114), .B(KEYINPUT42), .Z(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n780), .A2(new_n725), .A3(new_n618), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G131), .ZN(G33));
  NAND3_X1  g601(.A1(new_n780), .A2(new_n618), .A3(new_n700), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G134), .ZN(G36));
  AOI21_X1  g603(.A(new_n263), .B1(new_n637), .B2(new_n635), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT43), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OR3_X1    g606(.A1(new_n792), .A2(new_n624), .A3(new_n671), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n444), .A2(KEYINPUT45), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n444), .A2(KEYINPUT45), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(G469), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n452), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT46), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(KEYINPUT46), .A3(new_n452), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n450), .A3(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n803), .A2(new_n509), .A3(new_n719), .ZN(new_n804));
  INV_X1    g618(.A(new_n777), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n793), .B2(new_n794), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n795), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g622(.A(KEYINPUT115), .B(G137), .Z(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(G39));
  NAND2_X1  g624(.A1(new_n803), .A2(new_n509), .ZN(new_n811));
  AND2_X1   g625(.A1(KEYINPUT116), .A2(KEYINPUT47), .ZN(new_n812));
  NOR2_X1   g626(.A1(KEYINPUT116), .A2(KEYINPUT47), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n812), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n803), .A2(new_n509), .A3(new_n817), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n726), .A2(new_n678), .A3(new_n541), .A4(new_n777), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  AND4_X1   g639(.A1(new_n541), .A2(new_n706), .A3(new_n454), .A4(new_n509), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n731), .A2(new_n450), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT49), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n826), .A2(new_n713), .A3(new_n790), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n792), .A2(new_n690), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n732), .A2(new_n777), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n618), .A3(new_n831), .ZN(new_n832));
  XOR2_X1   g646(.A(KEYINPUT124), .B(KEYINPUT48), .Z(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n713), .A2(new_n541), .A3(new_n328), .ZN(new_n836));
  INV_X1    g650(.A(new_n831), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n838));
  OR3_X1    g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n836), .B2(new_n837), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n327), .B1(new_n841), .B2(new_n640), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n832), .A2(new_n834), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n761), .A2(new_n762), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n830), .A2(new_n743), .A3(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n835), .A2(new_n842), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n830), .A2(new_n767), .A3(new_n831), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n263), .A2(new_n638), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n839), .A2(new_n840), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n706), .A2(new_n707), .A3(new_n733), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT121), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n830), .A2(new_n852), .A3(new_n844), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n850), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n816), .A2(new_n818), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n827), .A2(new_n680), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n830), .A2(new_n844), .A3(new_n805), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT120), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n863), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n866), .A3(new_n861), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n858), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n861), .A2(KEYINPUT123), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n861), .A2(KEYINPUT123), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n872), .A3(new_n865), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n868), .B1(new_n873), .B2(new_n857), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n846), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n776), .A2(new_n509), .A3(new_n671), .A4(new_n695), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n713), .ZN(new_n878));
  INV_X1    g692(.A(new_n689), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n748), .A2(new_n878), .B1(new_n879), .B2(new_n725), .ZN(new_n880));
  AND4_X1   g694(.A1(KEYINPUT52), .A2(new_n770), .A3(new_n880), .A4(new_n703), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n766), .A2(new_n769), .B1(new_n697), .B2(new_n702), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT52), .B1(new_n882), .B2(new_n880), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n643), .A2(new_n333), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n627), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n655), .A2(KEYINPUT119), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n747), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n263), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT118), .B1(new_n890), .B2(new_n640), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n639), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n886), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n619), .B1(new_n344), .B2(new_n511), .ZN(new_n895));
  AOI211_X1 g709(.A(KEYINPUT95), .B(new_n510), .C1(new_n336), .C2(new_n343), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n897), .B2(new_n618), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n734), .B1(new_n742), .B2(new_n744), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n763), .A2(new_n899), .A3(new_n740), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n767), .A2(new_n725), .A3(new_n780), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n626), .B1(new_n605), .B2(new_n617), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n654), .A2(new_n671), .A3(new_n694), .A4(new_n777), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n887), .A4(new_n889), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n904), .A3(new_n788), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n785), .B2(new_n782), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n898), .A2(new_n900), .A3(new_n906), .A4(new_n673), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n876), .B1(new_n884), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n899), .A2(new_n740), .ZN(new_n909));
  INV_X1    g723(.A(new_n763), .ZN(new_n910));
  INV_X1    g724(.A(new_n905), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n786), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n891), .A2(new_n893), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n627), .A3(new_n885), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n621), .A2(new_n673), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n770), .A2(new_n880), .A3(new_n703), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT52), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n882), .A2(KEYINPUT52), .A3(new_n880), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n916), .A2(new_n921), .A3(KEYINPUT53), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n908), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n908), .A2(KEYINPUT54), .A3(new_n922), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n875), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(G952), .A2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n829), .B1(new_n927), .B2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n187), .A2(G952), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n495), .A2(new_n501), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(new_n499), .Z(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT55), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n884), .A2(new_n907), .A3(new_n876), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT53), .B1(new_n916), .B2(new_n921), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n536), .B(new_n505), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT56), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n536), .B1(new_n935), .B2(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT125), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n923), .A2(new_n942), .A3(new_n536), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n505), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(KEYINPUT126), .B(KEYINPUT56), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n933), .A2(new_n945), .ZN(new_n946));
  AOI211_X1 g760(.A(new_n930), .B(new_n939), .C1(new_n944), .C2(new_n946), .ZN(G51));
  AOI21_X1  g761(.A(new_n942), .B1(new_n923), .B2(new_n536), .ZN(new_n948));
  AOI211_X1 g762(.A(KEYINPUT125), .B(new_n318), .C1(new_n908), .C2(new_n922), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n798), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n451), .B(KEYINPUT57), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n925), .A2(new_n926), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n449), .B2(new_n448), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n930), .B1(new_n952), .B2(new_n955), .ZN(G54));
  AND2_X1   g770(.A1(KEYINPUT58), .A2(G475), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n255), .B1(new_n950), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n255), .A2(new_n957), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n941), .A2(new_n943), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n930), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n958), .A2(new_n962), .ZN(G60));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT59), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n925), .A2(new_n926), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n631), .A2(new_n633), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n961), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n966), .A2(new_n967), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT60), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n923), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n535), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n923), .A2(new_n669), .A3(new_n974), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(new_n961), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT61), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n976), .A2(KEYINPUT61), .A3(new_n961), .A4(new_n977), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(G66));
  AOI21_X1  g796(.A(new_n187), .B1(new_n330), .B2(G224), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n898), .A2(new_n900), .A3(new_n673), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n187), .ZN(new_n985));
  INV_X1    g799(.A(G898), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n931), .B1(new_n986), .B2(G953), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n985), .B(new_n987), .ZN(G69));
  INV_X1    g802(.A(new_n727), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n882), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n723), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n992));
  AOI22_X1  g806(.A1(new_n795), .A2(new_n807), .B1(new_n822), .B2(new_n823), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n618), .A2(new_n805), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n720), .B(new_n995), .C1(new_n891), .C2(new_n893), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT127), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n187), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n244), .A2(new_n245), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n590), .B(new_n1000), .Z(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(G900), .B2(G953), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n786), .A2(new_n788), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n748), .A2(new_n618), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1004), .B1(new_n804), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n993), .A2(new_n990), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1003), .B1(new_n1007), .B2(G953), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1010), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1002), .A2(new_n1012), .A3(new_n1008), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(G72));
  NAND2_X1  g828(.A1(G472), .A2(G902), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT63), .Z(new_n1016));
  OAI21_X1  g830(.A(new_n1016), .B1(new_n998), .B2(new_n984), .ZN(new_n1017));
  INV_X1    g831(.A(new_n591), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1017), .A2(new_n583), .A3(new_n1018), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n923), .B(new_n1016), .C1(new_n709), .C2(new_n609), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1016), .B1(new_n1007), .B2(new_n984), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1018), .A2(new_n583), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n930), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n1019), .A2(new_n1020), .A3(new_n1023), .ZN(G57));
endmodule


