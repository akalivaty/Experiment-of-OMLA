

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589;

  AND2_X1 U322 ( .A1(n570), .A2(n573), .ZN(n395) );
  INV_X1 U323 ( .A(n588), .ZN(n504) );
  NOR2_X1 U324 ( .A1(n484), .A2(n552), .ZN(n455) );
  XNOR2_X2 U325 ( .A(n394), .B(KEYINPUT41), .ZN(n573) );
  XNOR2_X1 U326 ( .A(G64GAT), .B(G92GAT), .ZN(n378) );
  XNOR2_X1 U327 ( .A(n434), .B(n433), .ZN(n435) );
  NOR2_X1 U328 ( .A1(n488), .A2(n487), .ZN(n506) );
  XNOR2_X1 U329 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U330 ( .A(n430), .B(n429), .Z(n290) );
  AND2_X1 U331 ( .A1(n392), .A2(n492), .ZN(n291) );
  XOR2_X1 U332 ( .A(n390), .B(n389), .Z(n292) );
  XNOR2_X1 U333 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U334 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n399) );
  XNOR2_X1 U335 ( .A(n432), .B(n376), .ZN(n377) );
  XNOR2_X1 U336 ( .A(n400), .B(n399), .ZN(n401) );
  INV_X1 U337 ( .A(KEYINPUT89), .ZN(n433) );
  NOR2_X1 U338 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U339 ( .A(n385), .B(n384), .ZN(n388) );
  XNOR2_X1 U340 ( .A(n391), .B(n292), .ZN(n492) );
  XNOR2_X1 U341 ( .A(n492), .B(KEYINPUT64), .ZN(n394) );
  INV_X1 U342 ( .A(G218GAT), .ZN(n459) );
  XNOR2_X1 U343 ( .A(n311), .B(n310), .ZN(n578) );
  XNOR2_X1 U344 ( .A(n459), .B(KEYINPUT62), .ZN(n460) );
  XNOR2_X1 U345 ( .A(n472), .B(KEYINPUT122), .ZN(n473) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U347 ( .A(n461), .B(n460), .ZN(G1355GAT) );
  XNOR2_X1 U348 ( .A(n474), .B(n473), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n496), .B(n495), .ZN(G1330GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n294) );
  XNOR2_X1 U351 ( .A(G106GAT), .B(G92GAT), .ZN(n293) );
  XNOR2_X1 U352 ( .A(n294), .B(n293), .ZN(n311) );
  XOR2_X1 U353 ( .A(KEYINPUT80), .B(KEYINPUT65), .Z(n296) );
  XNOR2_X1 U354 ( .A(G218GAT), .B(KEYINPUT81), .ZN(n295) );
  XNOR2_X1 U355 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U356 ( .A(n297), .B(KEYINPUT11), .Z(n299) );
  XOR2_X1 U357 ( .A(G99GAT), .B(G85GAT), .Z(n381) );
  XNOR2_X1 U358 ( .A(G134GAT), .B(n381), .ZN(n298) );
  XNOR2_X1 U359 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U360 ( .A(G36GAT), .B(G190GAT), .Z(n415) );
  XOR2_X1 U361 ( .A(KEYINPUT66), .B(n415), .Z(n301) );
  NAND2_X1 U362 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U363 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U364 ( .A(n303), .B(n302), .Z(n309) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n304) );
  XNOR2_X1 U366 ( .A(n304), .B(G29GAT), .ZN(n305) );
  XOR2_X1 U367 ( .A(n305), .B(KEYINPUT8), .Z(n307) );
  XNOR2_X1 U368 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n306) );
  XNOR2_X1 U369 ( .A(n307), .B(n306), .ZN(n352) );
  XOR2_X1 U370 ( .A(G50GAT), .B(G162GAT), .Z(n426) );
  XNOR2_X1 U371 ( .A(n352), .B(n426), .ZN(n308) );
  XNOR2_X1 U372 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U373 ( .A(KEYINPUT36), .B(n578), .Z(n489) );
  XOR2_X1 U374 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n313) );
  XNOR2_X1 U375 ( .A(G57GAT), .B(KEYINPUT96), .ZN(n312) );
  XNOR2_X1 U376 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U377 ( .A(KEYINPUT4), .B(n314), .Z(n316) );
  NAND2_X1 U378 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U379 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U380 ( .A(n317), .B(KEYINPUT97), .Z(n322) );
  XOR2_X1 U381 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n319) );
  XNOR2_X1 U382 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n318) );
  XNOR2_X1 U383 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U384 ( .A(G141GAT), .B(n320), .ZN(n439) );
  XOR2_X1 U385 ( .A(n439), .B(KEYINPUT98), .Z(n321) );
  XNOR2_X1 U386 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U387 ( .A(G85GAT), .B(G162GAT), .Z(n324) );
  XNOR2_X1 U388 ( .A(G29GAT), .B(G148GAT), .ZN(n323) );
  XNOR2_X1 U389 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U390 ( .A(n326), .B(n325), .Z(n334) );
  XOR2_X1 U391 ( .A(KEYINPUT0), .B(G134GAT), .Z(n328) );
  XNOR2_X1 U392 ( .A(KEYINPUT86), .B(G127GAT), .ZN(n327) );
  XNOR2_X1 U393 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U394 ( .A(G113GAT), .B(n329), .Z(n452) );
  XOR2_X1 U395 ( .A(KEYINPUT5), .B(G155GAT), .Z(n331) );
  XNOR2_X1 U396 ( .A(G1GAT), .B(G120GAT), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n452), .B(n332), .ZN(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n539) );
  INV_X1 U400 ( .A(KEYINPUT54), .ZN(n421) );
  XOR2_X1 U401 ( .A(G8GAT), .B(G113GAT), .Z(n336) );
  XNOR2_X1 U402 ( .A(G169GAT), .B(G197GAT), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U404 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n338) );
  XNOR2_X1 U405 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n337) );
  XNOR2_X1 U406 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U407 ( .A(n340), .B(n339), .Z(n347) );
  XOR2_X1 U408 ( .A(G36GAT), .B(G50GAT), .Z(n344) );
  XOR2_X1 U409 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n342) );
  XNOR2_X1 U410 ( .A(G15GAT), .B(G1GAT), .ZN(n341) );
  XNOR2_X1 U411 ( .A(n342), .B(n341), .ZN(n363) );
  XNOR2_X1 U412 ( .A(G22GAT), .B(n363), .ZN(n343) );
  XNOR2_X1 U413 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U414 ( .A(G141GAT), .B(n345), .ZN(n346) );
  XNOR2_X1 U415 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U416 ( .A(KEYINPUT75), .B(KEYINPUT67), .Z(n349) );
  NAND2_X1 U417 ( .A1(G229GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U419 ( .A(n351), .B(n350), .Z(n354) );
  XNOR2_X1 U420 ( .A(n352), .B(KEYINPUT70), .ZN(n353) );
  XOR2_X1 U421 ( .A(n354), .B(n353), .Z(n527) );
  INV_X1 U422 ( .A(n527), .ZN(n570) );
  XOR2_X1 U423 ( .A(KEYINPUT15), .B(KEYINPUT84), .Z(n356) );
  XNOR2_X1 U424 ( .A(G64GAT), .B(KEYINPUT85), .ZN(n355) );
  XNOR2_X1 U425 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U426 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n358) );
  XNOR2_X1 U427 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U429 ( .A(n360), .B(n359), .ZN(n371) );
  XOR2_X1 U430 ( .A(G8GAT), .B(G183GAT), .Z(n410) );
  XOR2_X1 U431 ( .A(G57GAT), .B(KEYINPUT13), .Z(n386) );
  XOR2_X1 U432 ( .A(n410), .B(n386), .Z(n362) );
  XNOR2_X1 U433 ( .A(G211GAT), .B(G78GAT), .ZN(n361) );
  XNOR2_X1 U434 ( .A(n362), .B(n361), .ZN(n367) );
  XOR2_X1 U435 ( .A(G22GAT), .B(G155GAT), .Z(n425) );
  XOR2_X1 U436 ( .A(n425), .B(n363), .Z(n365) );
  NAND2_X1 U437 ( .A1(G231GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U438 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U439 ( .A(n367), .B(n366), .Z(n369) );
  XNOR2_X1 U440 ( .A(G127GAT), .B(G71GAT), .ZN(n368) );
  XNOR2_X1 U441 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U442 ( .A(n371), .B(n370), .Z(n588) );
  NOR2_X1 U443 ( .A1(n504), .A2(n489), .ZN(n372) );
  XNOR2_X1 U444 ( .A(n372), .B(KEYINPUT45), .ZN(n392) );
  XOR2_X1 U445 ( .A(G120GAT), .B(G71GAT), .Z(n444) );
  XNOR2_X1 U446 ( .A(G106GAT), .B(G78GAT), .ZN(n373) );
  XNOR2_X1 U447 ( .A(n373), .B(G148GAT), .ZN(n432) );
  NAND2_X1 U448 ( .A1(G230GAT), .A2(G233GAT), .ZN(n375) );
  INV_X1 U449 ( .A(KEYINPUT31), .ZN(n374) );
  XNOR2_X1 U450 ( .A(n444), .B(n377), .ZN(n385) );
  INV_X1 U451 ( .A(n378), .ZN(n380) );
  XNOR2_X1 U452 ( .A(G176GAT), .B(G204GAT), .ZN(n379) );
  XNOR2_X1 U453 ( .A(n380), .B(n379), .ZN(n407) );
  XOR2_X1 U454 ( .A(n407), .B(n381), .Z(n383) );
  INV_X1 U455 ( .A(KEYINPUT78), .ZN(n382) );
  XNOR2_X1 U456 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U457 ( .A(n386), .B(KEYINPUT79), .ZN(n387) );
  XNOR2_X1 U458 ( .A(n388), .B(n387), .ZN(n391) );
  XOR2_X1 U459 ( .A(KEYINPUT77), .B(KEYINPUT33), .Z(n390) );
  XNOR2_X1 U460 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n389) );
  INV_X1 U461 ( .A(n492), .ZN(n584) );
  XNOR2_X1 U462 ( .A(n291), .B(KEYINPUT113), .ZN(n393) );
  NOR2_X1 U463 ( .A1(n570), .A2(n393), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n395), .B(KEYINPUT46), .ZN(n396) );
  NOR2_X1 U465 ( .A1(n588), .A2(n396), .ZN(n398) );
  INV_X1 U466 ( .A(n578), .ZN(n397) );
  NAND2_X1 U467 ( .A1(n398), .A2(n397), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n403), .B(KEYINPUT48), .ZN(n551) );
  XOR2_X1 U469 ( .A(KEYINPUT17), .B(KEYINPUT88), .Z(n405) );
  XNOR2_X1 U470 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U472 ( .A(G169GAT), .B(n406), .Z(n451) );
  XOR2_X1 U473 ( .A(KEYINPUT99), .B(n407), .Z(n409) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U476 ( .A(n411), .B(n410), .Z(n417) );
  XOR2_X1 U477 ( .A(KEYINPUT21), .B(G218GAT), .Z(n413) );
  XNOR2_X1 U478 ( .A(KEYINPUT91), .B(G211GAT), .ZN(n412) );
  XNOR2_X1 U479 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U480 ( .A(G197GAT), .B(n414), .Z(n430) );
  XNOR2_X1 U481 ( .A(n430), .B(n415), .ZN(n416) );
  XNOR2_X1 U482 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U483 ( .A(n451), .B(n418), .Z(n541) );
  INV_X1 U484 ( .A(n541), .ZN(n419) );
  NOR2_X1 U485 ( .A1(n551), .A2(n419), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n421), .B(n420), .ZN(n422) );
  NOR2_X1 U487 ( .A1(n539), .A2(n422), .ZN(n462) );
  XOR2_X1 U488 ( .A(KEYINPUT95), .B(KEYINPUT22), .Z(n424) );
  XNOR2_X1 U489 ( .A(KEYINPUT23), .B(KEYINPUT94), .ZN(n423) );
  XNOR2_X1 U490 ( .A(n424), .B(n423), .ZN(n438) );
  XOR2_X1 U491 ( .A(KEYINPUT90), .B(G204GAT), .Z(n428) );
  XNOR2_X1 U492 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U493 ( .A(n428), .B(n427), .ZN(n429) );
  NAND2_X1 U494 ( .A1(G228GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n290), .B(n431), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n432), .B(KEYINPUT24), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n484) );
  XOR2_X1 U499 ( .A(G176GAT), .B(G99GAT), .Z(n442) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(G190GAT), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U502 ( .A(n444), .B(n443), .Z(n446) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U505 ( .A(G183GAT), .B(KEYINPUT20), .Z(n448) );
  XNOR2_X1 U506 ( .A(G15GAT), .B(KEYINPUT87), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U508 ( .A(n450), .B(n449), .Z(n454) );
  XNOR2_X1 U509 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U510 ( .A(n454), .B(n453), .Z(n552) );
  XNOR2_X1 U511 ( .A(n455), .B(KEYINPUT26), .ZN(n568) );
  AND2_X1 U512 ( .A1(n462), .A2(n568), .ZN(n457) );
  INV_X1 U513 ( .A(KEYINPUT125), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n457), .B(n456), .ZN(n583) );
  INV_X1 U515 ( .A(n583), .ZN(n458) );
  NOR2_X1 U516 ( .A1(n489), .A2(n458), .ZN(n461) );
  INV_X1 U517 ( .A(n552), .ZN(n485) );
  NAND2_X1 U518 ( .A1(n462), .A2(n484), .ZN(n464) );
  INV_X1 U519 ( .A(KEYINPUT55), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n464), .B(n463), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n485), .A2(n465), .ZN(n466) );
  XNOR2_X1 U522 ( .A(n466), .B(KEYINPUT120), .ZN(n581) );
  NAND2_X1 U523 ( .A1(n581), .A2(n570), .ZN(n469) );
  INV_X1 U524 ( .A(KEYINPUT121), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n467), .B(G169GAT), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(G1348GAT) );
  NAND2_X1 U527 ( .A1(n581), .A2(n578), .ZN(n474) );
  XOR2_X1 U528 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n471) );
  XNOR2_X1 U529 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n541), .A2(n552), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n484), .A2(n475), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT25), .B(n476), .ZN(n480) );
  XOR2_X1 U534 ( .A(KEYINPUT27), .B(KEYINPUT100), .Z(n477) );
  XOR2_X1 U535 ( .A(n541), .B(n477), .Z(n482) );
  NAND2_X1 U536 ( .A1(n482), .A2(n568), .ZN(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT102), .B(n478), .Z(n479) );
  NOR2_X1 U538 ( .A1(n480), .A2(n479), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n539), .A2(n481), .ZN(n488) );
  NAND2_X1 U540 ( .A1(n482), .A2(n539), .ZN(n483) );
  XOR2_X1 U541 ( .A(KEYINPUT101), .B(n483), .Z(n550) );
  XOR2_X1 U542 ( .A(KEYINPUT28), .B(n484), .Z(n545) );
  INV_X1 U543 ( .A(n545), .ZN(n554) );
  NAND2_X1 U544 ( .A1(n554), .A2(n485), .ZN(n486) );
  NOR2_X1 U545 ( .A1(n550), .A2(n486), .ZN(n487) );
  NOR2_X1 U546 ( .A1(n506), .A2(n489), .ZN(n490) );
  NAND2_X1 U547 ( .A1(n504), .A2(n490), .ZN(n491) );
  XOR2_X1 U548 ( .A(KEYINPUT37), .B(n491), .Z(n538) );
  NAND2_X1 U549 ( .A1(n570), .A2(n492), .ZN(n509) );
  NOR2_X1 U550 ( .A1(n538), .A2(n509), .ZN(n493) );
  XOR2_X1 U551 ( .A(KEYINPUT38), .B(n493), .Z(n494) );
  XNOR2_X2 U552 ( .A(KEYINPUT107), .B(n494), .ZN(n525) );
  NAND2_X1 U553 ( .A1(n525), .A2(n552), .ZN(n496) );
  NAND2_X1 U554 ( .A1(n573), .A2(n581), .ZN(n499) );
  XOR2_X1 U555 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n497) );
  XNOR2_X1 U556 ( .A(n497), .B(G176GAT), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(G1349GAT) );
  NAND2_X1 U558 ( .A1(n583), .A2(n570), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n500), .B(KEYINPUT60), .ZN(n501) );
  XNOR2_X1 U560 ( .A(KEYINPUT59), .B(n501), .ZN(n503) );
  XOR2_X1 U561 ( .A(G197GAT), .B(KEYINPUT126), .Z(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(G1352GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT34), .B(KEYINPUT104), .Z(n512) );
  NOR2_X1 U564 ( .A1(n504), .A2(n578), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n505), .B(KEYINPUT16), .ZN(n508) );
  INV_X1 U566 ( .A(n506), .ZN(n507) );
  NAND2_X1 U567 ( .A1(n508), .A2(n507), .ZN(n529) );
  NOR2_X1 U568 ( .A1(n509), .A2(n529), .ZN(n510) );
  XOR2_X1 U569 ( .A(KEYINPUT103), .B(n510), .Z(n518) );
  NAND2_X1 U570 ( .A1(n518), .A2(n539), .ZN(n511) );
  XNOR2_X1 U571 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U572 ( .A(G1GAT), .B(n513), .Z(G1324GAT) );
  XOR2_X1 U573 ( .A(G8GAT), .B(KEYINPUT105), .Z(n515) );
  NAND2_X1 U574 ( .A1(n518), .A2(n541), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n515), .B(n514), .ZN(G1325GAT) );
  XOR2_X1 U576 ( .A(G15GAT), .B(KEYINPUT35), .Z(n517) );
  NAND2_X1 U577 ( .A1(n518), .A2(n552), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n517), .B(n516), .ZN(G1326GAT) );
  NAND2_X1 U579 ( .A1(n545), .A2(n518), .ZN(n519) );
  XNOR2_X1 U580 ( .A(n519), .B(KEYINPUT106), .ZN(n520) );
  XNOR2_X1 U581 ( .A(G22GAT), .B(n520), .ZN(G1327GAT) );
  XOR2_X1 U582 ( .A(G29GAT), .B(KEYINPUT39), .Z(n522) );
  NAND2_X1 U583 ( .A1(n539), .A2(n525), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n522), .B(n521), .ZN(G1328GAT) );
  NAND2_X1 U585 ( .A1(n525), .A2(n541), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(KEYINPUT108), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G36GAT), .B(n524), .ZN(G1329GAT) );
  NAND2_X1 U588 ( .A1(n545), .A2(n525), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G50GAT), .B(n526), .ZN(G1331GAT) );
  XNOR2_X1 U590 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n527), .A2(n573), .ZN(n528) );
  XOR2_X1 U592 ( .A(KEYINPUT109), .B(n528), .Z(n537) );
  NOR2_X1 U593 ( .A1(n529), .A2(n537), .ZN(n534) );
  NAND2_X1 U594 ( .A1(n539), .A2(n534), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1332GAT) );
  NAND2_X1 U596 ( .A1(n534), .A2(n541), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n532), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U598 ( .A1(n552), .A2(n534), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U600 ( .A(G78GAT), .B(KEYINPUT43), .Z(n536) );
  NAND2_X1 U601 ( .A1(n534), .A2(n545), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1335GAT) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n546) );
  NAND2_X1 U604 ( .A1(n546), .A2(n539), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n540), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U606 ( .A1(n546), .A2(n541), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(KEYINPUT110), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G92GAT), .B(n543), .ZN(G1337GAT) );
  NAND2_X1 U609 ( .A1(n552), .A2(n546), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n548) );
  NAND2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G106GAT), .B(n549), .ZN(G1339GAT) );
  NOR2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n567) );
  NAND2_X1 U616 ( .A1(n567), .A2(n552), .ZN(n553) );
  XOR2_X1 U617 ( .A(KEYINPUT114), .B(n553), .Z(n555) );
  NAND2_X1 U618 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U619 ( .A(n556), .B(KEYINPUT115), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n563), .A2(n570), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n557), .B(KEYINPUT116), .ZN(n558) );
  XNOR2_X1 U622 ( .A(G113GAT), .B(n558), .ZN(G1340GAT) );
  XOR2_X1 U623 ( .A(G120GAT), .B(KEYINPUT49), .Z(n560) );
  NAND2_X1 U624 ( .A1(n563), .A2(n573), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1341GAT) );
  NAND2_X1 U626 ( .A1(n588), .A2(n563), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(KEYINPUT50), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G127GAT), .B(n562), .ZN(G1342GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n578), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(G134GAT), .B(n566), .Z(G1343GAT) );
  XOR2_X1 U633 ( .A(G141GAT), .B(KEYINPUT119), .Z(n572) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT118), .B(n569), .Z(n579) );
  NAND2_X1 U636 ( .A1(n570), .A2(n579), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1344GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n575) );
  NAND2_X1 U639 ( .A1(n573), .A2(n579), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G148GAT), .B(n576), .ZN(G1345GAT) );
  NAND2_X1 U642 ( .A1(n579), .A2(n588), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n588), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U649 ( .A1(n583), .A2(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(G204GAT), .B(n587), .Z(G1353GAT) );
  NAND2_X1 U652 ( .A1(n588), .A2(n583), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
endmodule

