//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  AND3_X1   g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  OR3_X1    g0006(.A1(new_n206), .A2(KEYINPUT65), .A3(G13), .ZN(new_n207));
  OAI21_X1  g0007(.A(KEYINPUT65), .B1(new_n206), .B2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT67), .Z(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n223), .A2(G50), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n211), .B(new_n219), .C1(new_n222), .C2(new_n226), .ZN(G361));
  XOR2_X1   g0027(.A(G250), .B(G257), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT68), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n231), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G1698), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G232), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G238), .A3(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n249), .A2(G107), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT71), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n220), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n251), .A2(KEYINPUT71), .A3(new_n253), .A4(new_n254), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT69), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(new_n258), .B2(new_n220), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n267), .A2(KEYINPUT69), .A3(G1), .A4(G13), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n263), .A2(new_n266), .A3(G274), .A4(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n263), .A2(new_n265), .A3(new_n268), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n271), .B(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n270), .B1(new_n273), .B2(G244), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n261), .A2(new_n274), .A3(G190), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT72), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n275), .B(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n278), .A2(new_n220), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n264), .A2(G20), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G77), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n220), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n286), .A2(new_n288), .B1(new_n221), .B2(new_n202), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT15), .B(G87), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n221), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n285), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n284), .B(new_n293), .C1(G77), .C2(new_n280), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n261), .A2(new_n274), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(G200), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n277), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n261), .A2(new_n274), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n294), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT73), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n297), .A2(KEYINPUT73), .A3(new_n303), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n221), .B1(new_n201), .B2(new_n203), .ZN(new_n307));
  INV_X1    g0107(.A(G150), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n286), .A2(new_n291), .B1(new_n308), .B2(new_n288), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n285), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n280), .ZN(new_n311));
  INV_X1    g0111(.A(G50), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n283), .A2(G50), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n310), .B(new_n313), .C1(new_n281), .C2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT9), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n273), .A2(G226), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n252), .A2(G223), .A3(G1698), .ZN(new_n318));
  INV_X1    g0118(.A(G1698), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n252), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G222), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n318), .B1(new_n202), .B2(new_n252), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n270), .B1(new_n322), .B2(new_n259), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G200), .ZN(new_n325));
  INV_X1    g0125(.A(G190), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n316), .B(new_n325), .C1(new_n326), .C2(new_n324), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT10), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n325), .B2(KEYINPUT74), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n327), .B(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n324), .A2(new_n298), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n317), .A2(new_n323), .A3(new_n300), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(new_n315), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n305), .A2(new_n306), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G68), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n311), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT12), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n336), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n202), .B2(new_n291), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n282), .A2(G68), .A3(new_n283), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n338), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT11), .B1(new_n340), .B2(new_n285), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT14), .ZN(new_n347));
  NOR2_X1   g0147(.A1(G226), .A2(G1698), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n233), .B2(G1698), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n252), .B1(G33), .B2(G97), .ZN(new_n350));
  INV_X1    g0150(.A(new_n259), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n269), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n273), .B2(G238), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI211_X1 g0155(.A(KEYINPUT13), .B(new_n352), .C1(new_n273), .C2(G238), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n347), .B(G169), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n353), .B(new_n354), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n300), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n347), .B1(new_n358), .B2(G169), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n346), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(G200), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(new_n345), .C1(new_n326), .C2(new_n358), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n335), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(G58), .B(G68), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(G20), .B1(G159), .B2(new_n287), .ZN(new_n366));
  AOI21_X1  g0166(.A(G20), .B1(new_n246), .B2(new_n248), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  OAI21_X1  g0168(.A(G68), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n249), .A2(new_n370), .A3(new_n221), .ZN(new_n371));
  OAI211_X1 g0171(.A(KEYINPUT16), .B(new_n366), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n285), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n366), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n368), .A2(KEYINPUT75), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT75), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT7), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT76), .B1(new_n367), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT76), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(new_n370), .C1(new_n252), .C2(G20), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n247), .A2(KEYINPUT77), .A3(G33), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n246), .A2(KEYINPUT77), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n248), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n368), .A2(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n375), .B1(new_n389), .B2(G68), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n374), .B1(new_n390), .B2(KEYINPUT16), .ZN(new_n391));
  INV_X1    g0191(.A(new_n286), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n283), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n281), .B1(new_n393), .B2(KEYINPUT78), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n394), .A2(new_n395), .B1(new_n311), .B2(new_n286), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n391), .A2(KEYINPUT79), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT79), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n380), .A2(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n366), .B1(new_n399), .B2(new_n336), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n373), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n396), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n398), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n246), .A2(new_n248), .A3(G226), .A4(G1698), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT80), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n406), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n250), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n351), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n269), .B1(new_n271), .B2(new_n233), .ZN(new_n412));
  OAI21_X1  g0212(.A(G169), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n412), .ZN(new_n414));
  INV_X1    g0214(.A(G223), .ZN(new_n415));
  INV_X1    g0215(.A(G87), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n320), .A2(new_n415), .B1(new_n245), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n408), .B2(new_n407), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n414), .B(G179), .C1(new_n418), .C2(new_n351), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n397), .A2(new_n404), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n397), .A2(new_n404), .A3(new_n423), .A4(new_n420), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n402), .A2(new_n403), .ZN(new_n425));
  OAI21_X1  g0225(.A(G200), .B1(new_n411), .B2(new_n412), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n414), .B(G190), .C1(new_n418), .C2(new_n351), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT81), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n425), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n425), .A2(new_n428), .A3(new_n429), .A4(KEYINPUT17), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n422), .A2(new_n424), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n364), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(G97), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n311), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n264), .A2(G33), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n279), .A2(new_n280), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n440), .B2(new_n437), .ZN(new_n441));
  INV_X1    g0241(.A(G107), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(KEYINPUT6), .A3(G97), .ZN(new_n443));
  XOR2_X1   g0243(.A(G97), .B(G107), .Z(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(KEYINPUT6), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(G20), .B1(G77), .B2(new_n287), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n399), .B2(new_n442), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n441), .B1(new_n447), .B2(new_n285), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT82), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n246), .A2(new_n248), .A3(G244), .A4(new_n319), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT4), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n319), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n246), .A2(new_n248), .A3(G250), .A4(G1698), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n453), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT83), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n456), .A2(new_n455), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT83), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n454), .A4(new_n453), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n259), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT84), .ZN(new_n464));
  INV_X1    g0264(.A(G41), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(KEYINPUT84), .B2(G41), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n471), .A2(new_n263), .A3(new_n268), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(KEYINPUT85), .A3(G257), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n471), .A2(G257), .A3(new_n263), .A4(new_n268), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT85), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n263), .A2(G274), .A3(new_n268), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n473), .A2(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n463), .A2(new_n326), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(new_n476), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n477), .A2(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n351), .B1(new_n458), .B2(new_n461), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n480), .B1(new_n485), .B2(G200), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n463), .A2(G179), .A3(new_n479), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n485), .B2(new_n298), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n447), .A2(new_n285), .ZN(new_n489));
  INV_X1    g0289(.A(new_n441), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n450), .A2(new_n486), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n246), .A2(new_n248), .A3(G250), .A4(new_n319), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT95), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT95), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n252), .A2(new_n495), .A3(G250), .A4(new_n319), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n246), .A2(new_n248), .A3(G257), .A4(G1698), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G294), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n494), .A2(new_n496), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT96), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n497), .A2(new_n498), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT96), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(new_n494), .A4(new_n496), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n259), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n472), .A2(G264), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n482), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n298), .ZN(new_n507));
  OR3_X1    g0307(.A1(new_n280), .A2(KEYINPUT25), .A3(G107), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT25), .B1(new_n280), .B2(G107), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n509), .C1(new_n440), .C2(new_n442), .ZN(new_n510));
  XOR2_X1   g0310(.A(new_n510), .B(KEYINPUT94), .Z(new_n511));
  XNOR2_X1  g0311(.A(KEYINPUT92), .B(KEYINPUT22), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT93), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n416), .A2(G20), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n252), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G116), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n245), .A2(new_n516), .A3(G20), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT23), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n221), .B2(G107), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n442), .A2(KEYINPUT23), .A3(G20), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n252), .A2(new_n512), .A3(new_n514), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT93), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT22), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n252), .B2(new_n514), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n515), .B(new_n521), .C1(new_n523), .C2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT24), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n521), .A2(new_n515), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n529), .B(KEYINPUT24), .C1(new_n525), .C2(new_n523), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n530), .A3(new_n285), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n511), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n505), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n351), .B1(new_n499), .B2(KEYINPUT96), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n503), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(new_n300), .A3(new_n482), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n507), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n263), .A2(G274), .A3(new_n268), .A4(new_n470), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT86), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n246), .A2(new_n248), .A3(G244), .A4(G1698), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n246), .A2(new_n248), .A3(G238), .A4(new_n319), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(new_n245), .C2(new_n516), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n263), .A2(new_n268), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT87), .B1(new_n469), .B2(G1), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT87), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(new_n264), .A3(G45), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n544), .A2(new_n546), .A3(G250), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n542), .A2(new_n259), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(G169), .B1(new_n539), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n539), .A2(new_n548), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(new_n300), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G97), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n221), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G97), .A2(G107), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n416), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n336), .A2(G20), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n221), .A2(G33), .A3(G97), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n252), .A2(new_n558), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n285), .ZN(new_n562));
  INV_X1    g0362(.A(new_n290), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(new_n280), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT89), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n279), .B1(new_n557), .B2(new_n560), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT89), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n567), .A2(new_n568), .A3(new_n564), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n566), .A2(new_n569), .B1(new_n290), .B2(new_n440), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n551), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n440), .A2(new_n416), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n562), .A2(KEYINPUT89), .A3(new_n565), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n568), .B1(new_n567), .B2(new_n564), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n539), .A2(new_n548), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G200), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n539), .A2(G190), .A3(new_n548), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n537), .A2(new_n571), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n506), .A2(G200), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n535), .A2(G190), .A3(new_n482), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n511), .A4(new_n531), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n246), .A2(new_n248), .A3(G264), .A4(G1698), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n246), .A2(new_n248), .A3(G257), .A4(new_n319), .ZN(new_n585));
  INV_X1    g0385(.A(G303), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n584), .B(new_n585), .C1(new_n586), .C2(new_n252), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n259), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n471), .A2(G270), .A3(new_n263), .A4(new_n268), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n482), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT90), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n455), .B(new_n221), .C1(G33), .C2(new_n437), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n516), .A2(G20), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n285), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT20), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n280), .A2(G116), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n279), .A2(new_n280), .A3(new_n439), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(G116), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n298), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(KEYINPUT91), .A2(KEYINPUT21), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n588), .A2(new_n482), .A3(KEYINPUT90), .A4(new_n589), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n592), .A2(new_n601), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n590), .A2(new_n300), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n597), .A2(new_n600), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n263), .A2(G274), .A3(new_n268), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n589), .B1(new_n610), .B2(new_n471), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT90), .B1(new_n612), .B2(new_n588), .ZN(new_n613));
  INV_X1    g0413(.A(new_n604), .ZN(new_n614));
  OAI21_X1  g0414(.A(G190), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n607), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n592), .A2(G200), .A3(new_n604), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n592), .A2(new_n604), .A3(new_n601), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n602), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n609), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n492), .A2(new_n580), .A3(new_n583), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n436), .A2(new_n622), .ZN(G372));
  NAND2_X1  g0423(.A1(new_n573), .A2(new_n574), .ZN(new_n624));
  INV_X1    g0424(.A(new_n572), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n624), .A2(new_n625), .A3(new_n578), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT97), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n576), .B2(G200), .ZN(new_n628));
  INV_X1    g0428(.A(G200), .ZN(new_n629));
  AOI211_X1 g0429(.A(KEYINPUT97), .B(new_n629), .C1(new_n539), .C2(new_n548), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n626), .A2(new_n631), .B1(new_n570), .B2(new_n551), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n491), .A2(new_n449), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n448), .A2(KEYINPUT82), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n486), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n487), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n298), .B1(new_n463), .B2(new_n479), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n491), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n632), .A2(new_n635), .A3(new_n583), .A4(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n537), .A2(new_n620), .A3(new_n609), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n571), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n637), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(new_n487), .B1(new_n633), .B2(new_n634), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT26), .B1(new_n643), .B2(new_n632), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n571), .A2(new_n579), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n645), .A2(new_n638), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n435), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n333), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n391), .A2(new_n396), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n420), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT18), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n423), .A3(new_n420), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n363), .A2(new_n303), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(new_n361), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n432), .A2(new_n433), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n654), .B(new_n655), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n651), .B1(new_n659), .B2(new_n330), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n650), .A2(new_n660), .ZN(G369));
  NAND3_X1  g0461(.A1(new_n620), .A2(new_n608), .A3(new_n605), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n264), .A2(new_n221), .A3(G13), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(KEYINPUT98), .B(G343), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n616), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT99), .B1(new_n662), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n609), .A2(new_n618), .A3(new_n620), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n671), .B1(new_n672), .B2(new_n670), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n662), .A2(KEYINPUT99), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  INV_X1    g0477(.A(new_n669), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n532), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n583), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n680), .A2(new_n537), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n537), .A2(new_n678), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n662), .A2(new_n669), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n682), .B1(new_n683), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n689), .ZN(G399));
  INV_X1    g0490(.A(new_n209), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n555), .A2(new_n416), .A3(new_n516), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n692), .A2(new_n264), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n226), .B2(new_n692), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  INV_X1    g0496(.A(KEYINPUT100), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n535), .A2(new_n550), .A3(new_n606), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n463), .A2(new_n479), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n592), .A2(new_n576), .A3(new_n300), .A4(new_n604), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n485), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n700), .A2(KEYINPUT30), .B1(new_n702), .B2(new_n506), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n697), .B(new_n704), .C1(new_n698), .C2(new_n699), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n669), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n622), .A2(new_n678), .B1(new_n706), .B2(KEYINPUT31), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n700), .A2(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n506), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(G330), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT101), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT31), .B1(new_n710), .B2(new_n678), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n716), .B(new_n711), .C1(new_n622), .C2(new_n678), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT101), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(G330), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n633), .A2(new_n634), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n488), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n577), .A2(KEYINPUT97), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n576), .A2(new_n627), .A3(G200), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n575), .A2(new_n578), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n571), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT26), .B1(new_n722), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n448), .B1(new_n642), .B2(new_n487), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(new_n646), .A3(new_n571), .A4(new_n579), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n669), .B1(new_n641), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n649), .A2(new_n669), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(KEYINPUT29), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n720), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n696), .B1(new_n736), .B2(G1), .ZN(G364));
  INV_X1    g0537(.A(G13), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n264), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n692), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n221), .A2(G179), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G190), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G159), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT32), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n743), .A2(new_n326), .A3(G200), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n749), .B1(new_n442), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(G20), .A2(G179), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G58), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n752), .A2(new_n326), .A3(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n252), .B1(new_n754), .B2(new_n202), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n326), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n221), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n437), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n416), .ZN(new_n763));
  NOR4_X1   g0563(.A1(new_n751), .A2(new_n758), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n752), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(G190), .A3(G200), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n747), .A2(new_n748), .B1(new_n312), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n765), .A2(new_n326), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n767), .B1(G68), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G283), .ZN(new_n771));
  INV_X1    g0571(.A(G329), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n750), .A2(new_n771), .B1(new_n745), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT104), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n756), .A2(G322), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n775), .B(new_n249), .C1(new_n754), .C2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  INV_X1    g0578(.A(G326), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n760), .A2(new_n778), .B1(new_n766), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  OAI22_X1  g0581(.A1(new_n768), .A2(new_n781), .B1(new_n762), .B2(new_n586), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n777), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n764), .A2(new_n770), .B1(new_n774), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n220), .B1(G20), .B2(new_n298), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n742), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n209), .A2(G355), .A3(new_n252), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n691), .A2(new_n252), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n469), .B2(new_n226), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(KEYINPUT102), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n469), .B2(new_n243), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(KEYINPUT102), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n788), .B1(G116), .B2(new_n209), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n738), .A2(new_n245), .A3(KEYINPUT103), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT103), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(G13), .B2(G33), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n785), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n787), .B1(new_n795), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n801), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n676), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n676), .A2(G330), .ZN(new_n806));
  INV_X1    g0606(.A(new_n742), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n677), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(G396));
  INV_X1    g0609(.A(new_n720), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n302), .A2(new_n678), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n277), .A2(new_n296), .B1(new_n294), .B2(new_n678), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n813), .B2(new_n303), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n734), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n277), .A2(new_n296), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n294), .A2(new_n678), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n811), .B1(new_n818), .B2(new_n302), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n819), .B(new_n669), .C1(new_n641), .C2(new_n648), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n742), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n810), .B2(new_n821), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n799), .A2(new_n785), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT105), .Z(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n807), .B1(new_n826), .B2(new_n202), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G143), .A2(new_n756), .B1(new_n753), .B2(G159), .ZN(new_n828));
  INV_X1    g0628(.A(G137), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n829), .B2(new_n766), .C1(new_n308), .C2(new_n768), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT34), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n750), .A2(new_n336), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n252), .B1(new_n745), .B2(new_n834), .C1(new_n312), .C2(new_n762), .ZN(new_n835));
  INV_X1    g0635(.A(new_n760), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n833), .B(new_n835), .C1(G58), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n830), .A2(new_n831), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n832), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n750), .A2(new_n416), .B1(new_n766), .B2(new_n586), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n761), .B(new_n840), .C1(G283), .C2(new_n769), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n249), .B1(new_n762), .B2(new_n442), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT106), .Z(new_n843));
  OAI22_X1  g0643(.A1(new_n754), .A2(new_n516), .B1(new_n745), .B2(new_n776), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G294), .B2(new_n756), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n841), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n827), .B1(new_n786), .B2(new_n847), .C1(new_n819), .C2(new_n800), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n823), .A2(new_n848), .ZN(G384));
  OAI211_X1 g0649(.A(G116), .B(new_n222), .C1(new_n445), .C2(KEYINPUT35), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n850), .A2(KEYINPUT107), .B1(KEYINPUT35), .B2(new_n445), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(KEYINPUT107), .B2(new_n850), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT36), .Z(new_n853));
  OAI211_X1 g0653(.A(new_n226), .B(G77), .C1(new_n755), .C2(new_n336), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n201), .A2(G68), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n264), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  AND4_X1   g0657(.A1(new_n580), .A2(new_n492), .A3(new_n583), .A4(new_n621), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n715), .B1(new_n858), .B2(new_n669), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n711), .A2(KEYINPUT112), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT112), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n706), .A2(new_n861), .A3(KEYINPUT31), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n436), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n345), .A2(new_n669), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n361), .A2(new_n363), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n866), .B1(new_n361), .B2(new_n363), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n819), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n859), .B2(new_n863), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n397), .A2(new_n404), .A3(new_n667), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n425), .A2(new_n428), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n421), .A2(new_n871), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n871), .A2(new_n873), .A3(new_n653), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n872), .ZN(new_n876));
  INV_X1    g0676(.A(new_n871), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n654), .A2(new_n655), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n658), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(KEYINPUT110), .B(KEYINPUT38), .Z(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n367), .A2(new_n370), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n884), .B(G68), .C1(new_n368), .C2(new_n367), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT16), .B1(new_n885), .B2(new_n366), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n396), .B1(new_n373), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT108), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT108), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n396), .B(new_n889), .C1(new_n373), .C2(new_n886), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n667), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n434), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n888), .A2(new_n420), .A3(new_n890), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n873), .A2(new_n891), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n894), .B1(new_n874), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT111), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n893), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n899), .B1(new_n893), .B2(new_n898), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n883), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n870), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT40), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT109), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n893), .A2(new_n898), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n893), .B2(new_n898), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n874), .A2(new_n897), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n893), .A2(new_n909), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n907), .A2(new_n908), .B1(new_n910), .B2(KEYINPUT38), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n870), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n904), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n864), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n864), .A2(new_n914), .ZN(new_n916));
  INV_X1    g0716(.A(G330), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(new_n883), .C1(new_n900), .C2(new_n901), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n893), .B2(new_n909), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n893), .A2(new_n898), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT109), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n921), .B1(new_n923), .B2(new_n906), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n920), .B1(new_n924), .B2(new_n919), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n361), .A2(new_n678), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n361), .A2(new_n363), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n865), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n361), .A2(new_n363), .A3(new_n866), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n812), .B2(new_n820), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(new_n911), .B1(new_n878), .B2(new_n666), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n435), .A2(new_n735), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n660), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n936), .B(new_n938), .Z(new_n939));
  OAI22_X1  g0739(.A1(new_n918), .A2(new_n939), .B1(new_n264), .B2(new_n739), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n918), .A2(new_n939), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n857), .B1(new_n940), .B2(new_n941), .ZN(G367));
  OAI21_X1  g0742(.A(new_n802), .B1(new_n209), .B2(new_n290), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n231), .B2(new_n789), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT115), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n249), .B1(new_n754), .B2(new_n771), .ZN(new_n946));
  INV_X1    g0746(.A(G317), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n757), .A2(new_n586), .B1(new_n745), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n762), .A2(new_n516), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n946), .B(new_n948), .C1(KEYINPUT46), .C2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(KEYINPUT46), .B2(new_n949), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n750), .A2(new_n437), .B1(new_n768), .B2(new_n778), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n760), .A2(new_n442), .B1(new_n766), .B2(new_n776), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n750), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(G77), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n956), .B1(new_n755), .B2(new_n762), .C1(new_n336), .C2(new_n760), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n252), .B1(new_n757), .B2(new_n308), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n754), .A2(new_n201), .B1(new_n829), .B2(new_n745), .ZN(new_n959));
  INV_X1    g0759(.A(G143), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n960), .A2(new_n766), .B1(new_n768), .B2(new_n746), .ZN(new_n961));
  NOR4_X1   g0761(.A1(new_n957), .A2(new_n958), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT47), .Z(new_n964));
  AOI211_X1 g0764(.A(new_n807), .B(new_n945), .C1(new_n964), .C2(new_n785), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT116), .Z(new_n966));
  OR3_X1    g0766(.A1(new_n571), .A2(new_n575), .A3(new_n669), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n575), .A2(new_n669), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n727), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n966), .B1(new_n804), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n740), .B(KEYINPUT114), .Z(new_n971));
  OAI21_X1  g0771(.A(new_n492), .B1(new_n450), .B2(new_n669), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n643), .A2(new_n678), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n689), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT45), .B1(new_n689), .B2(new_n974), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT113), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n978), .B(KEYINPUT44), .C1(new_n689), .C2(new_n974), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n978), .A2(KEYINPUT44), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n978), .A2(KEYINPUT44), .ZN(new_n981));
  OR4_X1    g0781(.A1(new_n689), .A2(new_n974), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n977), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(new_n685), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n685), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n683), .B(new_n687), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(new_n677), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n736), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n736), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n692), .B(KEYINPUT41), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n971), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n993));
  INV_X1    g0793(.A(new_n974), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n638), .B1(new_n994), .B2(new_n537), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n669), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n683), .A2(new_n688), .ZN(new_n997));
  OAI21_X1  g0797(.A(KEYINPUT42), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n997), .A2(new_n994), .A3(KEYINPUT42), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n993), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n685), .A2(new_n974), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n970), .B1(new_n992), .B2(new_n1005), .ZN(G387));
  INV_X1    g0806(.A(new_n762), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n836), .A2(G283), .B1(new_n1007), .B2(G294), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G303), .A2(new_n753), .B1(new_n756), .B2(G317), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(KEYINPUT117), .B(G322), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1009), .B1(new_n776), .B2(new_n768), .C1(new_n766), .C2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT118), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1008), .B1(new_n1013), .B2(KEYINPUT48), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(KEYINPUT48), .B2(new_n1013), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT49), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n249), .B1(new_n745), .B2(new_n779), .C1(new_n516), .C2(new_n750), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n249), .B1(G50), .B2(new_n756), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n336), .B2(new_n754), .C1(new_n308), .C2(new_n745), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n836), .A2(new_n563), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n286), .B2(new_n768), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n762), .A2(new_n202), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n750), .A2(new_n437), .B1(new_n766), .B2(new_n746), .ZN(new_n1024));
  NOR4_X1   g0824(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n785), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n236), .A2(new_n469), .A3(new_n252), .ZN(new_n1027));
  OR3_X1    g0827(.A1(new_n286), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1028));
  OAI21_X1  g0828(.A(KEYINPUT50), .B1(new_n286), .B2(G50), .ZN(new_n1029));
  AOI21_X1  g0829(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n693), .B1(new_n1031), .B2(new_n249), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1033), .A2(new_n691), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n802), .B1(new_n442), .B2(new_n209), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1026), .B(new_n742), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n684), .B2(new_n801), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n988), .B2(new_n971), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n989), .A2(new_n692), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n736), .A2(new_n988), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(G393));
  NAND3_X1  g0841(.A1(new_n984), .A2(new_n985), .A3(new_n971), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n790), .A2(new_n240), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n802), .B1(new_n437), .B2(new_n209), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n742), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n754), .A2(new_n286), .B1(new_n201), .B2(new_n768), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT119), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1046), .A2(new_n1047), .B1(new_n202), .B2(new_n760), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1047), .B2(new_n1046), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT120), .Z(new_n1050));
  OAI22_X1  g0850(.A1(new_n757), .A2(new_n746), .B1(new_n766), .B2(new_n308), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT51), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n252), .B1(new_n745), .B2(new_n960), .C1(new_n416), .C2(new_n750), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G68), .B2(new_n1007), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1050), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n766), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1056), .A2(G317), .B1(G311), .B2(new_n756), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n249), .B1(new_n745), .B2(new_n1010), .C1(new_n754), .C2(new_n778), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n750), .A2(new_n442), .B1(new_n768), .B2(new_n586), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n760), .A2(new_n516), .B1(new_n762), .B2(new_n771), .ZN(new_n1061));
  OR3_X1    g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1055), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1045), .B1(new_n1063), .B2(new_n785), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n974), .B2(new_n804), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n986), .A2(new_n989), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n692), .B1(new_n986), .B2(new_n989), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1042), .B(new_n1065), .C1(new_n1066), .C2(new_n1067), .ZN(G390));
  NAND2_X1  g0868(.A1(new_n818), .A2(new_n302), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n669), .B(new_n1069), .C1(new_n641), .C2(new_n731), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1070), .A2(new_n812), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n926), .B(new_n902), .C1(new_n1071), .C2(new_n933), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n820), .A2(new_n812), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n927), .B1(new_n1073), .B2(new_n932), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1072), .B1(new_n925), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n917), .B1(new_n859), .B2(new_n863), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n814), .B1(new_n930), .B2(new_n931), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(KEYINPUT121), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n720), .A2(new_n819), .A3(new_n932), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1082), .B(new_n1072), .C1(new_n925), .C2(new_n1074), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT121), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1075), .A2(new_n1084), .A3(new_n1079), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1081), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n814), .B1(new_n714), .B2(new_n719), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1078), .B1(new_n1087), .B2(new_n932), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n1073), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n861), .B1(new_n706), .B2(KEYINPUT31), .ZN(new_n1090));
  AND4_X1   g0890(.A1(new_n861), .A2(new_n710), .A3(KEYINPUT31), .A4(new_n678), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(KEYINPUT122), .B(G330), .C1(new_n1092), .C2(new_n707), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n819), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1076), .A2(KEYINPUT122), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n933), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n1071), .A3(new_n1082), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1089), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n435), .A2(new_n1076), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n937), .A2(new_n1099), .A3(new_n660), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1086), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1100), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1104), .A2(new_n1081), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n692), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1085), .A2(new_n1083), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1084), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n925), .A2(new_n800), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n742), .B1(new_n825), .B2(new_n392), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n760), .A2(new_n202), .B1(new_n766), .B2(new_n771), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G107), .B2(new_n769), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n252), .B1(G116), .B2(new_n756), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n745), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1115), .A2(G294), .B1(G97), .B2(new_n753), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n763), .A2(new_n833), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1007), .A2(G150), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT53), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n836), .A2(G159), .B1(new_n1056), .B2(G128), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n201), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1122), .A2(new_n955), .B1(new_n769), .B2(G137), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n249), .B1(new_n1115), .B2(G125), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1126), .A2(new_n753), .B1(G132), .B2(new_n756), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1118), .B1(new_n1120), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1111), .B1(new_n1129), .B2(new_n785), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1109), .A2(new_n971), .B1(new_n1110), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1106), .A2(new_n1131), .ZN(G378));
  AOI21_X1  g0932(.A(new_n1100), .B1(new_n1109), .B2(new_n1104), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n936), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1077), .B1(new_n1092), .B2(new_n707), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n924), .A2(new_n1135), .A3(KEYINPUT40), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n912), .B1(new_n870), .B2(new_n902), .ZN(new_n1137));
  OAI21_X1  g0937(.A(G330), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n315), .A2(new_n667), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n334), .B(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n914), .A2(G330), .A3(new_n1142), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1134), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1134), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT57), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n692), .B1(new_n1133), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1101), .B1(new_n1086), .B2(new_n1102), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n936), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1134), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT57), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1149), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1143), .A2(new_n799), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1122), .A2(new_n799), .A3(new_n785), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n760), .A2(new_n336), .B1(new_n766), .B2(new_n516), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT123), .Z(new_n1160));
  NAND2_X1  g0960(.A1(new_n249), .A2(new_n465), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G107), .B2(new_n756), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1115), .A2(G283), .B1(new_n563), .B2(new_n753), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n750), .A2(new_n755), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1023), .B(new_n1164), .C1(G97), .C2(new_n769), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1160), .A2(new_n1162), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT58), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1161), .B(new_n312), .C1(G33), .C2(G41), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(G125), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1171), .A2(new_n766), .B1(new_n768), .B2(new_n834), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G128), .A2(new_n756), .B1(new_n753), .B2(G137), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n762), .B2(new_n1125), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(G150), .C2(new_n836), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n955), .A2(G159), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G33), .B(G41), .C1(new_n1115), .C2(G124), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1170), .B1(KEYINPUT58), .B2(new_n1167), .C1(new_n1177), .C2(new_n1181), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n807), .B(new_n1158), .C1(new_n1182), .C2(new_n785), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1154), .A2(new_n971), .B1(new_n1157), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1156), .A2(new_n1184), .ZN(G375));
  NAND3_X1  g0985(.A1(new_n1089), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1102), .A2(new_n991), .A3(new_n1186), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT124), .Z(new_n1188));
  OAI22_X1  g0988(.A1(new_n757), .A2(new_n771), .B1(new_n754), .B2(new_n442), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n252), .B(new_n1189), .C1(G303), .C2(new_n1115), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n516), .A2(new_n768), .B1(new_n766), .B2(new_n778), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G97), .B2(new_n1007), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1190), .A2(new_n956), .A3(new_n1021), .A4(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n760), .A2(new_n312), .B1(new_n762), .B2(new_n746), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G132), .B2(new_n1056), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n249), .B1(new_n1115), .B2(G128), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G137), .A2(new_n756), .B1(new_n753), .B2(G150), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1164), .B1(new_n769), .B2(new_n1126), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n786), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n807), .B(new_n1200), .C1(new_n336), .C2(new_n826), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n932), .B2(new_n800), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1071), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1087), .B2(new_n932), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1073), .A2(new_n1088), .B1(new_n1204), .B2(new_n1096), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n971), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1202), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1188), .A2(new_n1208), .ZN(G381));
  INV_X1    g1009(.A(G375), .ZN(new_n1210));
  INV_X1    g1010(.A(G390), .ZN(new_n1211));
  INV_X1    g1011(.A(G384), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(G393), .A2(G396), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(new_n1213), .A2(G387), .A3(G378), .A4(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1210), .A2(new_n1215), .A3(new_n1208), .A4(new_n1188), .ZN(G407));
  NAND2_X1  g1016(.A1(new_n1110), .A2(new_n1130), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1086), .B2(new_n1206), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n692), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1086), .B2(new_n1102), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1218), .B1(new_n1105), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(G213), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n668), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1210), .A2(new_n1221), .A3(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(G407), .A2(G213), .A3(new_n1224), .ZN(G409));
  XNOR2_X1  g1025(.A(G393), .B(G396), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT126), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1226), .A2(KEYINPUT126), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G387), .A2(new_n1211), .ZN(new_n1229));
  OAI211_X1 g1029(.A(G390), .B(new_n970), .C1(new_n992), .C2(new_n1005), .ZN(new_n1230));
  AND4_X1   g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1227), .A2(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT60), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1186), .B1(new_n1104), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1205), .A2(KEYINPUT60), .A3(new_n1100), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n692), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT125), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT125), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1235), .A2(new_n1239), .A3(new_n692), .A4(new_n1236), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G384), .B1(new_n1241), .B2(new_n1208), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1212), .B(new_n1207), .C1(new_n1238), .C2(new_n1240), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G378), .B(new_n1184), .C1(new_n1149), .C2(new_n1155), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1150), .A2(new_n991), .A3(new_n1154), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1154), .A2(new_n971), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1157), .A2(new_n1183), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1221), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1223), .B1(new_n1245), .B2(new_n1250), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1244), .A2(KEYINPUT62), .A3(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT62), .B1(new_n1244), .B2(new_n1251), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT127), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1245), .A2(new_n1250), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1223), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT60), .B1(new_n1205), .B2(new_n1100), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1219), .B1(new_n1258), .B2(new_n1186), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1239), .B1(new_n1259), .B2(new_n1236), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1240), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1208), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1212), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1241), .A2(G384), .A3(new_n1208), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1256), .A2(new_n1257), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT62), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1254), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1223), .A2(G2897), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1263), .A2(new_n1264), .A3(new_n1269), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1267), .A2(new_n1268), .A3(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1233), .B1(new_n1255), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT63), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1233), .B1(new_n1277), .B2(new_n1265), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1244), .A2(KEYINPUT63), .A3(new_n1251), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(new_n1268), .A3(new_n1274), .A4(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(G405));
  NAND2_X1  g1081(.A1(G375), .A2(new_n1221), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1245), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1244), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1282), .B(new_n1245), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(new_n1233), .ZN(G402));
endmodule


