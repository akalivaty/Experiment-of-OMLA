//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1037, new_n1038,
    new_n1039;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT16), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(new_n203), .B2(new_n202), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(G8gat), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G71gat), .B(G78gat), .Z(new_n208));
  NAND2_X1  g007(.A1(KEYINPUT97), .A2(KEYINPUT9), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G57gat), .B(G64gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n208), .B(new_n209), .C1(new_n212), .C2(new_n211), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT98), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT98), .B1(new_n214), .B2(new_n215), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT21), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n207), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G127gat), .B(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G231gat), .ZN(new_n224));
  INV_X1    g023(.A(G233gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n218), .A2(new_n219), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n227), .B1(new_n218), .B2(new_n219), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n223), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n230), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n228), .A3(new_n222), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT99), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n231), .B2(new_n233), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n221), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n231), .A2(new_n233), .ZN(new_n240));
  INV_X1    g039(.A(new_n235), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(new_n220), .A3(new_n236), .ZN(new_n243));
  XOR2_X1   g042(.A(G183gat), .B(G211gat), .Z(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n239), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n245), .B1(new_n239), .B2(new_n243), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G190gat), .B(G218gat), .ZN(new_n249));
  OR3_X1    g048(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n252), .B2(KEYINPUT91), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(KEYINPUT91), .B2(new_n250), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT92), .B(G29gat), .Z(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G36gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G50gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G43gat), .ZN(new_n259));
  INV_X1    g058(.A(G43gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G50gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT15), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  OR3_X1    g063(.A1(new_n258), .A2(KEYINPUT94), .A3(G43gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(KEYINPUT94), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n259), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT15), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n255), .A2(G36gat), .B1(new_n250), .B2(new_n251), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n262), .A2(KEYINPUT93), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n262), .A2(KEYINPUT93), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n269), .A2(new_n270), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT17), .B1(new_n264), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G99gat), .A2(G106gat), .ZN(new_n275));
  INV_X1    g074(.A(G85gat), .ZN(new_n276));
  INV_X1    g075(.A(G92gat), .ZN(new_n277));
  AOI22_X1  g076(.A1(KEYINPUT8), .A2(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n276), .B2(new_n277), .ZN(new_n280));
  NAND4_X1  g079(.A1(KEYINPUT101), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G99gat), .B(G106gat), .Z(new_n283));
  OR2_X1    g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n264), .A2(KEYINPUT17), .A3(new_n273), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT95), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n264), .A2(KEYINPUT95), .A3(KEYINPUT17), .A4(new_n273), .ZN(new_n291));
  AOI211_X1 g090(.A(new_n274), .B(new_n287), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n264), .A2(new_n273), .ZN(new_n293));
  NAND2_X1  g092(.A1(G232gat), .A2(G233gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n293), .A2(new_n287), .B1(KEYINPUT41), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n249), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n274), .B1(new_n290), .B2(new_n291), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n286), .ZN(new_n300));
  INV_X1    g099(.A(new_n249), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT102), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n298), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT103), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n295), .A2(KEYINPUT41), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT100), .ZN(new_n307));
  XOR2_X1   g106(.A(G134gat), .B(G162gat), .Z(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n304), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n305), .B1(new_n304), .B2(new_n309), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n303), .B1(new_n298), .B2(new_n302), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n304), .A2(new_n309), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT103), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n304), .A2(new_n305), .A3(new_n309), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n312), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n248), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT104), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n313), .B1(new_n310), .B2(new_n311), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(new_n312), .A3(new_n317), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT104), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n248), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G113gat), .B(G141gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT11), .ZN(new_n328));
  INV_X1    g127(.A(G169gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G197gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT12), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n299), .A2(new_n207), .ZN(new_n334));
  NAND2_X1  g133(.A1(G229gat), .A2(G233gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n206), .A2(new_n293), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n334), .A2(KEYINPUT18), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n206), .A2(new_n293), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT96), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT96), .B1(new_n206), .B2(new_n293), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(new_n338), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n335), .B(KEYINPUT13), .Z(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n336), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n346), .B1(new_n299), .B2(new_n207), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT18), .B1(new_n347), .B2(new_n335), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n333), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT18), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n352), .A2(new_n337), .A3(new_n344), .A4(new_n332), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G230gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n214), .A2(new_n215), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT98), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT98), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(new_n286), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT105), .B1(new_n282), .B2(new_n283), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n285), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n282), .A2(KEYINPUT105), .A3(new_n283), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n365), .A2(new_n214), .A3(new_n215), .A4(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n287), .B(KEYINPUT10), .C1(new_n216), .C2(new_n217), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n357), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G120gat), .B(G148gat), .Z(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(KEYINPUT108), .ZN(new_n372));
  XNOR2_X1  g171(.A(G176gat), .B(G204gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT106), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n362), .A2(new_n367), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(new_n357), .ZN(new_n378));
  AOI211_X1 g177(.A(KEYINPUT106), .B(new_n356), .C1(new_n362), .C2(new_n367), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(KEYINPUT107), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT107), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n375), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n356), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n374), .B(KEYINPUT109), .Z(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n326), .A2(new_n355), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT31), .B(G50gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(KEYINPUT89), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(KEYINPUT89), .ZN(new_n397));
  INV_X1    g196(.A(G228gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(new_n225), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G155gat), .B(G162gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G141gat), .B(G148gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(KEYINPUT2), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G155gat), .ZN(new_n405));
  INV_X1    g204(.A(G162gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT85), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(G162gat), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n405), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT2), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n401), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G141gat), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n413), .A2(KEYINPUT84), .A3(G148gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(G148gat), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT84), .B1(new_n413), .B2(G148gat), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n404), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(G211gat), .B(G218gat), .Z(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT79), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n423));
  INV_X1    g222(.A(G197gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(G204gat), .ZN(new_n425));
  INV_X1    g224(.A(G204gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(G197gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n423), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(G197gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n424), .A2(G204gat), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT78), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n422), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AOI211_X1 g234(.A(KEYINPUT79), .B(new_n433), .C1(new_n428), .C2(new_n431), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n421), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT78), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT78), .B1(new_n429), .B2(new_n430), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n434), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT79), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n432), .A2(new_n422), .A3(new_n434), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n420), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n437), .A2(new_n438), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT3), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n419), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n446), .B(new_n404), .C1(new_n412), .C2(new_n417), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n438), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT87), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(new_n451), .A3(new_n438), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n442), .A2(new_n420), .A3(new_n443), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n420), .B1(new_n442), .B2(new_n443), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT80), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT80), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(new_n437), .B2(new_n444), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n453), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n447), .B1(new_n459), .B2(KEYINPUT88), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT80), .B1(new_n454), .B2(new_n455), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n437), .A2(new_n457), .A3(new_n444), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n461), .A2(new_n462), .B1(new_n450), .B2(new_n452), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n400), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n446), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n418), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n456), .A2(new_n458), .ZN(new_n469));
  INV_X1    g268(.A(new_n449), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n468), .B(new_n400), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n466), .A2(G22gat), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G22gat), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n468), .B1(new_n463), .B2(new_n464), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n461), .A2(new_n462), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n476), .A2(new_n464), .A3(new_n453), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n399), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n474), .B1(new_n478), .B2(new_n471), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n396), .B(new_n397), .C1(new_n473), .C2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(G22gat), .B1(new_n466), .B2(new_n472), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n474), .A3(new_n471), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n481), .A2(KEYINPUT89), .A3(new_n482), .A4(new_n394), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT5), .ZN(new_n485));
  OR2_X1    g284(.A1(KEYINPUT73), .A2(G113gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(KEYINPUT73), .A2(G113gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(G120gat), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G113gat), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n489), .A2(G120gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT74), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n488), .A2(KEYINPUT74), .A3(new_n490), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(G127gat), .B(G134gat), .Z(new_n496));
  NOR2_X1   g295(.A1(new_n496), .A2(KEYINPUT1), .ZN(new_n497));
  XNOR2_X1  g296(.A(G113gat), .B(G120gat), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n498), .A2(KEYINPUT1), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n495), .A2(new_n497), .B1(new_n499), .B2(new_n496), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(KEYINPUT4), .A3(new_n419), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT4), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n488), .A2(KEYINPUT74), .A3(new_n490), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT74), .B1(new_n488), .B2(new_n490), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n497), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n499), .A2(new_n496), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n502), .B1(new_n507), .B2(new_n418), .ZN(new_n508));
  NAND2_X1  g307(.A1(G225gat), .A2(G233gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n418), .A2(KEYINPUT3), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n507), .A2(new_n510), .A3(new_n448), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n501), .A2(new_n508), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n509), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n500), .A2(new_n419), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n507), .A2(new_n418), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n485), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G1gat), .B(G29gat), .Z(new_n519));
  XNOR2_X1  g318(.A(G57gat), .B(G85gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n521), .B(new_n522), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n512), .A2(new_n485), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n523), .ZN(new_n526));
  INV_X1    g325(.A(new_n524), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(new_n517), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n518), .A2(KEYINPUT6), .A3(new_n523), .A4(new_n524), .ZN(new_n531));
  INV_X1    g330(.A(G183gat), .ZN(new_n532));
  OR2_X1    g331(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n533));
  NAND2_X1  g332(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n536));
  AOI21_X1  g335(.A(G190gat), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n534), .ZN(new_n538));
  NOR2_X1   g337(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n539));
  OAI21_X1  g338(.A(G183gat), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT69), .B1(new_n532), .B2(KEYINPUT27), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT28), .B1(new_n537), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G190gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT28), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT27), .B(G183gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT70), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n548), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G176gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n329), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(G169gat), .A2(G176gat), .ZN(new_n555));
  OAI22_X1  g354(.A1(new_n554), .A2(KEYINPUT71), .B1(new_n555), .B2(KEYINPUT26), .ZN(new_n556));
  NOR2_X1   g355(.A1(G169gat), .A2(G176gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT71), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT26), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G183gat), .A2(G190gat), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT72), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G169gat), .A2(G176gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n557), .A2(new_n558), .B1(new_n564), .B2(new_n559), .ZN(new_n565));
  NOR4_X1   g364(.A1(KEYINPUT71), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n566));
  OAI211_X1 g365(.A(KEYINPUT72), .B(new_n562), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI22_X1  g367(.A1(new_n544), .A2(new_n552), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT67), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(new_n557), .B2(KEYINPUT23), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT23), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n572), .B(KEYINPUT67), .C1(G169gat), .C2(G176gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n555), .B1(KEYINPUT23), .B2(new_n557), .ZN(new_n575));
  NOR2_X1   g374(.A1(G183gat), .A2(G190gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT24), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n574), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT25), .ZN(new_n583));
  AND2_X1   g382(.A1(G183gat), .A2(G190gat), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n576), .B1(new_n584), .B2(KEYINPUT24), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT66), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n562), .A2(KEYINPUT66), .A3(new_n578), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT25), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n589), .A2(new_n590), .A3(new_n574), .A4(new_n575), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n569), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G226gat), .A2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT81), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n596), .B(KEYINPUT82), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n536), .B(G183gat), .C1(new_n538), .C2(new_n539), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n601), .B(new_n545), .C1(new_n535), .C2(new_n541), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT28), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n546), .ZN(new_n605));
  INV_X1    g404(.A(new_n551), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n605), .B1(new_n606), .B2(new_n549), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT72), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n604), .A2(new_n607), .B1(new_n610), .B2(new_n567), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(new_n592), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n600), .B1(new_n612), .B2(KEYINPUT29), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n598), .B1(new_n613), .B2(KEYINPUT83), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n599), .B1(new_n594), .B2(new_n438), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT83), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n476), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G8gat), .B(G36gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G64gat), .B(G92gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n596), .B1(new_n612), .B2(KEYINPUT29), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n594), .A2(new_n599), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n469), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n618), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n530), .A2(new_n531), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n469), .A2(new_n624), .A3(new_n623), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n613), .A2(KEYINPUT83), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n616), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n598), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n629), .B1(new_n632), .B2(new_n476), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT37), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n622), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n469), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n634), .B1(new_n625), .B2(new_n476), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT38), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT38), .B1(new_n633), .B2(new_n634), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n618), .A2(new_n634), .A3(new_n626), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n621), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n628), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n501), .A2(new_n508), .A3(new_n511), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n513), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(KEYINPUT39), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n514), .A2(new_n515), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n646), .B(KEYINPUT39), .C1(new_n513), .C2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n649), .A3(new_n526), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n652), .A2(new_n525), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n615), .A2(new_n616), .B1(new_n594), .B2(new_n597), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n469), .B1(new_n654), .B2(new_n630), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n621), .B1(new_n655), .B2(new_n629), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(KEYINPUT30), .A3(new_n627), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT30), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n633), .A2(new_n658), .A3(new_n622), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n650), .A2(new_n651), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n653), .A2(new_n657), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n484), .A2(new_n644), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G227gat), .A2(G233gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT64), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT65), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n569), .A2(new_n593), .A3(new_n500), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n500), .B1(new_n569), .B2(new_n593), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n667), .B1(new_n668), .B2(KEYINPUT75), .ZN(new_n669));
  NOR4_X1   g468(.A1(new_n611), .A2(new_n507), .A3(new_n592), .A4(KEYINPUT75), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n666), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT32), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT76), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(G15gat), .B(G43gat), .Z(new_n675));
  XNOR2_X1  g474(.A(G71gat), .B(G99gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT76), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n507), .B1(new_n611), .B2(new_n592), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT75), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n670), .B1(new_n681), .B2(new_n667), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n678), .B(KEYINPUT32), .C1(new_n682), .C2(new_n666), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT33), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n682), .B2(new_n666), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n674), .A2(new_n677), .A3(new_n683), .A4(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n664), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n665), .A2(KEYINPUT34), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n688), .A2(KEYINPUT34), .B1(new_n682), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n669), .A2(new_n671), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n665), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT33), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(KEYINPUT32), .A3(new_n693), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n686), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n690), .B1(new_n686), .B2(new_n694), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT36), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT77), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(KEYINPUT77), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n697), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n683), .A2(new_n677), .A3(new_n685), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n678), .B1(new_n692), .B2(KEYINPUT32), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n694), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n690), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n686), .A2(new_n690), .A3(new_n694), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n700), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n657), .A2(new_n659), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n530), .A2(new_n531), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n480), .ZN(new_n714));
  INV_X1    g513(.A(new_n483), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n662), .A2(new_n702), .A3(new_n710), .A4(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n480), .A2(new_n707), .A3(new_n483), .A4(new_n708), .ZN(new_n718));
  OAI211_X1 g517(.A(KEYINPUT90), .B(KEYINPUT35), .C1(new_n718), .C2(new_n713), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT35), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n657), .A2(new_n659), .B1(new_n531), .B2(new_n530), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n484), .A2(new_n720), .A3(new_n697), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n697), .A2(new_n483), .A3(new_n480), .A4(new_n721), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT90), .B1(new_n724), .B2(KEYINPUT35), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n717), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n391), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n391), .A2(KEYINPUT110), .A3(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n712), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G1gat), .ZN(G1324gat));
  INV_X1    g533(.A(new_n711), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT16), .B(G8gat), .Z(new_n736));
  NAND3_X1  g535(.A1(new_n731), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n731), .A2(new_n735), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(G8gat), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n738), .B1(new_n737), .B2(new_n741), .ZN(G1325gat));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n709), .B1(new_n729), .B2(new_n730), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(G15gat), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n702), .A2(new_n710), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n731), .A2(G15gat), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n744), .A2(new_n743), .A3(G15gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(G1326gat));
  INV_X1    g550(.A(new_n484), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n731), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT43), .B(G22gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1327gat));
  INV_X1    g554(.A(new_n323), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n726), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n248), .A2(new_n355), .A3(new_n390), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n255), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(new_n732), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT45), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n726), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n717), .B(KEYINPUT112), .C1(new_n723), .C2(new_n725), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n321), .A2(new_n322), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n321), .B2(new_n322), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(KEYINPUT44), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n765), .A2(new_n766), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n757), .A2(KEYINPUT44), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n759), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n255), .B1(new_n776), .B2(new_n712), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n763), .A2(new_n777), .ZN(G1328gat));
  INV_X1    g577(.A(G36gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n760), .A2(new_n779), .A3(new_n735), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G36gat), .B1(new_n776), .B2(new_n711), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1329gat));
  NAND4_X1  g583(.A1(new_n775), .A2(G43gat), .A3(new_n747), .A4(new_n759), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n758), .A2(new_n697), .A3(new_n759), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n786), .A2(new_n260), .B1(KEYINPUT114), .B2(KEYINPUT47), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  OR2_X1    g587(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1330gat));
  INV_X1    g589(.A(KEYINPUT48), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n484), .A2(new_n258), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n760), .A2(new_n752), .ZN(new_n794));
  OAI221_X1 g593(.A(new_n791), .B1(new_n776), .B2(new_n793), .C1(new_n794), .C2(G50gat), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n776), .A2(new_n793), .ZN(new_n796));
  AOI21_X1  g595(.A(G50gat), .B1(new_n760), .B2(new_n752), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT48), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(G1331gat));
  AND2_X1   g598(.A1(new_n765), .A2(new_n766), .ZN(new_n800));
  INV_X1    g599(.A(new_n390), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n326), .A2(new_n354), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n732), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g605(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n807));
  AND2_X1   g606(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n808));
  NOR4_X1   g607(.A1(new_n803), .A2(new_n711), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n804), .A2(new_n735), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n807), .B2(new_n810), .ZN(G1333gat));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n800), .A2(new_n812), .A3(new_n697), .A4(new_n802), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n765), .A2(new_n697), .A3(new_n766), .A4(new_n802), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT115), .ZN(new_n815));
  AOI21_X1  g614(.A(G71gat), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n765), .A2(new_n747), .A3(new_n766), .A4(new_n802), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G71gat), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n816), .A2(KEYINPUT50), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n821));
  INV_X1    g620(.A(G71gat), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n814), .A2(KEYINPUT115), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n814), .A2(KEYINPUT115), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n821), .B1(new_n825), .B2(new_n818), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n820), .A2(new_n826), .ZN(G1334gat));
  NAND2_X1  g626(.A1(new_n804), .A2(new_n752), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g628(.A1(new_n248), .A2(new_n354), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n758), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n758), .A2(KEYINPUT51), .A3(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n835), .A2(new_n276), .A3(new_n732), .A4(new_n390), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n830), .A2(new_n390), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n773), .B2(new_n774), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(G85gat), .B1(new_n839), .B2(new_n712), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n836), .A2(new_n840), .ZN(G1336gat));
  OAI21_X1  g640(.A(G92gat), .B1(new_n839), .B2(new_n711), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n711), .A2(new_n801), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(G92gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n835), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n842), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n846), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n833), .B2(new_n834), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n277), .B1(new_n838), .B2(new_n735), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT52), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n852), .ZN(G1337gat));
  OAI21_X1  g652(.A(G99gat), .B1(new_n839), .B2(new_n746), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n709), .A2(new_n801), .A3(G99gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n835), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1338gat));
  OAI21_X1  g656(.A(G106gat), .B1(new_n839), .B2(new_n484), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n484), .A2(G106gat), .A3(new_n801), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n835), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n860), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n863), .B1(new_n833), .B2(new_n834), .ZN(new_n864));
  INV_X1    g663(.A(G106gat), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n865), .B1(new_n838), .B2(new_n752), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT53), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n862), .A2(new_n867), .ZN(G1339gat));
  NAND3_X1  g667(.A1(new_n368), .A2(new_n357), .A3(new_n369), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n386), .A2(KEYINPUT54), .A3(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n374), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n370), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT55), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n870), .A2(KEYINPUT55), .A3(new_n873), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n384), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n354), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880));
  INV_X1    g679(.A(new_n343), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n340), .B(new_n881), .C1(new_n341), .C2(new_n338), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT116), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n347), .A2(new_n335), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n331), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n353), .A3(new_n390), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n879), .A2(new_n880), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n880), .B1(new_n879), .B2(new_n886), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n769), .A2(new_n768), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n769), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n321), .A2(new_n322), .A3(new_n767), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n878), .A2(new_n353), .A3(new_n885), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n248), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  AND4_X1   g693(.A1(new_n320), .A2(new_n325), .A3(new_n355), .A4(new_n801), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n732), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n735), .ZN(new_n897));
  INV_X1    g696(.A(new_n718), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n898), .A3(new_n354), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G113gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n486), .A2(new_n487), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n899), .ZN(G1340gat));
  NAND3_X1  g701(.A1(new_n897), .A2(new_n898), .A3(new_n390), .ZN(new_n903));
  XNOR2_X1  g702(.A(KEYINPUT118), .B(G120gat), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n903), .B(new_n904), .ZN(G1341gat));
  NAND3_X1  g704(.A1(new_n897), .A2(new_n898), .A3(new_n248), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g706(.A1(new_n323), .A2(new_n735), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT119), .ZN(new_n909));
  NOR4_X1   g708(.A1(new_n896), .A2(G134gat), .A3(new_n718), .A4(new_n909), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT56), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n897), .A2(new_n898), .A3(new_n756), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G134gat), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1343gat));
  NOR2_X1   g713(.A1(new_n735), .A2(new_n712), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n746), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n752), .B1(new_n894), .B2(new_n895), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n355), .A2(new_n413), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n879), .A2(new_n886), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n323), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(KEYINPUT120), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n925), .B1(new_n323), .B2(new_n922), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n893), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n248), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n895), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n923), .B(KEYINPUT120), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n248), .B1(new_n932), .B2(new_n893), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT121), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n484), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n920), .B(new_n921), .C1(new_n935), .C2(new_n919), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n747), .A2(new_n484), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n897), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n413), .B1(new_n938), .B2(new_n355), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT58), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n936), .A2(new_n939), .A3(KEYINPUT58), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1344gat));
  OR3_X1    g743(.A1(new_n938), .A2(G148gat), .A3(new_n801), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G148gat), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n746), .B(new_n915), .C1(new_n917), .C2(KEYINPUT57), .ZN(new_n948));
  INV_X1    g747(.A(new_n895), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n949), .B1(new_n933), .B2(KEYINPUT121), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n929), .A2(new_n930), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n752), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n952), .B2(KEYINPUT57), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n947), .B1(new_n953), .B2(new_n390), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n756), .A2(new_n892), .ZN(new_n955));
  INV_X1    g754(.A(new_n923), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n928), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n949), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n919), .A3(new_n752), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n917), .A2(KEYINPUT57), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n916), .B(KEYINPUT122), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n959), .A2(new_n960), .A3(new_n390), .A4(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n946), .B1(new_n962), .B2(G148gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n945), .B1(new_n954), .B2(new_n963), .ZN(G1345gat));
  OAI21_X1  g763(.A(new_n920), .B1(new_n935), .B2(new_n919), .ZN(new_n965));
  OAI21_X1  g764(.A(G155gat), .B1(new_n965), .B2(new_n928), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n248), .A2(new_n405), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n938), .B2(new_n967), .ZN(G1346gat));
  AND2_X1   g767(.A1(new_n407), .A2(new_n409), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n965), .B2(new_n771), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n909), .A2(new_n970), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n937), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n971), .B1(new_n896), .B2(new_n973), .ZN(G1347gat));
  NAND2_X1  g773(.A1(new_n889), .A2(new_n893), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n928), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n732), .B1(new_n976), .B2(new_n949), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n718), .A2(new_n711), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(G169gat), .B1(new_n979), .B2(new_n354), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n711), .A2(new_n732), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(new_n697), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n484), .B1(new_n982), .B2(KEYINPUT123), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n983), .B1(KEYINPUT123), .B2(new_n982), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n984), .B1(new_n894), .B2(new_n895), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g786(.A(KEYINPUT124), .B(new_n984), .C1(new_n894), .C2(new_n895), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n355), .A2(new_n329), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n980), .B1(new_n989), .B2(new_n990), .ZN(G1348gat));
  NAND2_X1  g790(.A1(new_n977), .A2(new_n978), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n553), .B1(new_n992), .B2(new_n801), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n993), .A2(KEYINPUT125), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(KEYINPUT125), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n989), .A2(G176gat), .A3(new_n390), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(G1349gat));
  OAI211_X1 g796(.A(new_n979), .B(new_n248), .C1(new_n606), .C2(new_n549), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n987), .A2(new_n248), .A3(new_n988), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(G183gat), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(KEYINPUT60), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT60), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n998), .A2(new_n1003), .A3(new_n1000), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1002), .A2(new_n1004), .ZN(G1350gat));
  INV_X1    g804(.A(KEYINPUT61), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n987), .A2(new_n756), .A3(new_n988), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n1008));
  AND3_X1   g807(.A1(new_n1007), .A2(new_n1008), .A3(G190gat), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1008), .B1(new_n1007), .B2(G190gat), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1006), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1007), .A2(G190gat), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(KEYINPUT126), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1007), .A2(new_n1008), .A3(G190gat), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1013), .A2(KEYINPUT61), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n979), .A2(new_n545), .A3(new_n770), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1011), .A2(new_n1015), .A3(new_n1016), .ZN(G1351gat));
  NAND2_X1  g816(.A1(new_n977), .A2(new_n937), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n1018), .A2(new_n711), .ZN(new_n1019));
  AOI21_X1  g818(.A(G197gat), .B1(new_n1019), .B2(new_n354), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n746), .A2(new_n981), .ZN(new_n1021));
  INV_X1    g820(.A(new_n1021), .ZN(new_n1022));
  AND3_X1   g821(.A1(new_n959), .A2(new_n960), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n355), .A2(new_n424), .ZN(new_n1024));
  AOI21_X1  g823(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(G1352gat));
  NOR3_X1   g824(.A1(new_n1018), .A2(G204gat), .A3(new_n845), .ZN(new_n1026));
  XNOR2_X1  g825(.A(new_n1026), .B(KEYINPUT62), .ZN(new_n1027));
  NAND3_X1  g826(.A1(new_n959), .A2(new_n960), .A3(new_n390), .ZN(new_n1028));
  OAI21_X1  g827(.A(G204gat), .B1(new_n1028), .B2(new_n1021), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1027), .A2(new_n1029), .ZN(G1353gat));
  INV_X1    g829(.A(G211gat), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n1019), .A2(new_n1031), .A3(new_n248), .ZN(new_n1032));
  NAND4_X1  g831(.A1(new_n959), .A2(new_n960), .A3(new_n248), .A4(new_n1022), .ZN(new_n1033));
  AND3_X1   g832(.A1(new_n1033), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1034));
  AOI21_X1  g833(.A(KEYINPUT63), .B1(new_n1033), .B2(G211gat), .ZN(new_n1035));
  OAI21_X1  g834(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(G1354gat));
  AOI21_X1  g835(.A(G218gat), .B1(new_n1019), .B2(new_n770), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n756), .A2(G218gat), .ZN(new_n1038));
  XOR2_X1   g837(.A(new_n1038), .B(KEYINPUT127), .Z(new_n1039));
  AOI21_X1  g838(.A(new_n1037), .B1(new_n1023), .B2(new_n1039), .ZN(G1355gat));
endmodule


