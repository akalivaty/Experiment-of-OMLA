//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT77), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT75), .B1(new_n191), .B2(G107), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(G107), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n191), .A2(KEYINPUT75), .A3(G107), .ZN(new_n195));
  OAI21_X1  g009(.A(G101), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT2), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G113), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G116), .B(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n204), .A2(new_n207), .A3(new_n208), .A4(new_n193), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n196), .A2(new_n203), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT5), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  INV_X1    g026(.A(G116), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G119), .ZN(new_n214));
  INV_X1    g028(.A(G119), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G116), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(G116), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(G119), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT66), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n211), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n197), .B1(new_n214), .B2(new_n211), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT76), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT66), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n218), .B2(new_n219), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT5), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(new_n222), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n210), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n217), .A2(new_n198), .A3(new_n200), .A4(new_n220), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n203), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n204), .A2(new_n207), .A3(new_n193), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G101), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT4), .A3(new_n209), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n236), .A3(G101), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n232), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n190), .B1(new_n230), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n210), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n221), .A2(KEYINPUT76), .A3(new_n223), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n228), .B1(new_n227), .B2(new_n222), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n232), .A2(new_n235), .A3(new_n237), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(new_n189), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n239), .A2(new_n245), .A3(KEYINPUT6), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT1), .B1(new_n247), .B2(G146), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(G146), .ZN(new_n249));
  INV_X1    g063(.A(G146), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  OAI211_X1 g065(.A(G128), .B(new_n248), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT74), .B(G125), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n247), .A2(G146), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n254), .B(new_n255), .C1(KEYINPUT1), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n252), .A2(new_n253), .A3(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT0), .A4(G128), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT74), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT74), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G125), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n249), .A2(new_n251), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G128), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n259), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G224), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(G953), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n268), .B(new_n271), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n273));
  OAI211_X1 g087(.A(new_n190), .B(new_n273), .C1(new_n230), .C2(new_n238), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n246), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT79), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT79), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n246), .A2(new_n277), .A3(new_n272), .A4(new_n274), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  INV_X1    g094(.A(new_n268), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n271), .A2(KEYINPUT7), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT82), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n281), .B(new_n282), .C1(new_n283), .C2(new_n270), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT7), .B(new_n271), .C1(new_n268), .C2(KEYINPUT82), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT81), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT5), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n222), .A2(new_n288), .B1(new_n201), .B2(new_n202), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT80), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n209), .B(new_n196), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n222), .A2(new_n288), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n292), .A2(new_n290), .A3(new_n203), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n287), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OR2_X1    g108(.A1(new_n289), .A2(new_n290), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n196), .A2(new_n209), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n289), .A2(new_n290), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n295), .A2(new_n297), .A3(KEYINPUT81), .A4(new_n298), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n224), .A2(new_n229), .B1(new_n201), .B2(new_n202), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n294), .B(new_n299), .C1(new_n300), .C2(new_n297), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n189), .B(KEYINPUT8), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n286), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n245), .B1(new_n303), .B2(KEYINPUT83), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n305));
  AOI211_X1 g119(.A(new_n305), .B(new_n286), .C1(new_n301), .C2(new_n302), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n280), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n188), .B1(new_n279), .B2(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n301), .A2(new_n302), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n305), .B1(new_n309), .B2(new_n286), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n303), .A2(KEYINPUT83), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n245), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n276), .A2(new_n278), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n280), .A4(new_n187), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G478), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT15), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(KEYINPUT94), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n318), .B1(KEYINPUT94), .B2(new_n317), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT9), .B(G234), .ZN(new_n320));
  INV_X1    g134(.A(G217), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n320), .A2(new_n321), .A3(G953), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(G116), .B(G122), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(new_n206), .ZN(new_n325));
  XNOR2_X1  g139(.A(G128), .B(G143), .ZN(new_n326));
  INV_X1    g140(.A(G134), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT93), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n326), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n256), .A2(G143), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n327), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n330), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n335), .A3(new_n330), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n329), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n326), .B(new_n327), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n213), .A2(KEYINPUT14), .A3(G122), .ZN(new_n341));
  INV_X1    g155(.A(new_n324), .ZN(new_n342));
  OAI211_X1 g156(.A(G107), .B(new_n341), .C1(new_n342), .C2(KEYINPUT14), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n324), .A2(new_n206), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n323), .B1(new_n339), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n338), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(new_n336), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n345), .B(new_n322), .C1(new_n349), .C2(new_n329), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT70), .B(G902), .Z(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT95), .ZN(new_n354));
  INV_X1    g168(.A(new_n352), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(new_n347), .B2(new_n350), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT95), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n319), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n356), .A2(new_n357), .ZN(new_n360));
  INV_X1    g174(.A(new_n319), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n364));
  INV_X1    g178(.A(G237), .ZN(new_n365));
  INV_X1    g179(.A(G953), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(G214), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n247), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n365), .A2(new_n366), .A3(G143), .A4(G214), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G131), .ZN(new_n371));
  INV_X1    g185(.A(G131), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n372), .A3(new_n369), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n364), .B1(new_n374), .B2(KEYINPUT17), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT17), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n371), .A2(KEYINPUT88), .A3(new_n376), .A4(new_n373), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n370), .A2(KEYINPUT17), .A3(G131), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n261), .A2(new_n263), .A3(G140), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n260), .A2(G140), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(KEYINPUT16), .A2(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n264), .A2(new_n385), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n384), .A2(G146), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(G146), .B1(new_n384), .B2(new_n386), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n380), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n384), .A2(new_n386), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n250), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n384), .A2(G146), .A3(new_n386), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT87), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n370), .ZN(new_n395));
  NAND2_X1  g209(.A1(KEYINPUT18), .A2(G131), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT84), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n260), .A2(G140), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n383), .A2(new_n401), .A3(new_n250), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n382), .B1(new_n253), .B2(G140), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n250), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n404), .B1(new_n395), .B2(new_n396), .ZN(new_n405));
  OAI22_X1  g219(.A1(new_n379), .A2(new_n394), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G113), .B(G122), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(new_n191), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT19), .B1(new_n383), .B2(new_n401), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n403), .B2(KEYINPUT19), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n392), .B1(new_n411), .B2(G146), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT86), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT86), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n414), .B(new_n392), .C1(new_n411), .C2(G146), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n374), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n408), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n416), .B(new_n417), .C1(new_n400), .C2(new_n405), .ZN(new_n418));
  NOR2_X1   g232(.A1(G475), .A2(G902), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n419), .A2(KEYINPUT89), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(KEYINPUT89), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT20), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n409), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n409), .A2(new_n418), .A3(new_n419), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT20), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n409), .A2(new_n418), .A3(KEYINPUT90), .A4(new_n422), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G952), .ZN(new_n430));
  AOI211_X1 g244(.A(G953), .B(new_n430), .C1(G234), .C2(G237), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n366), .B(new_n352), .C1(G234), .C2(G237), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  XOR2_X1   g248(.A(KEYINPUT21), .B(G898), .Z(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT96), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n432), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n417), .A2(KEYINPUT91), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n406), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n406), .A2(new_n439), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n280), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n438), .B1(new_n442), .B2(G475), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n363), .A2(new_n429), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G214), .B1(G237), .B2(G902), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n315), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G110), .B(G140), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n366), .A2(G227), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n447), .B(new_n448), .Z(new_n449));
  NAND2_X1  g263(.A1(new_n252), .A2(new_n257), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n296), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT10), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n259), .B1(new_n265), .B2(new_n266), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n235), .A2(new_n454), .A3(new_n237), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT10), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n296), .B2(new_n450), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n452), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G137), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT11), .A3(G134), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n327), .A2(G137), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT11), .ZN(new_n463));
  OAI211_X1 g277(.A(KEYINPUT64), .B(new_n463), .C1(new_n327), .C2(G137), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n459), .A2(G134), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT64), .B1(new_n466), .B2(new_n463), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n462), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G131), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n462), .B(new_n372), .C1(new_n465), .C2(new_n467), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT67), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT67), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n458), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n458), .A2(new_n475), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n449), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n469), .A2(KEYINPUT67), .A3(new_n470), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT67), .B1(new_n469), .B2(new_n470), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n481), .A2(new_n455), .A3(new_n457), .A4(new_n452), .ZN(new_n482));
  INV_X1    g296(.A(new_n449), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n252), .A2(new_n257), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n209), .B2(new_n196), .ZN(new_n486));
  OAI221_X1 g300(.A(new_n484), .B1(new_n486), .B2(new_n451), .C1(new_n479), .C2(new_n480), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n471), .B1(new_n486), .B2(new_n451), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT12), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n482), .A2(new_n483), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n478), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G469), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n492), .A3(new_n352), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n280), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n487), .A2(new_n489), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n449), .B1(new_n496), .B2(new_n477), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n458), .A2(new_n475), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n482), .A2(new_n498), .A3(new_n483), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(G469), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n493), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G221), .B1(new_n320), .B2(G902), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n446), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n321), .B1(new_n352), .B2(G234), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n256), .B(G119), .C1(KEYINPUT72), .C2(KEYINPUT23), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT23), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(new_n215), .B2(G128), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT72), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n215), .B2(G128), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n513), .A2(G110), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  XOR2_X1   g329(.A(KEYINPUT24), .B(G110), .Z(new_n516));
  NOR2_X1   g330(.A1(new_n256), .A2(G119), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n215), .A2(G128), .ZN(new_n518));
  OR3_X1    g332(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT71), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT71), .B1(new_n517), .B2(new_n518), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n392), .B(new_n402), .C1(new_n515), .C2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n387), .A2(new_n388), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n519), .A2(new_n520), .A3(new_n516), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n513), .A2(new_n525), .A3(G110), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n525), .B1(new_n513), .B2(G110), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n522), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT22), .B(G137), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n366), .A2(G221), .A3(G234), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n522), .B(new_n532), .C1(new_n523), .C2(new_n528), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n352), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT25), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n537), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n507), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n534), .A2(new_n535), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n542), .A2(G902), .A3(new_n506), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n454), .B1(new_n479), .B2(new_n480), .ZN(new_n545));
  INV_X1    g359(.A(new_n232), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n466), .A2(new_n461), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G131), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n485), .A2(new_n470), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT28), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT68), .ZN(new_n553));
  INV_X1    g367(.A(new_n470), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n252), .A2(new_n548), .A3(new_n257), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n485), .A2(new_n470), .A3(KEYINPUT68), .A4(new_n548), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n545), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(new_n546), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n552), .B1(new_n560), .B2(KEYINPUT28), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n365), .A2(new_n366), .A3(G210), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n562), .B(KEYINPUT27), .Z(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT26), .B(G101), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n563), .B(new_n564), .Z(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT29), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n355), .B1(new_n561), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n545), .A2(new_n558), .A3(KEYINPUT30), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT30), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n453), .B1(new_n469), .B2(new_n470), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n549), .B1(new_n572), .B2(KEYINPUT65), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT65), .ZN(new_n574));
  AOI211_X1 g388(.A(new_n574), .B(new_n453), .C1(new_n469), .C2(new_n470), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n571), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n570), .A2(new_n576), .A3(new_n232), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT69), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n570), .A2(new_n576), .A3(KEYINPUT69), .A4(new_n232), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n545), .A2(new_n546), .A3(new_n558), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(new_n565), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT28), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n232), .B1(new_n573), .B2(new_n575), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n587), .A2(new_n552), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n567), .B1(new_n588), .B2(new_n566), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n569), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G472), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n566), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n582), .A2(new_n565), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT31), .B1(new_n581), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT31), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n596), .B(new_n593), .C1(new_n579), .C2(new_n580), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n592), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT32), .ZN(new_n599));
  NOR2_X1   g413(.A1(G472), .A2(G902), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n599), .B1(new_n598), .B2(new_n600), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n591), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n505), .A2(new_n544), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  AND2_X1   g420(.A1(new_n588), .A2(new_n566), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n581), .A2(new_n594), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n596), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n581), .A2(new_n594), .A3(KEYINPUT31), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G472), .B1(new_n611), .B2(new_n355), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n598), .A2(new_n600), .ZN(new_n613));
  INV_X1    g427(.A(new_n544), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n503), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n612), .A2(KEYINPUT97), .A3(new_n615), .A4(new_n613), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n356), .B2(G478), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n353), .A2(KEYINPUT100), .A3(new_n316), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n624));
  AND3_X1   g438(.A1(new_n347), .A2(new_n350), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n347), .A2(new_n350), .B1(new_n626), .B2(KEYINPUT33), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n355), .A2(new_n316), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n622), .A2(new_n623), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n442), .A2(G475), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n438), .B(new_n630), .C1(new_n429), .C2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n308), .A2(new_n633), .A3(new_n314), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n279), .A2(new_n307), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(KEYINPUT98), .A3(new_n187), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n632), .A2(new_n634), .A3(new_n445), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT101), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n620), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT34), .B(G104), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NOR2_X1   g455(.A1(new_n314), .A2(new_n633), .ZN(new_n642));
  INV_X1    g456(.A(new_n445), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT20), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n409), .A2(new_n418), .A3(new_n645), .A4(new_n419), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n427), .A2(new_n646), .A3(KEYINPUT102), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n426), .A2(new_n648), .A3(KEYINPUT20), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n443), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n650), .A2(new_n651), .A3(new_n363), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n644), .A2(new_n634), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n618), .A2(new_n619), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  INV_X1    g470(.A(new_n540), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n506), .B1(new_n657), .B2(new_n538), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT103), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n529), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n280), .A3(new_n507), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n501), .A3(new_n502), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n446), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n612), .A2(new_n613), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT104), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT37), .B(G110), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  INV_X1    g485(.A(new_n600), .ZN(new_n672));
  OAI21_X1  g486(.A(KEYINPUT32), .B1(new_n611), .B2(new_n672), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n673), .A2(new_n601), .B1(G472), .B2(new_n590), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n644), .A2(new_n634), .A3(new_n665), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n432), .B1(new_n434), .B2(G900), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n647), .A2(new_n649), .A3(new_n631), .A4(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n363), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  XNOR2_X1  g495(.A(new_n677), .B(KEYINPUT39), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n503), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n363), .B1(new_n429), .B2(new_n631), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n658), .A2(new_n662), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n445), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n673), .A2(new_n601), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n583), .A2(new_n566), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n280), .B1(new_n560), .B2(new_n565), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n315), .B(KEYINPUT38), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n685), .A2(new_n686), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n691), .A2(new_n696), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G143), .ZN(G45));
  AOI21_X1  g514(.A(new_n630), .B1(new_n429), .B2(new_n631), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(new_n677), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n676), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n637), .B(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n614), .B1(new_n692), .B2(new_n591), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n355), .B1(new_n478), .B2(new_n490), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n492), .ZN(new_n709));
  AOI211_X1 g523(.A(G469), .B(new_n355), .C1(new_n478), .C2(new_n490), .ZN(new_n710));
  INV_X1    g524(.A(new_n502), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(KEYINPUT106), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(KEYINPUT106), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n706), .A2(new_n707), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND4_X1  g532(.A1(new_n604), .A2(new_n653), .A3(new_n544), .A4(new_n715), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  NAND2_X1  g534(.A1(new_n444), .A2(new_n663), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n692), .B2(new_n591), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n634), .A2(new_n636), .A3(new_n445), .A4(new_n712), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n644), .A2(KEYINPUT107), .A3(new_n634), .A4(new_n712), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n722), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n723), .B1(new_n722), .B2(new_n728), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT109), .B(G119), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G21));
  NAND2_X1  g547(.A1(new_n612), .A2(KEYINPUT110), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n735), .B(G472), .C1(new_n611), .C2(new_n355), .ZN(new_n736));
  OAI22_X1  g550(.A1(new_n595), .A2(new_n597), .B1(new_n561), .B2(new_n565), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n734), .A2(new_n736), .B1(new_n600), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n713), .A2(new_n714), .A3(new_n437), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n634), .A2(new_n636), .A3(new_n445), .A4(new_n688), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(new_n544), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NAND4_X1  g557(.A1(new_n738), .A2(new_n663), .A3(new_n728), .A4(new_n702), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  NAND3_X1  g559(.A1(new_n308), .A2(new_n445), .A3(new_n314), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n308), .A2(KEYINPUT113), .A3(new_n445), .A4(new_n314), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n499), .A2(KEYINPUT112), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n482), .A2(new_n498), .A3(new_n751), .A4(new_n483), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n497), .A2(KEYINPUT111), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(new_n449), .C1(new_n496), .C2(new_n477), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n753), .A2(new_n754), .A3(G469), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n494), .B1(new_n708), .B2(new_n492), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n711), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n748), .A2(new_n702), .A3(new_n749), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT42), .B1(new_n707), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n674), .A2(new_n760), .A3(new_n763), .A4(new_n614), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n372), .ZN(G33));
  AND4_X1   g580(.A1(new_n679), .A2(new_n748), .A3(new_n749), .A4(new_n759), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n707), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  AND2_X1   g583(.A1(new_n429), .A2(new_n631), .ZN(new_n770));
  INV_X1    g584(.A(new_n630), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(KEYINPUT43), .Z(new_n773));
  AND3_X1   g587(.A1(new_n773), .A2(new_n667), .A3(new_n663), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT44), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n753), .A2(new_n754), .A3(KEYINPUT45), .A4(new_n756), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n497), .A2(new_n499), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n776), .B(G469), .C1(KEYINPUT45), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n495), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(KEYINPUT46), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n493), .B1(new_n780), .B2(KEYINPUT46), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n502), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(new_n683), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n748), .A2(new_n749), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n774), .A2(KEYINPUT44), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n775), .A2(new_n785), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  XNOR2_X1  g604(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n783), .B(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n674), .A2(new_n787), .A3(new_n614), .A4(new_n702), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  NAND3_X1  g609(.A1(new_n544), .A2(new_n445), .A3(new_n502), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT115), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n772), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT116), .Z(new_n799));
  NOR2_X1   g613(.A1(new_n709), .A2(new_n710), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT49), .Z(new_n801));
  OR4_X1    g615(.A1(new_n696), .A2(new_n799), .A3(new_n697), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n712), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n432), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n773), .A2(new_n787), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n805), .A2(new_n614), .A3(new_n674), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT48), .Z(new_n807));
  NAND2_X1  g621(.A1(new_n738), .A2(new_n544), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n773), .A2(new_n431), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n728), .ZN(new_n811));
  INV_X1    g625(.A(new_n696), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n544), .A2(new_n812), .A3(new_n787), .A4(new_n804), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n430), .B(G953), .C1(new_n813), .C2(new_n701), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n807), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n738), .A2(new_n663), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n805), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n697), .A2(new_n445), .A3(new_n803), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n810), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT50), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n770), .A2(new_n630), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n817), .B(new_n820), .C1(new_n813), .C2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n808), .A2(new_n809), .A3(new_n786), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n792), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n800), .A2(new_n711), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n792), .B2(new_n825), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n824), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT51), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n792), .A2(new_n827), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n831), .B1(new_n832), .B2(new_n824), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n815), .B(new_n830), .C1(new_n823), .C2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n315), .A2(new_n445), .A3(new_n437), .ZN(new_n836));
  INV_X1    g650(.A(new_n358), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n361), .B1(new_n837), .B2(new_n360), .ZN(new_n838));
  INV_X1    g652(.A(new_n362), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT117), .B1(new_n359), .B2(new_n362), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n701), .B1(new_n770), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n836), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n618), .A2(new_n845), .A3(new_n619), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n742), .A2(new_n846), .A3(new_n719), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n666), .A2(new_n667), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n604), .A2(new_n544), .A3(new_n715), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n605), .B(new_n848), .C1(new_n638), .C2(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n731), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n744), .A2(new_n680), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n759), .A2(new_n689), .A3(new_n677), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n740), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n676), .A2(new_n702), .B1(new_n858), .B2(new_n696), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n852), .A2(new_n853), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n680), .A3(new_n744), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT52), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n748), .A2(new_n749), .A3(new_n759), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n738), .A2(new_n663), .A3(new_n702), .A4(new_n863), .ZN(new_n864));
  OR3_X1    g678(.A1(new_n664), .A2(new_n843), .A3(new_n678), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n786), .A2(new_n865), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n707), .A2(new_n767), .B1(new_n866), .B2(new_n604), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n864), .B(new_n867), .C1(new_n762), .C2(new_n764), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n851), .A2(new_n860), .A3(new_n862), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n668), .B1(new_n707), .B2(new_n505), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n873), .B(new_n716), .C1(new_n729), .C2(new_n730), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n874), .A2(new_n868), .A3(new_n847), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(KEYINPUT53), .A3(new_n860), .A4(new_n862), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n835), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n872), .A2(new_n878), .A3(new_n876), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n870), .A2(KEYINPUT119), .A3(new_n871), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT54), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n834), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n802), .B1(new_n883), .B2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n366), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n879), .A2(new_n880), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n352), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT56), .B1(new_n889), .B2(new_n188), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n246), .A2(new_n274), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT121), .Z(new_n892));
  XOR2_X1   g706(.A(new_n272), .B(KEYINPUT55), .Z(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n887), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n890), .B2(new_n894), .ZN(G51));
  XNOR2_X1  g710(.A(new_n494), .B(KEYINPUT57), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n879), .A2(KEYINPUT54), .A3(new_n880), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n899), .B2(new_n881), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n491), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n901), .A2(KEYINPUT122), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n778), .B(KEYINPUT123), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n901), .A2(KEYINPUT122), .B1(new_n889), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n886), .B1(new_n902), .B2(new_n904), .ZN(G54));
  NAND3_X1  g719(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n409), .A2(new_n418), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n886), .ZN(G60));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n911));
  INV_X1    g725(.A(new_n628), .ZN(new_n912));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT59), .Z(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n888), .A2(new_n835), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(new_n898), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n911), .B1(new_n918), .B2(new_n886), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n915), .B1(new_n899), .B2(new_n881), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(KEYINPUT124), .A3(new_n887), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n912), .B1(new_n882), .B2(new_n914), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n919), .A2(new_n921), .A3(new_n925), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(G63));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT60), .Z(new_n929));
  NAND3_X1  g743(.A1(new_n879), .A2(new_n880), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n886), .B1(new_n930), .B2(new_n542), .ZN(new_n931));
  INV_X1    g745(.A(new_n661), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n930), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g748(.A(new_n366), .B1(new_n436), .B2(G224), .ZN(new_n935));
  INV_X1    g749(.A(new_n851), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n366), .ZN(new_n937));
  INV_X1    g751(.A(G898), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n892), .B1(new_n938), .B2(G953), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n937), .B(new_n939), .ZN(G69));
  AOI21_X1  g754(.A(new_n366), .B1(G227), .B2(G900), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n784), .A2(new_n740), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n707), .B1(new_n942), .B2(new_n767), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n794), .A3(new_n789), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n852), .A2(new_n703), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n765), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n366), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n570), .A2(new_n576), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(new_n411), .ZN(new_n949));
  NAND2_X1  g763(.A1(G900), .A2(G953), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n941), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n786), .A2(new_n685), .A3(new_n844), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n707), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n794), .A2(new_n789), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n852), .A2(new_n699), .A3(new_n703), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(KEYINPUT62), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n959));
  AOI21_X1  g773(.A(G953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n951), .B1(new_n960), .B2(new_n949), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n953), .B(new_n961), .Z(G72));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n608), .B1(new_n584), .B2(new_n965), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n583), .A2(KEYINPUT127), .A3(new_n565), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n872), .B2(new_n876), .ZN(new_n969));
  INV_X1    g783(.A(new_n964), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n946), .B2(new_n851), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n583), .A2(new_n566), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n887), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n958), .A2(new_n851), .A3(new_n959), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n964), .ZN(new_n975));
  AOI211_X1 g789(.A(new_n969), .B(new_n973), .C1(new_n693), .C2(new_n975), .ZN(G57));
endmodule


