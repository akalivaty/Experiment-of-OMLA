

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n620, n621, n622, n623, n624,
         n625, n626, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788;

  INV_X1 U380 ( .A(KEYINPUT41), .ZN(n360) );
  XNOR2_X1 U381 ( .A(G137), .B(G140), .ZN(n515) );
  INV_X1 U382 ( .A(G237), .ZN(n450) );
  XNOR2_X1 U383 ( .A(G101), .B(G107), .ZN(n488) );
  XNOR2_X1 U384 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n460) );
  INV_X1 U385 ( .A(G107), .ZN(n442) );
  XNOR2_X2 U386 ( .A(n394), .B(n395), .ZN(n597) );
  NAND2_X4 U387 ( .A1(n652), .A2(G953), .ZN(n722) );
  XNOR2_X2 U388 ( .A(n617), .B(n616), .ZN(n689) );
  XNOR2_X2 U389 ( .A(n359), .B(n626), .ZN(n635) );
  NAND2_X1 U390 ( .A1(n624), .A2(n625), .ZN(n359) );
  XNOR2_X2 U391 ( .A(n540), .B(KEYINPUT6), .ZN(n607) );
  AND2_X2 U392 ( .A1(n543), .A2(n748), .ZN(n552) );
  XNOR2_X2 U393 ( .A(n361), .B(n360), .ZN(n779) );
  NOR2_X4 U394 ( .A1(n767), .A2(n618), .ZN(n361) );
  XOR2_X2 U395 ( .A(n711), .B(KEYINPUT59), .Z(n712) );
  XOR2_X2 U396 ( .A(KEYINPUT62), .B(n695), .Z(n696) );
  XNOR2_X2 U397 ( .A(n648), .B(n649), .ZN(n650) );
  XNOR2_X2 U398 ( .A(n449), .B(G902), .ZN(n637) );
  XNOR2_X2 U399 ( .A(KEYINPUT67), .B(KEYINPUT22), .ZN(n482) );
  NAND2_X2 U400 ( .A1(n362), .A2(n441), .ZN(n483) );
  XNOR2_X2 U401 ( .A(n396), .B(n393), .ZN(n362) );
  XNOR2_X1 U402 ( .A(G116), .B(KEYINPUT5), .ZN(n500) );
  NAND2_X1 U403 ( .A1(G234), .A2(G237), .ZN(n452) );
  INV_X1 U404 ( .A(KEYINPUT15), .ZN(n449) );
  AND2_X1 U405 ( .A1(n555), .A2(n554), .ZN(n765) );
  INV_X1 U406 ( .A(G902), .ZN(n400) );
  XNOR2_X2 U407 ( .A(n409), .B(KEYINPUT80), .ZN(n731) );
  NOR2_X2 U408 ( .A1(n621), .A2(n583), .ZN(n409) );
  NAND2_X2 U409 ( .A1(n581), .A2(n458), .ZN(n396) );
  XNOR2_X2 U410 ( .A(n397), .B(n410), .ZN(n581) );
  XOR2_X1 U411 ( .A(G131), .B(G140), .Z(n490) );
  BUF_X2 U412 ( .A(G128), .Z(n657) );
  NOR2_X2 U413 ( .A1(G953), .A2(G237), .ZN(n499) );
  NOR2_X1 U414 ( .A1(n381), .A2(n382), .ZN(n602) );
  NAND2_X1 U415 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U416 ( .A1(n433), .A2(KEYINPUT36), .ZN(n432) );
  XNOR2_X1 U417 ( .A(KEYINPUT42), .B(n388), .ZN(n787) );
  XNOR2_X1 U418 ( .A(n407), .B(n406), .ZN(n557) );
  AND2_X1 U419 ( .A1(n779), .A2(n622), .ZN(n388) );
  XNOR2_X1 U420 ( .A(n609), .B(KEYINPUT111), .ZN(n433) );
  OR2_X1 U421 ( .A1(n620), .A2(n582), .ZN(n583) );
  XNOR2_X1 U422 ( .A(n530), .B(n363), .ZN(n611) );
  XNOR2_X1 U423 ( .A(n630), .B(KEYINPUT38), .ZN(n763) );
  XNOR2_X1 U424 ( .A(n471), .B(n470), .ZN(n555) );
  XNOR2_X1 U425 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U426 ( .A(n423), .B(n374), .ZN(n534) );
  XNOR2_X1 U427 ( .A(n460), .B(n459), .ZN(n512) );
  XOR2_X2 U428 ( .A(KEYINPUT70), .B(KEYINPUT97), .Z(n489) );
  XNOR2_X2 U429 ( .A(G113), .B(G143), .ZN(n421) );
  XNOR2_X2 U430 ( .A(G137), .B(G134), .ZN(n484) );
  XNOR2_X2 U431 ( .A(G110), .B(G119), .ZN(n509) );
  XNOR2_X1 U432 ( .A(KEYINPUT1), .B(KEYINPUT92), .ZN(n363) );
  XNOR2_X1 U433 ( .A(KEYINPUT86), .B(KEYINPUT45), .ZN(n570) );
  XNOR2_X1 U434 ( .A(n364), .B(KEYINPUT82), .ZN(n639) );
  NAND2_X1 U435 ( .A1(n365), .A2(n679), .ZN(n364) );
  XNOR2_X2 U436 ( .A(n741), .B(n636), .ZN(n679) );
  NOR2_X4 U437 ( .A1(n635), .A2(n634), .ZN(n741) );
  XNOR2_X1 U438 ( .A(n366), .B(KEYINPUT83), .ZN(n365) );
  NAND2_X1 U439 ( .A1(n642), .A2(n637), .ZN(n366) );
  XNOR2_X2 U440 ( .A(n368), .B(n367), .ZN(n663) );
  XNOR2_X2 U441 ( .A(n494), .B(KEYINPUT16), .ZN(n367) );
  XNOR2_X2 U442 ( .A(n372), .B(G110), .ZN(n494) );
  XNOR2_X2 U443 ( .A(n505), .B(n465), .ZN(n368) );
  XNOR2_X2 U444 ( .A(n371), .B(n442), .ZN(n465) );
  XNOR2_X2 U445 ( .A(n370), .B(n369), .ZN(n505) );
  XNOR2_X2 U446 ( .A(G119), .B(KEYINPUT3), .ZN(n369) );
  XNOR2_X2 U447 ( .A(G113), .B(G101), .ZN(n370) );
  XNOR2_X2 U448 ( .A(G122), .B(G116), .ZN(n371) );
  XNOR2_X2 U449 ( .A(G104), .B(KEYINPUT94), .ZN(n372) );
  XNOR2_X1 U450 ( .A(n396), .B(n393), .ZN(n373) );
  NOR2_X2 U451 ( .A1(n390), .A2(n526), .ZN(n527) );
  BUF_X2 U452 ( .A(n597), .Z(n630) );
  XNOR2_X1 U453 ( .A(n422), .B(n421), .ZN(n420) );
  XNOR2_X1 U454 ( .A(G122), .B(G104), .ZN(n422) );
  XNOR2_X1 U455 ( .A(n418), .B(KEYINPUT11), .ZN(n417) );
  INV_X1 U456 ( .A(KEYINPUT12), .ZN(n418) );
  XNOR2_X1 U457 ( .A(KEYINPUT103), .B(KEYINPUT102), .ZN(n416) );
  INV_X1 U458 ( .A(KEYINPUT0), .ZN(n393) );
  INV_X1 U459 ( .A(n497), .ZN(n401) );
  XNOR2_X1 U460 ( .A(G131), .B(KEYINPUT100), .ZN(n502) );
  INV_X1 U461 ( .A(n745), .ZN(n645) );
  INV_X1 U462 ( .A(KEYINPUT65), .ZN(n640) );
  INV_X1 U463 ( .A(KEYINPUT107), .ZN(n437) );
  NOR2_X1 U464 ( .A1(n614), .A2(n613), .ZN(n625) );
  INV_X1 U465 ( .A(KEYINPUT34), .ZN(n406) );
  INV_X1 U466 ( .A(KEYINPUT19), .ZN(n410) );
  XNOR2_X1 U467 ( .A(KEYINPUT70), .B(KEYINPUT23), .ZN(n510) );
  XOR2_X1 U468 ( .A(G134), .B(KEYINPUT104), .Z(n461) );
  XOR2_X1 U469 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n466) );
  XNOR2_X1 U470 ( .A(n419), .B(n415), .ZN(n475) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n420), .B(n472), .ZN(n419) );
  NOR2_X1 U473 ( .A1(n630), .A2(n426), .ZN(n425) );
  NAND2_X1 U474 ( .A1(n762), .A2(KEYINPUT36), .ZN(n426) );
  AND2_X1 U475 ( .A1(n430), .A2(n429), .ZN(n428) );
  INV_X1 U476 ( .A(KEYINPUT36), .ZN(n429) );
  NAND2_X1 U477 ( .A1(n401), .A2(n400), .ZN(n399) );
  INV_X1 U478 ( .A(G478), .ZN(n469) );
  NOR2_X1 U479 ( .A1(n780), .A2(n436), .ZN(n781) );
  XOR2_X1 U480 ( .A(KEYINPUT13), .B(G475), .Z(n374) );
  XNOR2_X1 U481 ( .A(KEYINPUT87), .B(KEYINPUT35), .ZN(n375) );
  XOR2_X1 U482 ( .A(KEYINPUT91), .B(KEYINPUT33), .Z(n376) );
  AND2_X1 U483 ( .A1(n563), .A2(KEYINPUT44), .ZN(n377) );
  XNOR2_X2 U484 ( .A(n530), .B(KEYINPUT1), .ZN(n378) );
  XNOR2_X1 U485 ( .A(n530), .B(KEYINPUT1), .ZN(n543) );
  BUF_X1 U486 ( .A(n465), .Z(n379) );
  AND2_X2 U487 ( .A1(n534), .A2(n555), .ZN(n734) );
  BUF_X1 U488 ( .A(n564), .Z(n566) );
  XNOR2_X1 U489 ( .A(n496), .B(n507), .ZN(n719) );
  AND2_X1 U490 ( .A1(n546), .A2(n607), .ZN(n547) );
  BUF_X1 U491 ( .A(n581), .Z(n380) );
  NOR2_X1 U492 ( .A1(n731), .A2(n384), .ZN(n381) );
  AND2_X1 U493 ( .A1(n383), .A2(n585), .ZN(n382) );
  INV_X1 U494 ( .A(n586), .ZN(n383) );
  OR2_X1 U495 ( .A1(KEYINPUT81), .A2(n586), .ZN(n384) );
  BUF_X1 U496 ( .A(n633), .Z(n385) );
  XNOR2_X2 U497 ( .A(n408), .B(KEYINPUT39), .ZN(n633) );
  INV_X1 U498 ( .A(n373), .ZN(n528) );
  XNOR2_X1 U499 ( .A(n483), .B(n482), .ZN(n386) );
  XNOR2_X1 U500 ( .A(n483), .B(n482), .ZN(n548) );
  BUF_X1 U501 ( .A(n691), .Z(n387) );
  XNOR2_X1 U502 ( .A(n405), .B(n550), .ZN(n691) );
  NAND2_X1 U503 ( .A1(n615), .A2(n440), .ZN(n408) );
  BUF_X1 U504 ( .A(n772), .Z(n389) );
  XNOR2_X1 U505 ( .A(n553), .B(n376), .ZN(n772) );
  NAND2_X1 U506 ( .A1(n386), .A2(n498), .ZN(n390) );
  NAND2_X1 U507 ( .A1(n548), .A2(n498), .ZN(n539) );
  NAND2_X1 U508 ( .A1(n404), .A2(n403), .ZN(n402) );
  BUF_X1 U509 ( .A(n676), .Z(n391) );
  AND2_X1 U510 ( .A1(n559), .A2(n377), .ZN(n565) );
  NOR2_X1 U511 ( .A1(n647), .A2(n637), .ZN(n394) );
  AND2_X1 U512 ( .A1(n451), .A2(G210), .ZN(n395) );
  NOR2_X2 U513 ( .A1(n597), .A2(n610), .ZN(n397) );
  XNOR2_X1 U514 ( .A(n537), .B(n437), .ZN(n413) );
  OR2_X4 U515 ( .A1(n402), .A2(n398), .ZN(n530) );
  NOR2_X1 U516 ( .A1(n719), .A2(n399), .ZN(n398) );
  NAND2_X1 U517 ( .A1(n497), .A2(G902), .ZN(n403) );
  NAND2_X1 U518 ( .A1(n719), .A2(n497), .ZN(n404) );
  NAND2_X1 U519 ( .A1(n772), .A2(n435), .ZN(n407) );
  NAND2_X1 U520 ( .A1(n547), .A2(n386), .ZN(n405) );
  NAND2_X1 U521 ( .A1(n411), .A2(n569), .ZN(n571) );
  XNOR2_X1 U522 ( .A(n412), .B(KEYINPUT89), .ZN(n411) );
  NAND2_X1 U523 ( .A1(n414), .A2(n413), .ZN(n412) );
  NAND2_X1 U524 ( .A1(n439), .A2(n438), .ZN(n414) );
  OR2_X2 U525 ( .A1(n590), .A2(n610), .ZN(n592) );
  AND2_X2 U526 ( .A1(n595), .A2(n594), .ZN(n615) );
  NAND2_X1 U527 ( .A1(n661), .A2(n691), .ZN(n564) );
  INV_X1 U528 ( .A(n534), .ZN(n554) );
  NAND2_X1 U529 ( .A1(n711), .A2(n400), .ZN(n423) );
  NAND2_X1 U530 ( .A1(n433), .A2(n762), .ZN(n628) );
  NAND2_X1 U531 ( .A1(n427), .A2(n424), .ZN(n612) );
  NAND2_X1 U532 ( .A1(n433), .A2(n425), .ZN(n424) );
  NOR2_X1 U533 ( .A1(n432), .A2(n428), .ZN(n427) );
  NAND2_X1 U534 ( .A1(n431), .A2(n762), .ZN(n430) );
  INV_X1 U535 ( .A(n630), .ZN(n431) );
  XNOR2_X2 U536 ( .A(n462), .B(n434), .ZN(n487) );
  XNOR2_X2 U537 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n434) );
  XNOR2_X2 U538 ( .A(G143), .B(G128), .ZN(n462) );
  INV_X1 U539 ( .A(n528), .ZN(n435) );
  INV_X1 U540 ( .A(n389), .ZN(n436) );
  INV_X1 U541 ( .A(n559), .ZN(n693) );
  XNOR2_X2 U542 ( .A(n558), .B(n375), .ZN(n559) );
  NAND2_X1 U543 ( .A1(n565), .A2(n566), .ZN(n438) );
  NAND2_X1 U544 ( .A1(n562), .A2(KEYINPUT66), .ZN(n439) );
  BUF_X1 U545 ( .A(n717), .Z(n705) );
  NOR2_X2 U546 ( .A1(n689), .A2(n787), .ZN(n623) );
  NAND2_X1 U547 ( .A1(n602), .A2(n601), .ZN(n604) );
  BUF_X1 U548 ( .A(n642), .Z(n666) );
  AND2_X1 U549 ( .A1(n763), .A2(n748), .ZN(n440) );
  AND2_X1 U550 ( .A1(n765), .A2(n750), .ZN(n441) );
  INV_X1 U551 ( .A(KEYINPUT75), .ZN(n603) );
  NAND2_X1 U552 ( .A1(n611), .A2(n578), .ZN(n545) );
  INV_X1 U553 ( .A(KEYINPUT85), .ZN(n636) );
  XNOR2_X1 U554 ( .A(n469), .B(KEYINPUT105), .ZN(n470) );
  INV_X1 U555 ( .A(KEYINPUT40), .ZN(n616) );
  INV_X1 U556 ( .A(KEYINPUT56), .ZN(n654) );
  BUF_X1 U557 ( .A(n661), .Z(n662) );
  XNOR2_X2 U558 ( .A(G146), .B(G125), .ZN(n473) );
  XNOR2_X1 U559 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n443) );
  XNOR2_X1 U560 ( .A(n473), .B(n443), .ZN(n446) );
  INV_X2 U561 ( .A(G953), .ZN(n680) );
  NAND2_X1 U562 ( .A1(n680), .A2(G224), .ZN(n444) );
  XNOR2_X1 U563 ( .A(n444), .B(KEYINPUT77), .ZN(n445) );
  XNOR2_X1 U564 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U565 ( .A(n487), .B(n447), .ZN(n448) );
  XNOR2_X1 U566 ( .A(n663), .B(n448), .ZN(n647) );
  NAND2_X1 U567 ( .A1(n400), .A2(n450), .ZN(n451) );
  AND2_X1 U568 ( .A1(n451), .A2(G214), .ZN(n610) );
  XNOR2_X1 U569 ( .A(n452), .B(KEYINPUT14), .ZN(n455) );
  NAND2_X1 U570 ( .A1(G952), .A2(n455), .ZN(n453) );
  XOR2_X1 U571 ( .A(KEYINPUT95), .B(n453), .Z(n778) );
  NOR2_X1 U572 ( .A1(G953), .A2(n778), .ZN(n454) );
  XNOR2_X1 U573 ( .A(n454), .B(KEYINPUT96), .ZN(n575) );
  NAND2_X1 U574 ( .A1(G902), .A2(n455), .ZN(n572) );
  INV_X1 U575 ( .A(G898), .ZN(n456) );
  NAND2_X1 U576 ( .A1(n456), .A2(G953), .ZN(n664) );
  NOR2_X1 U577 ( .A1(n572), .A2(n664), .ZN(n457) );
  OR2_X1 U578 ( .A1(n575), .A2(n457), .ZN(n458) );
  NAND2_X1 U579 ( .A1(n680), .A2(G234), .ZN(n459) );
  NAND2_X1 U580 ( .A1(n512), .A2(G217), .ZN(n464) );
  XNOR2_X1 U581 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n464), .B(n463), .ZN(n468) );
  XOR2_X1 U583 ( .A(n466), .B(n379), .Z(n467) );
  XNOR2_X1 U584 ( .A(n468), .B(n467), .ZN(n706) );
  NOR2_X1 U585 ( .A1(G902), .A2(n706), .ZN(n471) );
  NAND2_X1 U586 ( .A1(G214), .A2(n499), .ZN(n472) );
  XNOR2_X1 U587 ( .A(n473), .B(KEYINPUT10), .ZN(n518) );
  INV_X1 U588 ( .A(n490), .ZN(n474) );
  XNOR2_X1 U589 ( .A(n518), .B(n474), .ZN(n677) );
  XNOR2_X1 U590 ( .A(n475), .B(n677), .ZN(n711) );
  INV_X1 U591 ( .A(n637), .ZN(n476) );
  NAND2_X1 U592 ( .A1(n476), .A2(G234), .ZN(n477) );
  XNOR2_X1 U593 ( .A(n477), .B(KEYINPUT20), .ZN(n521) );
  INV_X1 U594 ( .A(n521), .ZN(n479) );
  INV_X1 U595 ( .A(G221), .ZN(n478) );
  OR2_X1 U596 ( .A1(n479), .A2(n478), .ZN(n481) );
  INV_X1 U597 ( .A(KEYINPUT21), .ZN(n480) );
  XNOR2_X1 U598 ( .A(n481), .B(n480), .ZN(n750) );
  XNOR2_X1 U599 ( .A(n484), .B(KEYINPUT71), .ZN(n485) );
  INV_X1 U600 ( .A(n485), .ZN(n486) );
  XNOR2_X2 U601 ( .A(n487), .B(n486), .ZN(n676) );
  XNOR2_X2 U602 ( .A(n676), .B(G146), .ZN(n507) );
  XNOR2_X1 U603 ( .A(n489), .B(n488), .ZN(n493) );
  NAND2_X1 U604 ( .A1(n680), .A2(G227), .ZN(n491) );
  XNOR2_X1 U605 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U606 ( .A(n493), .B(n492), .ZN(n495) );
  XNOR2_X1 U607 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U608 ( .A(KEYINPUT74), .B(G469), .ZN(n497) );
  INV_X1 U609 ( .A(n378), .ZN(n498) );
  NAND2_X1 U610 ( .A1(n499), .A2(G210), .ZN(n501) );
  XNOR2_X1 U611 ( .A(n501), .B(n500), .ZN(n503) );
  XNOR2_X1 U612 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U613 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U614 ( .A(n507), .B(n506), .ZN(n694) );
  OR2_X2 U615 ( .A1(n694), .A2(G902), .ZN(n508) );
  XNOR2_X2 U616 ( .A(n508), .B(G472), .ZN(n540) );
  XNOR2_X1 U617 ( .A(n509), .B(KEYINPUT24), .ZN(n511) );
  XNOR2_X1 U618 ( .A(n511), .B(n510), .ZN(n514) );
  NAND2_X1 U619 ( .A1(n512), .A2(G221), .ZN(n513) );
  XNOR2_X1 U620 ( .A(n514), .B(n513), .ZN(n520) );
  XNOR2_X1 U621 ( .A(n657), .B(KEYINPUT98), .ZN(n516) );
  XNOR2_X1 U622 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U623 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U624 ( .A(n520), .B(n519), .ZN(n702) );
  OR2_X1 U625 ( .A1(n702), .A2(G902), .ZN(n525) );
  NAND2_X1 U626 ( .A1(n521), .A2(G217), .ZN(n523) );
  XNOR2_X1 U627 ( .A(KEYINPUT99), .B(KEYINPUT25), .ZN(n522) );
  XNOR2_X1 U628 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X2 U629 ( .A(n525), .B(n524), .ZN(n751) );
  NAND2_X1 U630 ( .A1(n607), .A2(n751), .ZN(n526) );
  XNOR2_X1 U631 ( .A(n527), .B(KEYINPUT106), .ZN(n687) );
  AND2_X1 U632 ( .A1(n751), .A2(n750), .ZN(n748) );
  NAND2_X1 U633 ( .A1(n552), .A2(n540), .ZN(n757) );
  NOR2_X1 U634 ( .A1(n528), .A2(n757), .ZN(n529) );
  XOR2_X1 U635 ( .A(KEYINPUT31), .B(n529), .Z(n737) );
  NAND2_X1 U636 ( .A1(n530), .A2(n748), .ZN(n531) );
  NOR2_X1 U637 ( .A1(n531), .A2(n540), .ZN(n532) );
  NAND2_X1 U638 ( .A1(n435), .A2(n532), .ZN(n533) );
  XNOR2_X1 U639 ( .A(n533), .B(KEYINPUT101), .ZN(n725) );
  NOR2_X1 U640 ( .A1(n737), .A2(n725), .ZN(n535) );
  NOR2_X1 U641 ( .A1(n555), .A2(n534), .ZN(n736) );
  NOR2_X1 U642 ( .A1(n736), .A2(n734), .ZN(n768) );
  NOR2_X1 U643 ( .A1(n535), .A2(n768), .ZN(n536) );
  NOR2_X1 U644 ( .A1(n687), .A2(n536), .ZN(n537) );
  INV_X1 U645 ( .A(KEYINPUT110), .ZN(n538) );
  XNOR2_X1 U646 ( .A(n539), .B(n538), .ZN(n542) );
  XNOR2_X1 U647 ( .A(n540), .B(KEYINPUT109), .ZN(n590) );
  INV_X1 U648 ( .A(n751), .ZN(n578) );
  AND2_X1 U649 ( .A1(n590), .A2(n578), .ZN(n541) );
  NAND2_X1 U650 ( .A1(n542), .A2(n541), .ZN(n661) );
  INV_X1 U651 ( .A(KEYINPUT108), .ZN(n544) );
  XNOR2_X1 U652 ( .A(n545), .B(n544), .ZN(n546) );
  INV_X1 U653 ( .A(KEYINPUT79), .ZN(n549) );
  XNOR2_X1 U654 ( .A(n549), .B(KEYINPUT32), .ZN(n550) );
  INV_X1 U655 ( .A(n564), .ZN(n560) );
  INV_X1 U656 ( .A(n607), .ZN(n551) );
  NAND2_X1 U657 ( .A1(n551), .A2(n552), .ZN(n553) );
  NOR2_X1 U658 ( .A1(n555), .A2(n554), .ZN(n596) );
  XNOR2_X1 U659 ( .A(n596), .B(KEYINPUT78), .ZN(n556) );
  NAND2_X1 U660 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U661 ( .A1(n561), .A2(KEYINPUT44), .ZN(n562) );
  INV_X1 U662 ( .A(KEYINPUT66), .ZN(n563) );
  XOR2_X1 U663 ( .A(KEYINPUT90), .B(n566), .Z(n568) );
  NOR2_X1 U664 ( .A1(n693), .A2(KEYINPUT44), .ZN(n567) );
  NAND2_X1 U665 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U666 ( .A(n571), .B(n570), .ZN(n642) );
  NOR2_X1 U667 ( .A1(G900), .A2(n572), .ZN(n573) );
  AND2_X1 U668 ( .A1(G953), .A2(n573), .ZN(n574) );
  OR2_X1 U669 ( .A1(n575), .A2(n574), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n593), .A2(n750), .ZN(n576) );
  XNOR2_X1 U671 ( .A(n576), .B(KEYINPUT73), .ZN(n577) );
  NAND2_X1 U672 ( .A1(n578), .A2(n577), .ZN(n605) );
  NOR2_X1 U673 ( .A1(n590), .A2(n605), .ZN(n580) );
  XNOR2_X1 U674 ( .A(KEYINPUT113), .B(KEYINPUT28), .ZN(n579) );
  XNOR2_X1 U675 ( .A(n580), .B(n579), .ZN(n621) );
  INV_X1 U676 ( .A(n530), .ZN(n620) );
  INV_X1 U677 ( .A(n380), .ZN(n582) );
  INV_X1 U678 ( .A(n768), .ZN(n584) );
  NAND2_X1 U679 ( .A1(n584), .A2(KEYINPUT47), .ZN(n585) );
  NOR2_X1 U680 ( .A1(KEYINPUT81), .A2(KEYINPUT47), .ZN(n586) );
  INV_X1 U681 ( .A(n731), .ZN(n589) );
  NOR2_X1 U682 ( .A1(n768), .A2(KEYINPUT47), .ZN(n587) );
  NOR2_X1 U683 ( .A1(n587), .A2(KEYINPUT81), .ZN(n588) );
  NOR2_X1 U684 ( .A1(n589), .A2(n588), .ZN(n600) );
  INV_X1 U685 ( .A(KEYINPUT30), .ZN(n591) );
  XNOR2_X1 U686 ( .A(n592), .B(n591), .ZN(n595) );
  AND2_X1 U687 ( .A1(n530), .A2(n593), .ZN(n594) );
  NAND2_X1 U688 ( .A1(n596), .A2(n748), .ZN(n598) );
  NOR2_X1 U689 ( .A1(n598), .A2(n630), .ZN(n599) );
  AND2_X1 U690 ( .A1(n615), .A2(n599), .ZN(n730) );
  NOR2_X1 U691 ( .A1(n600), .A2(n730), .ZN(n601) );
  XNOR2_X1 U692 ( .A(n604), .B(n603), .ZN(n614) );
  INV_X1 U693 ( .A(n605), .ZN(n606) );
  NAND2_X1 U694 ( .A1(n734), .A2(n606), .ZN(n608) );
  OR2_X1 U695 ( .A1(n608), .A2(n607), .ZN(n609) );
  INV_X1 U696 ( .A(n610), .ZN(n762) );
  NAND2_X1 U697 ( .A1(n612), .A2(n611), .ZN(n739) );
  XOR2_X1 U698 ( .A(KEYINPUT88), .B(n739), .Z(n613) );
  NAND2_X1 U699 ( .A1(n633), .A2(n734), .ZN(n617) );
  INV_X1 U700 ( .A(n765), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n763), .A2(n762), .ZN(n767) );
  NOR2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U703 ( .A(n623), .B(KEYINPUT46), .ZN(n624) );
  XNOR2_X1 U704 ( .A(KEYINPUT72), .B(KEYINPUT48), .ZN(n626) );
  NOR2_X1 U705 ( .A1(n628), .A2(n378), .ZN(n629) );
  XOR2_X1 U706 ( .A(KEYINPUT43), .B(n629), .Z(n631) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n632), .B(KEYINPUT112), .ZN(n788) );
  NAND2_X1 U709 ( .A1(n385), .A2(n736), .ZN(n660) );
  NAND2_X1 U710 ( .A1(n788), .A2(n660), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n637), .A2(KEYINPUT2), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(n646) );
  NAND2_X1 U714 ( .A1(n741), .A2(KEYINPUT2), .ZN(n643) );
  INV_X1 U715 ( .A(n666), .ZN(n742) );
  NOR2_X1 U716 ( .A1(n643), .A2(n742), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n644), .B(KEYINPUT76), .ZN(n745) );
  AND2_X2 U718 ( .A1(n646), .A2(n645), .ZN(n717) );
  NAND2_X1 U719 ( .A1(n717), .A2(G210), .ZN(n651) );
  BUF_X1 U720 ( .A(n647), .Z(n648) );
  XNOR2_X1 U721 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n651), .B(n650), .ZN(n653) );
  INV_X1 U723 ( .A(G952), .ZN(n652) );
  NAND2_X1 U724 ( .A1(n653), .A2(n722), .ZN(n655) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(G51) );
  NAND2_X1 U726 ( .A1(n725), .A2(n734), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n656), .B(G104), .ZN(G6) );
  XNOR2_X1 U728 ( .A(n657), .B(KEYINPUT29), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n731), .A2(n736), .ZN(n658) );
  XOR2_X1 U730 ( .A(n659), .B(n658), .Z(G30) );
  XNOR2_X1 U731 ( .A(n660), .B(G134), .ZN(G36) );
  XNOR2_X1 U732 ( .A(n662), .B(G110), .ZN(G12) );
  BUF_X1 U733 ( .A(n663), .Z(n665) );
  NAND2_X1 U734 ( .A1(n665), .A2(n664), .ZN(n674) );
  NAND2_X1 U735 ( .A1(n666), .A2(n680), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n667), .B(KEYINPUT124), .ZN(n672) );
  XOR2_X1 U737 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n669) );
  NAND2_X1 U738 ( .A1(G224), .A2(G953), .ZN(n668) );
  XNOR2_X1 U739 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U740 ( .A1(n670), .A2(G898), .ZN(n671) );
  NAND2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U742 ( .A(n674), .B(n673), .Z(G69) );
  INV_X1 U743 ( .A(KEYINPUT70), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n391), .B(n675), .ZN(n678) );
  XNOR2_X1 U745 ( .A(n678), .B(n677), .ZN(n682) );
  XOR2_X1 U746 ( .A(n682), .B(n679), .Z(n681) );
  NAND2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n686) );
  XNOR2_X1 U748 ( .A(G227), .B(n682), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n683), .A2(G900), .ZN(n684) );
  NAND2_X1 U750 ( .A1(n684), .A2(G953), .ZN(n685) );
  NAND2_X1 U751 ( .A1(n686), .A2(n685), .ZN(G72) );
  XOR2_X1 U752 ( .A(n687), .B(G101), .Z(G3) );
  XNOR2_X1 U753 ( .A(G131), .B(KEYINPUT127), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n689), .B(n688), .ZN(G33) );
  XNOR2_X1 U755 ( .A(G119), .B(KEYINPUT126), .ZN(n690) );
  XNOR2_X1 U756 ( .A(n387), .B(n690), .ZN(G21) );
  XNOR2_X1 U757 ( .A(G122), .B(KEYINPUT125), .ZN(n692) );
  XNOR2_X1 U758 ( .A(n693), .B(n692), .ZN(G24) );
  NAND2_X1 U759 ( .A1(n717), .A2(G472), .ZN(n697) );
  BUF_X1 U760 ( .A(n694), .Z(n695) );
  XNOR2_X1 U761 ( .A(n697), .B(n696), .ZN(n698) );
  NAND2_X1 U762 ( .A1(n698), .A2(n722), .ZN(n701) );
  XOR2_X1 U763 ( .A(KEYINPUT114), .B(KEYINPUT63), .Z(n699) );
  XNOR2_X1 U764 ( .A(n699), .B(KEYINPUT93), .ZN(n700) );
  XNOR2_X1 U765 ( .A(n701), .B(n700), .ZN(G57) );
  NAND2_X1 U766 ( .A1(n705), .A2(G217), .ZN(n703) );
  XNOR2_X1 U767 ( .A(n703), .B(n702), .ZN(n704) );
  INV_X1 U768 ( .A(n722), .ZN(n709) );
  NOR2_X1 U769 ( .A1(n704), .A2(n709), .ZN(G66) );
  NAND2_X1 U770 ( .A1(n705), .A2(G478), .ZN(n708) );
  XNOR2_X1 U771 ( .A(n706), .B(KEYINPUT122), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n708), .B(n707), .ZN(n710) );
  NOR2_X1 U773 ( .A1(n710), .A2(n709), .ZN(G63) );
  NAND2_X1 U774 ( .A1(n717), .A2(G475), .ZN(n713) );
  XNOR2_X1 U775 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U776 ( .A1(n714), .A2(n722), .ZN(n716) );
  XOR2_X1 U777 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n715) );
  XNOR2_X1 U778 ( .A(n716), .B(n715), .ZN(G60) );
  NAND2_X1 U779 ( .A1(n717), .A2(G469), .ZN(n721) );
  XNOR2_X1 U780 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n718) );
  XNOR2_X1 U781 ( .A(n721), .B(n720), .ZN(n723) );
  NAND2_X1 U782 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U783 ( .A(n724), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U784 ( .A1(n725), .A2(n736), .ZN(n727) );
  XOR2_X1 U785 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n726) );
  XNOR2_X1 U786 ( .A(n727), .B(n726), .ZN(n729) );
  XOR2_X1 U787 ( .A(G107), .B(KEYINPUT115), .Z(n728) );
  XNOR2_X1 U788 ( .A(n729), .B(n728), .ZN(G9) );
  XOR2_X1 U789 ( .A(G143), .B(n730), .Z(G45) );
  NAND2_X1 U790 ( .A1(n731), .A2(n734), .ZN(n732) );
  XNOR2_X1 U791 ( .A(n732), .B(KEYINPUT116), .ZN(n733) );
  XNOR2_X1 U792 ( .A(G146), .B(n733), .ZN(G48) );
  NAND2_X1 U793 ( .A1(n737), .A2(n734), .ZN(n735) );
  XNOR2_X1 U794 ( .A(n735), .B(G113), .ZN(G15) );
  NAND2_X1 U795 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U796 ( .A(n738), .B(G116), .ZN(G18) );
  XOR2_X1 U797 ( .A(G125), .B(n739), .Z(n740) );
  XNOR2_X1 U798 ( .A(n740), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U799 ( .A(KEYINPUT85), .B(n741), .ZN(n743) );
  NOR2_X1 U800 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U801 ( .A1(n744), .A2(KEYINPUT2), .ZN(n746) );
  NOR2_X1 U802 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U803 ( .A(KEYINPUT84), .B(n747), .Z(n784) );
  NOR2_X1 U804 ( .A1(n378), .A2(n748), .ZN(n749) );
  XOR2_X1 U805 ( .A(KEYINPUT50), .B(n749), .Z(n755) );
  NOR2_X1 U806 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U807 ( .A(KEYINPUT49), .B(n752), .Z(n753) );
  NOR2_X1 U808 ( .A1(n753), .A2(n540), .ZN(n754) );
  NAND2_X1 U809 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U810 ( .A(KEYINPUT117), .B(n756), .Z(n758) );
  AND2_X1 U811 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U812 ( .A(n759), .B(KEYINPUT51), .ZN(n760) );
  XNOR2_X1 U813 ( .A(n760), .B(KEYINPUT118), .ZN(n761) );
  NAND2_X1 U814 ( .A1(n761), .A2(n779), .ZN(n774) );
  NOR2_X1 U815 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U816 ( .A(n764), .B(KEYINPUT119), .ZN(n766) );
  NAND2_X1 U817 ( .A1(n766), .A2(n765), .ZN(n770) );
  OR2_X1 U818 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U819 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U820 ( .A1(n389), .A2(n771), .ZN(n773) );
  NAND2_X1 U821 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U822 ( .A(n775), .B(KEYINPUT120), .ZN(n776) );
  XOR2_X1 U823 ( .A(KEYINPUT52), .B(n776), .Z(n777) );
  NOR2_X1 U824 ( .A1(n778), .A2(n777), .ZN(n782) );
  INV_X1 U825 ( .A(n779), .ZN(n780) );
  NOR2_X1 U826 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U827 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U828 ( .A1(n785), .A2(G953), .ZN(n786) );
  XNOR2_X1 U829 ( .A(n786), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U830 ( .A(n787), .B(G137), .Z(G39) );
  XNOR2_X1 U831 ( .A(G140), .B(n788), .ZN(G42) );
endmodule

