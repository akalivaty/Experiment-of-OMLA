//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G137), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(G137), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n194), .A3(new_n197), .A4(new_n192), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n205), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n193), .A2(G134), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n190), .A2(G137), .ZN(new_n213));
  OAI21_X1  g027(.A(G131), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n198), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n201), .A2(new_n203), .A3(new_n216), .A4(G128), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n218), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(new_n219), .B2(new_n209), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n199), .A2(new_n211), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g035(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n222));
  OAI21_X1  g036(.A(new_n188), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g037(.A1(KEYINPUT2), .A2(G113), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT2), .A2(G113), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n224), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G116), .B(G119), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n229), .B(new_n224), .C1(new_n226), .C2(new_n227), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n221), .A2(KEYINPUT30), .ZN(new_n234));
  INV_X1    g048(.A(new_n222), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n220), .A2(new_n198), .A3(new_n214), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n196), .A2(new_n198), .B1(new_n208), .B2(new_n210), .ZN(new_n237));
  OAI211_X1 g051(.A(KEYINPUT65), .B(new_n235), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n223), .A2(new_n233), .A3(new_n234), .A4(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT31), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(G101), .ZN(new_n243));
  NOR2_X1   g057(.A1(G237), .A2(G953), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G210), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n243), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n233), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n199), .A2(new_n211), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n220), .A2(new_n198), .A3(new_n214), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n240), .A2(new_n241), .A3(new_n246), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n249), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT65), .B1(new_n252), .B2(new_n235), .ZN(new_n253));
  AOI211_X1 g067(.A(new_n188), .B(new_n222), .C1(new_n248), .C2(new_n249), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n255), .A2(KEYINPUT67), .A3(new_n233), .A4(new_n234), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n239), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n256), .A2(new_n246), .A3(new_n250), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT31), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n236), .B2(new_n237), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n248), .A2(KEYINPUT68), .A3(new_n249), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(new_n247), .ZN(new_n266));
  INV_X1    g080(.A(new_n246), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n250), .A2(new_n268), .A3(KEYINPUT28), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n251), .A2(new_n260), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT32), .ZN(new_n272));
  NOR2_X1   g086(.A1(G472), .A2(G902), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n272), .B1(new_n271), .B2(new_n273), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G472), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n278));
  AOI211_X1 g092(.A(KEYINPUT28), .B(new_n233), .C1(new_n262), .C2(new_n263), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n250), .A2(new_n268), .A3(KEYINPUT28), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT29), .B(new_n246), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n266), .A2(new_n269), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n284), .A2(KEYINPUT69), .A3(KEYINPUT29), .A4(new_n246), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g100(.A(KEYINPUT70), .B(G902), .Z(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n278), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  AOI211_X1 g103(.A(KEYINPUT71), .B(new_n287), .C1(new_n283), .C2(new_n285), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n256), .A2(new_n267), .A3(new_n250), .A4(new_n258), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n284), .A2(new_n267), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n277), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n187), .B1(new_n276), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n271), .A2(new_n273), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT32), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n286), .A2(new_n288), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT71), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n286), .A2(new_n278), .A3(new_n288), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n296), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G472), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n302), .A2(KEYINPUT72), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G116), .B(G122), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT92), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n310), .ZN(new_n313));
  INV_X1    g127(.A(G107), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n202), .A2(G128), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n218), .A2(G143), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(new_n190), .ZN(new_n319));
  INV_X1    g133(.A(G116), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT14), .A3(G122), .ZN(new_n321));
  XOR2_X1   g135(.A(G116), .B(G122), .Z(new_n322));
  OAI211_X1 g136(.A(G107), .B(new_n321), .C1(new_n322), .C2(KEYINPUT14), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n315), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(new_n190), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT13), .ZN(new_n326));
  OAI21_X1  g140(.A(G134), .B1(new_n316), .B2(KEYINPUT13), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n313), .ZN(new_n329));
  OAI21_X1  g143(.A(G107), .B1(new_n329), .B2(new_n311), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n328), .B1(new_n330), .B2(new_n315), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT93), .B1(new_n324), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n315), .ZN(new_n333));
  INV_X1    g147(.A(new_n328), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT93), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n315), .A2(new_n319), .A3(new_n323), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  XOR2_X1   g152(.A(KEYINPUT9), .B(G234), .Z(new_n339));
  INV_X1    g153(.A(G953), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(G217), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n332), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n335), .A2(new_n337), .ZN(new_n343));
  INV_X1    g157(.A(new_n341), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(KEYINPUT93), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n288), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT94), .ZN(new_n347));
  INV_X1    g161(.A(G478), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n347), .B1(KEYINPUT15), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(KEYINPUT15), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n346), .B2(KEYINPUT94), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n349), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G475), .ZN(new_n353));
  INV_X1    g167(.A(G902), .ZN(new_n354));
  NAND2_X1  g168(.A1(KEYINPUT75), .A2(G125), .ZN(new_n355));
  INV_X1    g169(.A(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(KEYINPUT75), .A2(G125), .A3(G140), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT16), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT16), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n356), .A3(G125), .ZN(new_n362));
  AOI21_X1  g176(.A(G146), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n361), .B1(new_n357), .B2(new_n358), .ZN(new_n364));
  INV_X1    g178(.A(new_n362), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n364), .A2(new_n200), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT90), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G143), .ZN(new_n369));
  INV_X1    g183(.A(G237), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n340), .A3(G214), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(G143), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n202), .A2(KEYINPUT90), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(G214), .B2(new_n244), .ZN(new_n375));
  OAI21_X1  g189(.A(G131), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT17), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n371), .A2(new_n369), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n244), .A2(G214), .B1(new_n368), .B2(G143), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n378), .B(new_n197), .C1(new_n379), .C2(new_n369), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT17), .B(G131), .C1(new_n373), .C2(new_n375), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n367), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G113), .B(G122), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n384), .B(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G125), .B(G140), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n200), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(new_n359), .B2(new_n200), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n371), .A2(new_n372), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n374), .ZN(new_n391));
  AND4_X1   g205(.A1(KEYINPUT18), .A2(new_n391), .A3(G131), .A4(new_n378), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n391), .A2(new_n378), .B1(KEYINPUT18), .B2(G131), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n383), .A2(new_n386), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n360), .A2(G146), .A3(new_n362), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT76), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n366), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n376), .A2(new_n380), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n387), .A2(KEYINPUT19), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT19), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n357), .B2(new_n358), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n200), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n397), .A2(new_n399), .A3(new_n400), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n386), .B1(new_n405), .B2(new_n394), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n353), .B(new_n354), .C1(new_n395), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT20), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT91), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT91), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n410), .A3(KEYINPUT20), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n407), .A2(KEYINPUT20), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n386), .B1(new_n383), .B2(new_n394), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n354), .B1(new_n395), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G475), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G952), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(G953), .ZN(new_n419));
  INV_X1    g233(.A(G234), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(new_n370), .ZN(new_n421));
  AOI211_X1 g235(.A(new_n340), .B(new_n288), .C1(G234), .C2(G237), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT21), .B(G898), .Z(new_n424));
  OAI21_X1  g238(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n425), .B(KEYINPUT95), .Z(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n352), .A2(new_n417), .A3(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(G119), .B(G128), .Z(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT73), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT24), .B(G110), .Z(new_n431));
  AOI21_X1  g245(.A(new_n367), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT23), .B1(new_n218), .B2(G119), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT74), .B1(new_n218), .B2(G119), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G110), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n397), .A2(new_n399), .A3(new_n388), .ZN(new_n438));
  OAI22_X1  g252(.A1(new_n430), .A2(new_n431), .B1(new_n435), .B2(G110), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n438), .A2(KEYINPUT77), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT77), .B1(new_n438), .B2(new_n439), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT78), .B(KEYINPUT22), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(G137), .ZN(new_n444));
  INV_X1    g258(.A(G221), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n445), .A2(new_n420), .A3(G953), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n444), .B(new_n446), .Z(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n437), .B(new_n447), .C1(new_n440), .C2(new_n441), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT25), .B1(new_n451), .B2(new_n287), .ZN(new_n452));
  OAI21_X1  g266(.A(G217), .B1(new_n287), .B2(new_n420), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT25), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n449), .A2(new_n455), .A3(new_n288), .A4(new_n450), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n454), .A2(G902), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n449), .A2(new_n458), .A3(new_n450), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n298), .A2(new_n308), .A3(new_n428), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n445), .B1(new_n339), .B2(new_n354), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n464));
  INV_X1    g278(.A(new_n217), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT80), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT80), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n468), .B(KEYINPUT1), .C1(new_n202), .C2(G146), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(G128), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n465), .B1(new_n470), .B2(new_n204), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n385), .A2(G107), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n385), .A2(G107), .ZN(new_n474));
  OAI21_X1  g288(.A(G101), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT3), .B1(new_n385), .B2(G107), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n314), .A3(G104), .ZN(new_n478));
  INV_X1    g292(.A(G101), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n476), .A2(new_n478), .A3(new_n479), .A4(new_n472), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n471), .A2(KEYINPUT81), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT81), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n469), .A2(G128), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n468), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n204), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n217), .ZN(new_n487));
  INV_X1    g301(.A(new_n481), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI22_X1  g303(.A1(new_n482), .A2(new_n489), .B1(new_n488), .B2(new_n220), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT12), .B1(new_n490), .B2(new_n199), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n488), .A2(new_n220), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT81), .B1(new_n471), .B2(new_n481), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n487), .A2(new_n483), .A3(new_n488), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT12), .ZN(new_n496));
  INV_X1    g310(.A(new_n199), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n464), .B1(new_n491), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT10), .B1(new_n493), .B2(new_n494), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n476), .A2(new_n478), .A3(new_n472), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G101), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(KEYINPUT4), .A3(new_n480), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT4), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n504), .A3(G101), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n211), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n488), .A2(KEYINPUT10), .A3(new_n220), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n500), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n497), .ZN(new_n510));
  XNOR2_X1  g324(.A(G110), .B(G140), .ZN(new_n511));
  INV_X1    g325(.A(G227), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(G953), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n511), .B(new_n513), .Z(new_n514));
  NAND3_X1  g328(.A1(new_n490), .A2(KEYINPUT12), .A3(new_n199), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n496), .B1(new_n495), .B2(new_n497), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT83), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n499), .A2(new_n510), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT82), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n199), .B1(new_n500), .B2(new_n508), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n510), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n514), .ZN(new_n522));
  OAI211_X1 g336(.A(KEYINPUT82), .B(new_n199), .C1(new_n500), .C2(new_n508), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G469), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n288), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT84), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n287), .B1(new_n518), .B2(new_n524), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(KEYINPUT84), .A3(new_n526), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n515), .A2(new_n516), .B1(new_n509), .B2(new_n497), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT79), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n522), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n521), .B(new_n523), .C1(new_n533), .C2(KEYINPUT79), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n354), .B(new_n535), .C1(new_n536), .C2(new_n522), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G469), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n463), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  OR3_X1    g353(.A1(new_n220), .A2(KEYINPUT87), .A3(G125), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n208), .A2(G125), .A3(new_n210), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT87), .B1(new_n220), .B2(G125), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n340), .A2(G224), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n233), .A2(new_n505), .A3(new_n503), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT5), .ZN(new_n547));
  INV_X1    g361(.A(G119), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(G116), .ZN(new_n549));
  OAI211_X1 g363(.A(G113), .B(new_n549), .C1(new_n230), .C2(new_n547), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n488), .A2(new_n232), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G122), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT86), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n552), .A2(new_n554), .B1(new_n555), .B2(KEYINPUT6), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(KEYINPUT6), .ZN(new_n557));
  AOI211_X1 g371(.A(new_n553), .B(new_n557), .C1(new_n546), .C2(new_n551), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n546), .A2(new_n553), .A3(new_n551), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n545), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n550), .A2(new_n232), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n481), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT88), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n551), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n553), .B(KEYINPUT8), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n562), .A2(KEYINPUT88), .A3(new_n481), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n541), .A2(KEYINPUT89), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n571), .A2(new_n541), .A3(new_n540), .A4(new_n542), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n543), .A2(new_n570), .A3(new_n569), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n568), .A2(new_n572), .A3(new_n573), .A4(new_n560), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n354), .ZN(new_n575));
  OAI21_X1  g389(.A(G210), .B1(G237), .B2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n561), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n574), .A2(new_n354), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n552), .A2(new_n554), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n557), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n552), .A2(new_n555), .A3(KEYINPUT6), .A4(new_n554), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n560), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n545), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n576), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G214), .B1(G237), .B2(G902), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT85), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n539), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n462), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n479), .ZN(G3));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n271), .A2(new_n288), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n596), .A2(G472), .B1(new_n273), .B2(new_n271), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n539), .A2(new_n595), .A3(new_n461), .A4(new_n597), .ZN(new_n598));
  AND4_X1   g412(.A1(KEYINPUT84), .A2(new_n525), .A3(new_n526), .A4(new_n288), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT84), .B1(new_n530), .B2(new_n526), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n538), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n463), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n601), .A2(new_n597), .A3(new_n602), .A4(new_n461), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT96), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT33), .B1(new_n342), .B2(new_n345), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n343), .A2(KEYINPUT98), .A3(new_n341), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n341), .A2(KEYINPUT98), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n335), .A2(new_n337), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n607), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(G478), .B(new_n288), .C1(new_n606), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n346), .A2(new_n348), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n417), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n617), .B(new_n577), .C1(new_n561), .C2(new_n575), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n588), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n587), .B2(KEYINPUT97), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n616), .A2(new_n426), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n605), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  INV_X1    g439(.A(new_n411), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n410), .B1(new_n407), .B2(KEYINPUT20), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT99), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n409), .A2(new_n629), .A3(new_n411), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n416), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n412), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n426), .B(KEYINPUT100), .Z(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(new_n620), .A3(new_n352), .A4(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n605), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NOR2_X1   g452(.A1(new_n448), .A2(KEYINPUT36), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n442), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n442), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n458), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n457), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n428), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n539), .A2(new_n645), .A3(new_n591), .A4(new_n597), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G110), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  OAI21_X1  g463(.A(new_n421), .B1(new_n423), .B2(G900), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n632), .A2(new_n352), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n298), .A2(new_n308), .A3(new_n620), .A4(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n529), .A2(new_n531), .B1(G469), .B2(new_n537), .ZN(new_n654));
  INV_X1    g468(.A(new_n644), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n654), .A2(new_n463), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(new_n218), .ZN(G30));
  INV_X1    g473(.A(new_n539), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n650), .B(KEYINPUT39), .Z(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n352), .A2(new_n417), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n663), .B2(KEYINPUT40), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n587), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n587), .A2(new_n667), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(KEYINPUT38), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(KEYINPUT38), .ZN(new_n673));
  INV_X1    g487(.A(new_n588), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n267), .B1(new_n240), .B2(new_n250), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n250), .A2(new_n268), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n354), .B1(new_n678), .B2(new_n246), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n644), .B1(new_n302), .B2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n664), .A2(new_n666), .A3(new_n675), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  INV_X1    g497(.A(new_n650), .ZN(new_n684));
  AOI221_X4 g498(.A(new_n684), .B1(new_n612), .B2(new_n613), .C1(new_n413), .C2(new_n416), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n620), .A3(KEYINPUT103), .ZN(new_n686));
  AND4_X1   g500(.A1(new_n602), .A2(new_n686), .A3(new_n601), .A4(new_n644), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n688));
  INV_X1    g502(.A(new_n685), .ZN(new_n689));
  INV_X1    g503(.A(new_n620), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n687), .A2(new_n298), .A3(new_n308), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  AND3_X1   g507(.A1(new_n298), .A2(new_n461), .A3(new_n308), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n530), .A2(new_n526), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n532), .A2(new_n602), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n694), .A2(new_n695), .A3(new_n622), .A4(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n298), .A2(new_n697), .A3(new_n308), .A4(new_n461), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT104), .B1(new_n699), .B2(new_n621), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT41), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G113), .ZN(G15));
  NOR2_X1   g517(.A1(new_n699), .A2(new_n634), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n320), .ZN(G18));
  NAND4_X1  g519(.A1(new_n298), .A2(new_n308), .A3(new_n620), .A4(new_n645), .ZN(new_n706));
  INV_X1    g520(.A(new_n697), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n548), .ZN(G21));
  NAND2_X1  g523(.A1(new_n596), .A2(G472), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n246), .B1(new_n284), .B2(KEYINPUT105), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(KEYINPUT105), .B2(new_n284), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n251), .A2(new_n260), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n273), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n460), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n690), .A2(new_n665), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n697), .A2(new_n716), .A3(new_n633), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NOR2_X1   g533(.A1(new_n715), .A2(new_n655), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n697), .A2(new_n720), .A3(new_n620), .A4(new_n685), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  OAI21_X1  g536(.A(KEYINPUT106), .B1(new_n654), .B2(new_n463), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n460), .B1(new_n302), .B2(new_n307), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n578), .A2(new_n586), .A3(new_n674), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n650), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n615), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n727), .A2(KEYINPUT42), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n601), .A2(new_n729), .A3(new_n602), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n723), .A2(new_n724), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n723), .A2(new_n725), .A3(new_n730), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n298), .A2(new_n461), .A3(new_n308), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n732), .A2(new_n733), .A3(new_n689), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n731), .B1(new_n734), .B2(KEYINPUT42), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT107), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  NOR3_X1   g551(.A1(new_n732), .A2(new_n733), .A3(new_n651), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n190), .ZN(G36));
  OR2_X1    g553(.A1(new_n536), .A2(new_n522), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n535), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT45), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n740), .A2(new_n743), .A3(new_n535), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n744), .A3(G469), .ZN(new_n745));
  NAND2_X1  g559(.A1(G469), .A2(G902), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n745), .A2(KEYINPUT46), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT46), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  INV_X1    g562(.A(new_n532), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n750), .A2(new_n463), .A3(new_n661), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n725), .B(KEYINPUT109), .Z(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n614), .A2(new_n413), .A3(new_n416), .ZN(new_n754));
  XNOR2_X1  g568(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(KEYINPUT108), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n756), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n760), .A2(new_n597), .A3(new_n655), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n753), .B1(new_n761), .B2(KEYINPUT44), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n751), .B(new_n762), .C1(KEYINPUT44), .C2(new_n761), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n750), .B2(new_n463), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n748), .A2(new_n749), .ZN(new_n767));
  OAI211_X1 g581(.A(KEYINPUT47), .B(new_n602), .C1(new_n767), .C2(new_n747), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n461), .B1(new_n298), .B2(new_n308), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n727), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n692), .B(new_n721), .C1(new_n657), .C2(new_n653), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n681), .A2(new_n717), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n539), .A2(new_n650), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n773), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n298), .A2(new_n308), .A3(new_n691), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n539), .A2(new_n644), .A3(new_n686), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n721), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n658), .ZN(new_n783));
  INV_X1    g597(.A(new_n777), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n782), .A2(new_n783), .A3(KEYINPUT52), .A4(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n778), .A2(new_n785), .A3(KEYINPUT113), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n781), .A2(new_n658), .A3(new_n773), .A4(new_n777), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n352), .B1(new_n631), .B2(new_n412), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n656), .A2(new_n298), .A3(new_n308), .A4(new_n792), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n710), .A2(new_n616), .A3(new_n644), .A4(new_n714), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n723), .A2(new_n730), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n726), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n791), .B1(new_n738), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n726), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n276), .A2(new_n297), .A3(new_n187), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT72), .B1(new_n302), .B2(new_n307), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n601), .A2(new_n602), .A3(new_n644), .A4(new_n792), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n723), .A2(new_n730), .A3(new_n794), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n798), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n732), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n694), .A3(new_n652), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(KEYINPUT111), .A3(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n797), .A2(new_n807), .A3(new_n735), .ZN(new_n808));
  INV_X1    g622(.A(new_n352), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n615), .B1(new_n809), .B2(new_n417), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(new_n591), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n598), .A2(new_n604), .A3(new_n633), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n646), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n812), .A2(new_n593), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n718), .B1(new_n699), .B2(new_n634), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n708), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n814), .A2(new_n701), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n808), .A2(new_n817), .A3(KEYINPUT112), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n797), .A2(new_n807), .A3(new_n735), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n814), .A2(new_n701), .A3(new_n816), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n790), .A2(new_n818), .A3(new_n819), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n781), .A2(new_n658), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(new_n825), .B2(new_n784), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT114), .B1(new_n826), .B2(new_n787), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n778), .A2(new_n785), .A3(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n827), .A2(new_n829), .A3(new_n817), .A4(new_n808), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT53), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n824), .A2(new_n831), .A3(KEYINPUT54), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT115), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n824), .A2(new_n831), .A3(new_n834), .A4(KEYINPUT54), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n701), .A2(new_n816), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n838), .A2(KEYINPUT116), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n819), .A3(new_n821), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n838), .A2(KEYINPUT116), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n814), .A3(new_n841), .A4(new_n790), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n830), .A2(new_n819), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n532), .A2(new_n696), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n463), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n766), .A2(new_n768), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n760), .ZN(new_n849));
  INV_X1    g663(.A(new_n421), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n716), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n753), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT117), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n674), .B1(new_n672), .B2(new_n673), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n855), .A2(new_n851), .A3(new_n707), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT50), .B1(new_n856), .B2(KEYINPUT118), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT50), .ZN(new_n859));
  INV_X1    g673(.A(new_n851), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n697), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n858), .B(new_n859), .C1(new_n861), .C2(new_n855), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n697), .A2(new_n850), .A3(new_n725), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n302), .A2(new_n680), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n864), .A2(new_n460), .A3(new_n865), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n866), .A2(new_n417), .A3(new_n614), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n864), .A2(new_n760), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT119), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n720), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n854), .A2(new_n863), .A3(new_n867), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n848), .A2(new_n853), .B1(new_n857), .B2(new_n862), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(KEYINPUT51), .A3(new_n867), .A4(new_n870), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n419), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n724), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT48), .Z(new_n878));
  NOR2_X1   g692(.A1(new_n866), .A2(new_n615), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n861), .A2(new_n690), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n876), .A2(new_n878), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n836), .A2(new_n837), .A3(new_n845), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n418), .A2(new_n340), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n881), .A2(new_n833), .A3(new_n845), .A4(new_n835), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT120), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n672), .A2(new_n673), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n846), .B(KEYINPUT49), .Z(new_n888));
  NOR4_X1   g702(.A1(new_n460), .A2(new_n754), .A3(new_n463), .A4(new_n590), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT110), .Z(new_n890));
  OR4_X1    g704(.A1(new_n887), .A2(new_n888), .A3(new_n890), .A4(new_n865), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n891), .ZN(G75));
  AOI21_X1  g706(.A(new_n288), .B1(new_n842), .B2(new_n844), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n577), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n583), .A2(new_n584), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n561), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT55), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n894), .B2(new_n895), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n340), .A2(G952), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(G51));
  NOR2_X1   g716(.A1(new_n746), .A2(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n842), .A2(new_n844), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n903), .B1(new_n905), .B2(new_n845), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n746), .A2(KEYINPUT57), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n525), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n893), .A2(G469), .A3(new_n742), .A4(new_n744), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n901), .B1(new_n909), .B2(new_n910), .ZN(G54));
  NAND3_X1  g725(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n395), .A2(new_n406), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n901), .ZN(new_n915));
  INV_X1    g729(.A(new_n913), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .A4(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT121), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n914), .A2(new_n920), .A3(new_n915), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(G60));
  OR2_X1    g736(.A1(new_n606), .A2(new_n611), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT122), .Z(new_n924));
  NAND3_X1  g738(.A1(new_n833), .A2(new_n845), .A3(new_n835), .ZN(new_n925));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT59), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n924), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n924), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n927), .B(new_n930), .C1(new_n905), .C2(new_n845), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n929), .A2(new_n931), .A3(new_n901), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT60), .Z(new_n934));
  NAND2_X1  g748(.A1(new_n904), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n451), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n904), .A2(new_n641), .A3(new_n642), .A4(new_n934), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n915), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G66));
  AOI21_X1  g754(.A(new_n340), .B1(new_n424), .B2(G224), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n822), .B2(new_n340), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n559), .B(new_n560), .C1(G898), .C2(new_n340), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n942), .B(new_n943), .Z(G69));
  NAND4_X1  g758(.A1(new_n694), .A2(new_n662), .A3(new_n725), .A4(new_n810), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n771), .A2(new_n763), .A3(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n774), .B(KEYINPUT123), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n682), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n947), .A2(KEYINPUT62), .A3(new_n682), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n340), .ZN(new_n953));
  NAND3_X1  g767(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n255), .A2(new_n234), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n401), .A2(new_n403), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n955), .B(new_n956), .Z(new_n957));
  NAND3_X1  g771(.A1(new_n953), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n512), .A2(G900), .A3(G953), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n751), .A2(new_n717), .A3(new_n724), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT124), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n735), .A3(new_n947), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n771), .A2(new_n806), .A3(new_n763), .ZN(new_n963));
  OR3_X1    g777(.A1(new_n962), .A2(KEYINPUT125), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT125), .B1(new_n962), .B2(new_n963), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n959), .B1(new_n966), .B2(G953), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n958), .B1(new_n967), .B2(new_n957), .ZN(G72));
  NAND3_X1  g782(.A1(new_n964), .A2(new_n817), .A3(new_n965), .ZN(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n277), .A2(new_n354), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(new_n971), .Z(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n901), .B1(new_n974), .B2(new_n294), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n952), .A2(new_n817), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n676), .B1(new_n976), .B2(new_n972), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n979), .B(new_n676), .C1(new_n976), .C2(new_n972), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n824), .A2(new_n831), .A3(new_n293), .A4(new_n973), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n982), .A2(new_n676), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n975), .A2(new_n981), .A3(new_n983), .ZN(G57));
endmodule


