//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1209, new_n1210, new_n1211, new_n1212, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0008(.A(KEYINPUT65), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n209), .B1(new_n210), .B2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G13), .ZN(new_n212));
  NAND4_X1  g0012(.A1(new_n212), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n231), .A2(G50), .A3(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n216), .B(new_n227), .C1(new_n230), .C2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  AOI21_X1  g0051(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G1), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT5), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT5), .A2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n252), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n262), .B1(new_n257), .B2(new_n258), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n265), .A2(G274), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n260), .A2(G270), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G33), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n269), .A2(new_n271), .A3(G264), .A4(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n269), .A2(new_n271), .A3(G257), .A4(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G303), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n272), .B(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n252), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n267), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G200), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G116), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n281), .A2(new_n228), .B1(G20), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G283), .ZN(new_n284));
  INV_X1    g0084(.A(G97), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n284), .B(new_n229), .C1(G33), .C2(new_n285), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n283), .A2(KEYINPUT20), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT20), .B1(new_n283), .B2(new_n286), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n281), .A2(new_n228), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n282), .B1(new_n261), .B2(G33), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n212), .A2(new_n229), .A3(G1), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n212), .A2(G1), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n295), .A2(KEYINPUT70), .A3(G20), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n291), .B(new_n292), .C1(new_n294), .C2(new_n296), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n298), .A2(new_n299), .A3(new_n282), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n267), .A2(new_n278), .A3(G190), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n280), .A2(new_n289), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n297), .B(new_n300), .C1(new_n288), .C2(new_n287), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(new_n279), .A3(G169), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT21), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n267), .A2(new_n278), .A3(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n304), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n304), .A2(new_n279), .A3(KEYINPUT21), .A4(G169), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n303), .A2(new_n307), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT84), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n309), .A2(new_n310), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT84), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(new_n314), .A3(new_n307), .A4(new_n303), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G20), .A2(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G150), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT8), .B(G58), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n229), .A2(G33), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT68), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n322), .A2(new_n323), .B1(G20), .B2(new_n203), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(KEYINPUT68), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n291), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT69), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n293), .A2(new_n290), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n202), .B1(new_n261), .B2(G20), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n328), .A2(new_n329), .B1(new_n202), .B2(new_n293), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n326), .A2(KEYINPUT69), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(KEYINPUT9), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT9), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n331), .B2(new_n333), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n276), .A2(G222), .A3(new_n273), .ZN(new_n338));
  INV_X1    g0138(.A(G77), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n276), .A2(G1698), .ZN(new_n340));
  INV_X1    g0140(.A(G223), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n338), .B1(new_n339), .B2(new_n276), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n252), .ZN(new_n343));
  AOI21_X1  g0143(.A(G1), .B1(new_n256), .B2(new_n253), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(new_n265), .A3(G274), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n265), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n346), .B1(G226), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT71), .B(G200), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n353), .B1(new_n355), .B2(new_n351), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n335), .A2(new_n337), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT10), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n332), .A2(new_n334), .ZN(new_n359));
  INV_X1    g0159(.A(G169), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n351), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n359), .B(new_n361), .C1(G179), .C2(new_n351), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n319), .B1(new_n261), .B2(G20), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n328), .B1(new_n293), .B2(new_n319), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n276), .B2(G20), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n270), .A2(G33), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT7), .B(new_n229), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT76), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n269), .A2(new_n271), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n229), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n374), .B2(new_n366), .ZN(new_n375));
  OAI21_X1  g0175(.A(G68), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G58), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n218), .ZN(new_n378));
  OAI21_X1  g0178(.A(G20), .B1(new_n378), .B2(new_n201), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n317), .A2(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT16), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n276), .A2(new_n366), .A3(G20), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT7), .B1(new_n373), .B2(new_n229), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n290), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n365), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT77), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT77), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(new_n365), .C1(new_n383), .C2(new_n388), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n265), .A2(G232), .A3(new_n347), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n345), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n269), .A2(new_n271), .A3(G226), .A4(G1698), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n269), .A2(new_n271), .A3(G223), .A4(new_n273), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n395), .B(new_n396), .C1(new_n268), .C2(new_n220), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n394), .B1(new_n397), .B2(new_n252), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(G169), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT78), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n345), .A2(new_n393), .A3(KEYINPUT78), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(G179), .B1(new_n397), .B2(new_n252), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n399), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n390), .A2(new_n392), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT18), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n397), .A2(new_n252), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n352), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n410), .A2(new_n403), .B1(new_n398), .B2(G200), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n365), .B(new_n411), .C1(new_n383), .C2(new_n388), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT79), .B1(new_n412), .B2(KEYINPUT80), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n367), .A2(new_n370), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n381), .B1(new_n414), .B2(G68), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n291), .B1(new_n415), .B2(KEYINPUT16), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n376), .A2(new_n382), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(KEYINPUT16), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT79), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(new_n419), .A3(new_n365), .A4(new_n411), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n413), .A2(new_n420), .A3(KEYINPUT17), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  OAI211_X1 g0222(.A(KEYINPUT79), .B(new_n422), .C1(new_n412), .C2(KEYINPUT80), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n390), .A2(new_n424), .A3(new_n392), .A4(new_n406), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n408), .A2(new_n421), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n345), .B1(new_n219), .B2(new_n348), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n269), .A2(new_n271), .A3(G232), .A4(G1698), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT73), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n276), .A2(KEYINPUT73), .A3(G232), .A4(G1698), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G97), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n276), .A2(G226), .A3(new_n273), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n430), .A2(new_n431), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n427), .B1(new_n434), .B2(new_n252), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT13), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI211_X1 g0237(.A(KEYINPUT13), .B(new_n427), .C1(new_n434), .C2(new_n252), .ZN(new_n438));
  OAI21_X1  g0238(.A(G169), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(KEYINPUT14), .B(G169), .C1(new_n437), .C2(new_n438), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n438), .B(KEYINPUT74), .ZN(new_n444));
  INV_X1    g0244(.A(G179), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n437), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n317), .A2(G50), .ZN(new_n449));
  XOR2_X1   g0249(.A(new_n449), .B(KEYINPUT75), .Z(new_n450));
  OAI22_X1  g0250(.A1(new_n320), .A2(new_n339), .B1(new_n229), .B2(G68), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n290), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT11), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n294), .A2(new_n296), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(new_n290), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n261), .A2(G20), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(G68), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT12), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n295), .A2(new_n460), .A3(G20), .A4(new_n218), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n294), .A2(new_n296), .A3(G68), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(new_n460), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n454), .A2(new_n455), .A3(new_n459), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n448), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n437), .A2(new_n352), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n444), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n464), .ZN(new_n468));
  OAI21_X1  g0268(.A(G200), .B1(new_n437), .B2(new_n438), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n349), .A2(G244), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n276), .A2(G232), .A3(new_n273), .ZN(new_n473));
  INV_X1    g0273(.A(G107), .ZN(new_n474));
  OAI221_X1 g0274(.A(new_n473), .B1(new_n474), .B2(new_n276), .C1(new_n340), .C2(new_n219), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n346), .B(new_n472), .C1(new_n475), .C2(new_n252), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n445), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT72), .ZN(new_n478));
  INV_X1    g0278(.A(new_n319), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n479), .A2(new_n317), .B1(G20), .B2(G77), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT15), .B(G87), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n320), .B2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(new_n290), .B1(new_n339), .B2(new_n456), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n457), .A2(G77), .A3(new_n458), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n476), .B2(G169), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n476), .A2(G190), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n489), .B(new_n490), .C1(new_n354), .C2(new_n476), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NOR4_X1   g0292(.A1(new_n363), .A2(new_n426), .A3(new_n471), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n259), .A2(new_n254), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(G257), .A3(new_n265), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n266), .A2(new_n263), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n269), .A2(new_n271), .A3(G244), .A4(new_n273), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(KEYINPUT81), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(KEYINPUT81), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n276), .A2(G244), .A3(new_n273), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n500), .A2(new_n284), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n497), .B1(new_n504), .B2(new_n252), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT82), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n505), .A2(new_n506), .A3(G190), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n505), .B2(G190), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G200), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(G107), .B1(new_n371), .B2(new_n375), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n474), .A2(KEYINPUT6), .A3(G97), .ZN(new_n513));
  XOR2_X1   g0313(.A(G97), .B(G107), .Z(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(G20), .B1(G77), .B2(new_n317), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n291), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n293), .A2(new_n285), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n328), .B1(G1), .B2(new_n268), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(new_n285), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n511), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n517), .A2(new_n520), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n505), .A2(G169), .ZN(new_n523));
  AOI211_X1 g0323(.A(G179), .B(new_n497), .C1(new_n252), .C2(new_n504), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n509), .A2(new_n521), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n269), .A2(new_n271), .A3(new_n229), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT22), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n276), .A2(new_n529), .A3(new_n229), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n268), .A2(new_n282), .A3(G20), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n229), .B2(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n474), .A2(KEYINPUT23), .A3(G20), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n531), .A2(new_n532), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n532), .B1(new_n531), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n290), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n519), .A2(new_n474), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n293), .A2(new_n474), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n542), .B(KEYINPUT25), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n269), .A2(new_n271), .A3(G257), .A4(G1698), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n269), .A2(new_n271), .A3(G250), .A4(new_n273), .ZN(new_n547));
  INV_X1    g0347(.A(G294), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n547), .C1(new_n268), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n252), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n260), .A2(G264), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n550), .A2(new_n496), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n445), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n549), .A2(new_n252), .B1(new_n260), .B2(G264), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n496), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n360), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n545), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n552), .A2(G200), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n555), .A2(G190), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n540), .B(new_n544), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n219), .A2(new_n273), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(G244), .B2(new_n273), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n562), .A2(new_n373), .B1(new_n268), .B2(new_n282), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n252), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n265), .A2(G274), .A3(new_n254), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT83), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n265), .A2(KEYINPUT83), .A3(G274), .A4(new_n254), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n252), .A2(new_n221), .A3(new_n254), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n564), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n360), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n276), .A2(new_n229), .A3(G68), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n229), .B1(new_n432), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(G87), .B2(new_n206), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n575), .B1(new_n320), .B2(new_n285), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n574), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n290), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n456), .A2(new_n481), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n519), .C2(new_n481), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n570), .B1(new_n563), .B2(new_n252), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(new_n445), .A3(new_n569), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n573), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n328), .B(G87), .C1(G1), .C2(new_n268), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n580), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n572), .A2(new_n355), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n583), .A2(G190), .A3(new_n569), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AND4_X1   g0390(.A1(new_n557), .A2(new_n560), .A3(new_n585), .A4(new_n590), .ZN(new_n591));
  AND4_X1   g0391(.A1(new_n316), .A2(new_n493), .A3(new_n526), .A4(new_n591), .ZN(G372));
  NAND2_X1  g0392(.A1(new_n389), .A2(new_n406), .ZN(new_n593));
  XNOR2_X1  g0393(.A(new_n593), .B(new_n424), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n487), .A2(new_n470), .B1(new_n448), .B2(new_n464), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n421), .A2(new_n423), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT86), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(KEYINPUT86), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n358), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n601), .A2(new_n362), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n590), .A2(new_n585), .A3(KEYINPUT85), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT85), .B1(new_n590), .B2(new_n585), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n557), .A2(new_n307), .A3(new_n313), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n526), .A2(new_n605), .A3(new_n560), .A4(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT26), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n522), .A2(new_n525), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n605), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n590), .A2(new_n585), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT26), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n607), .A2(new_n611), .A3(new_n585), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n493), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n602), .A2(new_n615), .ZN(G369));
  NAND2_X1  g0416(.A1(new_n313), .A2(new_n307), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n295), .A2(new_n229), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n618), .A2(KEYINPUT27), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(KEYINPUT27), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(G213), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G343), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n304), .A2(new_n623), .ZN(new_n624));
  MUX2_X1   g0424(.A(new_n617), .B(new_n316), .S(new_n624), .Z(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G330), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n545), .A2(new_n553), .A3(new_n556), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n623), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n545), .A2(new_n623), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n557), .A2(new_n560), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(KEYINPUT87), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n557), .A2(new_n623), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT87), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n631), .B(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n623), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n617), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n635), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n634), .A2(new_n641), .ZN(G399));
  INV_X1    g0442(.A(new_n214), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(G41), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n645), .A2(G1), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n234), .B2(new_n644), .ZN(new_n648));
  XOR2_X1   g0448(.A(new_n648), .B(KEYINPUT28), .Z(new_n649));
  INV_X1    g0449(.A(KEYINPUT31), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n279), .A2(new_n572), .A3(new_n445), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n651), .A2(new_n505), .A3(new_n552), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n564), .A2(new_n569), .A3(new_n571), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n308), .A2(new_n505), .A3(new_n554), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT30), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n583), .A2(new_n550), .A3(new_n551), .A4(new_n569), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n267), .A2(new_n278), .A3(G179), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT30), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(new_n505), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n652), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n623), .B1(new_n661), .B2(KEYINPUT88), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT88), .ZN(new_n663));
  AOI211_X1 g0463(.A(new_n663), .B(new_n652), .C1(new_n655), .C2(new_n660), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n650), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n316), .A2(new_n591), .A3(new_n526), .A4(new_n638), .ZN(new_n666));
  INV_X1    g0466(.A(new_n652), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n654), .A2(KEYINPUT30), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n659), .B1(new_n658), .B2(new_n505), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(KEYINPUT31), .A3(new_n623), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n665), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n608), .B1(new_n609), .B2(new_n612), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT89), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n605), .A2(KEYINPUT26), .A3(new_n610), .ZN(new_n677));
  OAI211_X1 g0477(.A(KEYINPUT89), .B(new_n608), .C1(new_n609), .C2(new_n612), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n607), .A2(new_n585), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n638), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n614), .A2(new_n638), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n673), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n649), .B1(new_n687), .B2(G1), .ZN(G364));
  NOR2_X1   g0488(.A1(new_n212), .A2(G20), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n261), .B1(new_n689), .B2(G45), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n644), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n228), .B1(G20), .B2(new_n360), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n352), .A2(G179), .A3(G200), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n229), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n373), .B1(new_n697), .B2(new_n548), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n229), .A2(G190), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(G179), .A3(new_n510), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n445), .A3(new_n510), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n701), .A2(G311), .B1(new_n703), .B2(G329), .ZN(new_n704));
  INV_X1    g0504(.A(G326), .ZN(new_n705));
  NOR4_X1   g0505(.A1(new_n229), .A2(new_n445), .A3(new_n352), .A4(new_n510), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n704), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n355), .A2(new_n445), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n229), .B1(new_n709), .B2(KEYINPUT91), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(KEYINPUT91), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n352), .ZN(new_n712));
  AOI211_X1 g0512(.A(new_n698), .B(new_n708), .C1(new_n712), .C2(G303), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n229), .A2(new_n445), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(new_n352), .A3(G200), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g0516(.A(KEYINPUT33), .B(G317), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(KEYINPUT93), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n717), .A2(KEYINPUT93), .ZN(new_n719));
  INV_X1    g0519(.A(G322), .ZN(new_n720));
  NOR4_X1   g0520(.A1(new_n229), .A2(new_n445), .A3(new_n352), .A4(G200), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n718), .A2(new_n719), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT94), .ZN(new_n724));
  INV_X1    g0524(.A(G283), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n711), .A2(G190), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n713), .B(new_n724), .C1(new_n725), .C2(new_n727), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n276), .B1(new_n722), .B2(new_n377), .C1(new_n202), .C2(new_n707), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n697), .A2(new_n285), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(G68), .B2(new_n716), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(KEYINPUT92), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n729), .B(new_n732), .C1(G77), .C2(new_n701), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n712), .A2(G87), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n726), .A2(G107), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT32), .ZN(new_n736));
  INV_X1    g0536(.A(G159), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n736), .B1(new_n702), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n703), .A2(KEYINPUT32), .A3(G159), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n731), .A2(KEYINPUT92), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n733), .A2(new_n734), .A3(new_n735), .A4(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n695), .B1(new_n728), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n694), .ZN(new_n746));
  NAND3_X1  g0546(.A1(G355), .A2(new_n214), .A3(new_n276), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n250), .A2(G45), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT90), .Z(new_n749));
  NOR2_X1   g0549(.A1(new_n643), .A2(new_n276), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(G45), .B2(new_n233), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n747), .B1(G116), .B2(new_n214), .C1(new_n749), .C2(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n693), .B(new_n742), .C1(new_n746), .C2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n745), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n753), .B1(new_n625), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n626), .A2(new_n693), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n625), .A2(G330), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(G396));
  NAND2_X1  g0558(.A1(new_n485), .A2(new_n623), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n491), .B(new_n759), .C1(new_n478), .C2(new_n486), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(new_n488), .B2(new_n759), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n684), .B(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n673), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT96), .Z(new_n764));
  AOI21_X1  g0564(.A(new_n692), .B1(new_n762), .B2(new_n673), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n707), .A2(new_n275), .B1(new_n282), .B2(new_n700), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(G283), .B2(new_n716), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT95), .Z(new_n769));
  NAND2_X1  g0569(.A1(new_n712), .A2(G107), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n373), .B1(new_n722), .B2(new_n548), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n730), .B(new_n771), .C1(G311), .C2(new_n703), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n726), .A2(G87), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n769), .A2(new_n770), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G132), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n276), .B1(new_n702), .B2(new_n775), .C1(new_n697), .C2(new_n377), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G159), .A2(new_n701), .B1(new_n706), .B2(G137), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n716), .A2(G150), .B1(new_n721), .B2(G143), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT34), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n780), .B2(new_n779), .ZN(new_n782));
  INV_X1    g0582(.A(new_n712), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n202), .A2(new_n783), .B1(new_n727), .B2(new_n218), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n774), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n694), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n694), .A2(new_n743), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n693), .B1(new_n339), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n786), .B(new_n788), .C1(new_n761), .C2(new_n744), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n766), .A2(new_n789), .ZN(G384));
  NOR2_X1   g0590(.A1(new_n689), .A2(new_n261), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n670), .A2(new_n663), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n667), .B(KEYINPUT88), .C1(new_n668), .C2(new_n669), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n792), .A2(KEYINPUT31), .A3(new_n623), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n665), .A2(new_n666), .A3(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n795), .A2(new_n761), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n464), .A2(new_n623), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n441), .A2(new_n442), .B1(new_n444), .B2(new_n446), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n470), .B(new_n797), .C1(new_n798), .C2(new_n468), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT98), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n465), .A2(KEYINPUT98), .A3(new_n470), .A4(new_n797), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n470), .A2(new_n798), .ZN(new_n804));
  INV_X1    g0604(.A(new_n797), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n415), .A2(KEYINPUT16), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n365), .B1(new_n388), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n621), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n426), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n621), .B(KEYINPUT100), .Z(new_n813));
  NAND3_X1  g0613(.A1(new_n390), .A2(new_n392), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT37), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n407), .A2(new_n814), .A3(new_n815), .A4(new_n412), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n809), .A2(new_n406), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT99), .ZN(new_n818));
  AND3_X1   g0618(.A1(new_n817), .A2(new_n818), .A3(new_n412), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(new_n817), .B2(new_n412), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n819), .A2(new_n820), .A3(new_n811), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n816), .B1(new_n821), .B2(new_n815), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n812), .A2(new_n822), .A3(KEYINPUT38), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT38), .B1(new_n812), .B2(new_n822), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n796), .B(new_n807), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT40), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT101), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n825), .A2(KEYINPUT101), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n594), .A2(new_n421), .A3(new_n423), .ZN(new_n832));
  INV_X1    g0632(.A(new_n814), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n593), .A2(new_n412), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT37), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n816), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT38), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n812), .A2(new_n822), .A3(KEYINPUT38), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n826), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n801), .A2(new_n802), .B1(new_n805), .B2(new_n804), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n795), .A2(new_n761), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n831), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n493), .A2(new_n795), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(G330), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n846), .B2(new_n847), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n683), .A2(new_n685), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n493), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n602), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n594), .A2(new_n813), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n614), .A2(new_n761), .A3(new_n638), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n487), .A2(new_n638), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n842), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n812), .A2(new_n822), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n840), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n855), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n823), .B2(new_n838), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n861), .A2(KEYINPUT39), .A3(new_n840), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n465), .A2(new_n623), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n854), .B(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n791), .B1(new_n851), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n870), .B2(new_n851), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n515), .B(KEYINPUT97), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT35), .ZN(new_n874));
  OAI211_X1 g0674(.A(G116), .B(new_n230), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n874), .B2(new_n873), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT36), .Z(new_n877));
  NOR3_X1   g0677(.A1(new_n233), .A2(new_n339), .A3(new_n378), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n218), .A2(G50), .ZN(new_n879));
  OAI211_X1 g0679(.A(G1), .B(new_n212), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n872), .A2(new_n877), .A3(new_n880), .ZN(G367));
  NOR3_X1   g0681(.A1(new_n243), .A2(new_n643), .A3(new_n276), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n746), .B1(new_n214), .B2(new_n481), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n692), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n697), .A2(new_n218), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(G150), .B2(new_n721), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT108), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n276), .B1(new_n715), .B2(new_n737), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n706), .A2(G143), .ZN(new_n889));
  XOR2_X1   g0689(.A(KEYINPUT109), .B(G137), .Z(new_n890));
  OAI22_X1  g0690(.A1(new_n702), .A2(new_n890), .B1(new_n700), .B2(new_n202), .ZN(new_n891));
  NOR4_X1   g0691(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n891), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n892), .B1(new_n377), .B2(new_n783), .C1(new_n339), .C2(new_n727), .ZN(new_n893));
  OAI221_X1 g0693(.A(new_n373), .B1(new_n474), .B2(new_n697), .C1(new_n722), .C2(new_n275), .ZN(new_n894));
  INV_X1    g0694(.A(G317), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n715), .A2(new_n548), .B1(new_n702), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(G311), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n707), .A2(new_n897), .B1(new_n725), .B2(new_n700), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n894), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n726), .A2(G97), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n783), .A2(new_n282), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n899), .B(new_n900), .C1(new_n901), .C2(KEYINPUT46), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n901), .A2(KEYINPUT46), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n893), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT47), .Z(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(new_n695), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n587), .A2(new_n638), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n585), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n605), .B2(new_n908), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n884), .B(new_n906), .C1(new_n745), .C2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT44), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n522), .A2(new_n623), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n526), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n609), .B2(new_n638), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n913), .B1(new_n641), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n916), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n632), .A2(new_n639), .ZN(new_n919));
  OAI211_X1 g0719(.A(KEYINPUT44), .B(new_n918), .C1(new_n919), .C2(new_n635), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n922));
  NAND3_X1  g0722(.A1(new_n641), .A2(new_n916), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n641), .A2(new_n916), .ZN(new_n924));
  INV_X1    g0724(.A(new_n922), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n921), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n633), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n637), .A2(new_n640), .ZN(new_n929));
  OR3_X1    g0729(.A1(new_n929), .A2(new_n919), .A3(new_n626), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n626), .B1(new_n929), .B2(new_n919), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n932), .A2(new_n686), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n921), .A2(new_n634), .A3(new_n923), .A4(new_n926), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n928), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT107), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT107), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n928), .A2(new_n934), .A3(new_n937), .A4(new_n933), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n687), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n644), .B(KEYINPUT41), .Z(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n691), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n634), .A2(new_n918), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT43), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n910), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n526), .A2(new_n627), .A3(new_n914), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n623), .B1(new_n948), .B2(new_n609), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n637), .A2(new_n640), .A3(new_n916), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(KEYINPUT42), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT42), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n919), .A2(new_n952), .A3(new_n916), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n947), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT105), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n910), .A2(new_n946), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT102), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n955), .B1(new_n954), .B2(new_n958), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT103), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n951), .A2(new_n953), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n957), .C1(new_n964), .C2(new_n947), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT103), .B1(new_n954), .B2(new_n958), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT104), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n962), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n965), .A2(new_n966), .ZN(new_n970));
  INV_X1    g0770(.A(new_n961), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n959), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT104), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n945), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n968), .B1(new_n962), .B2(new_n967), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n970), .A2(new_n972), .A3(KEYINPUT104), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n976), .A3(new_n944), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n912), .B1(new_n943), .B2(new_n978), .ZN(G387));
  OR3_X1    g0779(.A1(new_n239), .A2(new_n253), .A3(new_n276), .ZN(new_n980));
  OAI21_X1  g0780(.A(KEYINPUT50), .B1(new_n319), .B2(G50), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n981), .B(new_n253), .C1(new_n218), .C2(new_n339), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n319), .A2(KEYINPUT50), .A3(G50), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n373), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n646), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n643), .B1(new_n980), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n746), .B1(new_n474), .B2(new_n214), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G322), .A2(new_n706), .B1(new_n721), .B2(G317), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n275), .B2(new_n700), .C1(new_n897), .C2(new_n715), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT48), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n725), .B2(new_n697), .C1(new_n548), .C2(new_n783), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT111), .Z(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT49), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n373), .B1(new_n705), .B2(new_n702), .C1(new_n727), .C2(new_n282), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n992), .B2(KEYINPUT49), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n373), .B1(new_n703), .B2(G150), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n900), .B(new_n996), .C1(new_n783), .C2(new_n339), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT110), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n697), .A2(new_n481), .B1(new_n700), .B2(new_n218), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n722), .A2(new_n202), .B1(new_n319), .B2(new_n715), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(G159), .C2(new_n706), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n993), .A2(new_n995), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n692), .B1(new_n986), .B2(new_n987), .C1(new_n1002), .C2(new_n695), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n632), .B2(new_n745), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n932), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1004), .B1(new_n691), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n933), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n644), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1005), .A2(new_n687), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(G393));
  NAND2_X1  g0810(.A1(new_n918), .A2(new_n745), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT112), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n247), .A2(new_n750), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n746), .B1(new_n285), .B2(new_n214), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n692), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n712), .A2(G283), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G317), .A2(new_n706), .B1(new_n721), .B2(G311), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT52), .Z(new_n1018));
  OAI22_X1  g0818(.A1(new_n702), .A2(new_n720), .B1(new_n700), .B2(new_n548), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n373), .B1(new_n697), .B2(new_n282), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(G303), .C2(new_n716), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n735), .A2(new_n1016), .A3(new_n1018), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(G150), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n707), .A2(new_n1023), .B1(new_n722), .B2(new_n737), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT51), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n276), .B1(new_n697), .B2(new_n339), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n715), .A2(new_n202), .B1(new_n700), .B2(new_n319), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n712), .A2(G68), .B1(G143), .B2(new_n703), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n773), .B(new_n1030), .C1(new_n1032), .C2(KEYINPUT113), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1032), .A2(KEYINPUT113), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1022), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1015), .B1(new_n1035), .B2(new_n694), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1012), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n928), .A2(new_n934), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1037), .B1(new_n1038), .B2(new_n690), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n645), .B1(new_n1038), .B2(new_n1007), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1039), .B1(new_n939), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(G390));
  OAI21_X1  g0842(.A(new_n276), .B1(new_n727), .B2(new_n202), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1043), .A2(KEYINPUT116), .ZN(new_n1044));
  INV_X1    g0844(.A(G128), .ZN(new_n1045));
  INV_X1    g0845(.A(G125), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n707), .A2(new_n1045), .B1(new_n1046), .B2(new_n702), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n722), .A2(new_n775), .B1(new_n715), .B2(new_n890), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(KEYINPUT54), .B(G143), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n697), .A2(new_n737), .B1(new_n700), .B2(new_n1049), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1043), .A2(KEYINPUT116), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n712), .A2(G150), .ZN(new_n1053));
  XOR2_X1   g0853(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1054));
  XNOR2_X1  g0854(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1044), .A2(new_n1051), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n373), .B1(new_n339), .B2(new_n697), .C1(new_n722), .C2(new_n282), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n715), .A2(new_n474), .B1(new_n702), .B2(new_n548), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n707), .A2(new_n725), .B1(new_n285), .B2(new_n700), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n734), .B(new_n1060), .C1(new_n727), .C2(new_n218), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n695), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n693), .B(new_n1062), .C1(new_n319), .C2(new_n787), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n865), .A2(new_n866), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1063), .B1(new_n1065), .B2(new_n744), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n796), .A2(new_n807), .A3(G330), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n638), .B(new_n761), .C1(new_n679), .C2(new_n680), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n857), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n807), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n867), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n839), .A2(new_n840), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n856), .A2(new_n857), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n807), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n865), .A2(new_n866), .B1(new_n1076), .B2(new_n1072), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1068), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1072), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1064), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n672), .A2(G330), .A3(new_n761), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1081), .A2(new_n842), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1078), .A2(new_n1085), .A3(KEYINPUT114), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT114), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n1088), .A3(new_n1068), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n807), .B1(new_n796), .B2(G330), .ZN(new_n1091));
  OR3_X1    g0891(.A1(new_n1091), .A2(new_n1082), .A3(new_n1070), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1081), .A2(new_n842), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1067), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1075), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n493), .A2(G330), .A3(new_n795), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1096), .A2(new_n602), .A3(new_n853), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n644), .B1(new_n1090), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1066), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT115), .B1(new_n1090), .B2(new_n691), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT115), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1104), .B(new_n690), .C1(new_n1086), .C2(new_n1089), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1102), .A2(new_n1106), .ZN(G378));
  NAND2_X1  g0907(.A1(new_n359), .A2(new_n810), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n358), .A2(new_n362), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n358), .B2(new_n362), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  OR3_X1    g0912(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1112), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(G330), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n841), .B2(new_n844), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1115), .B1(new_n831), .B2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n828), .B(KEYINPUT40), .C1(new_n862), .C2(new_n844), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT101), .B1(new_n825), .B2(new_n826), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1117), .B(new_n1115), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n869), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1117), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1115), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n869), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n1127), .A3(new_n1121), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1123), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n691), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n693), .B1(new_n202), .B2(new_n787), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n722), .A2(new_n1045), .B1(new_n775), .B2(new_n715), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n701), .A2(G137), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n1023), .B2(new_n697), .C1(new_n1046), .C2(new_n707), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1049), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1132), .B(new_n1134), .C1(new_n712), .C2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT59), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n726), .A2(G159), .ZN(new_n1140));
  AOI211_X1 g0940(.A(G33), .B(G41), .C1(new_n703), .C2(G124), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n783), .A2(new_n339), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n727), .A2(new_n377), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n276), .A2(G41), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n218), .B2(new_n697), .C1(new_n722), .C2(new_n474), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G283), .A2(new_n703), .B1(new_n706), .B2(G116), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n285), .B2(new_n715), .C1(new_n481), .C2(new_n700), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1149), .A2(KEYINPUT58), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(KEYINPUT58), .ZN(new_n1151));
  AOI211_X1 g0951(.A(G50), .B(new_n1145), .C1(new_n268), .C2(new_n256), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT118), .Z(new_n1153));
  AND4_X1   g0953(.A1(new_n1142), .A2(new_n1150), .A3(new_n1151), .A4(new_n1153), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1131), .B1(new_n695), .B2(new_n1154), .C1(new_n1115), .C2(new_n744), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1130), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n853), .A2(new_n602), .A3(new_n1097), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT119), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(KEYINPUT114), .B(new_n1067), .C1(new_n1080), .C2(new_n1084), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1088), .B1(new_n1087), .B2(new_n1068), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n1085), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1160), .B1(new_n1163), .B2(new_n1098), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1129), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1126), .A2(new_n1127), .A3(new_n1121), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1127), .B1(new_n1126), .B2(new_n1121), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT57), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1159), .B1(new_n1090), .B2(new_n1099), .ZN(new_n1171));
  OAI211_X1 g0971(.A(KEYINPUT120), .B(new_n644), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1166), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n1164), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT120), .B1(new_n1175), .B2(new_n644), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1157), .B1(new_n1173), .B2(new_n1176), .ZN(G375));
  NAND2_X1  g0977(.A1(new_n1096), .A2(new_n691), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n373), .B1(new_n481), .B2(new_n697), .C1(new_n722), .C2(new_n725), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n702), .A2(new_n275), .B1(new_n700), .B2(new_n474), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n707), .A2(new_n548), .B1(new_n282), .B2(new_n715), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n783), .B2(new_n285), .C1(new_n339), .C2(new_n727), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1144), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n702), .A2(new_n1045), .B1(new_n700), .B2(new_n1023), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n716), .B2(new_n1135), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT121), .B1(new_n707), .B2(new_n775), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n707), .A2(KEYINPUT121), .A3(new_n775), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n276), .B1(new_n722), .B2(new_n890), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n697), .A2(new_n202), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .A4(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n783), .A2(new_n737), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1183), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n695), .B1(new_n1194), .B2(KEYINPUT122), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(KEYINPUT122), .B2(new_n1194), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n693), .B1(new_n218), .B2(new_n787), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n807), .C2(new_n744), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1178), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT123), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1199), .B(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1096), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1158), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n942), .A3(new_n1098), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1204), .ZN(G381));
  OR2_X1    g1005(.A1(G393), .A2(G396), .ZN(new_n1206));
  OR4_X1    g1006(.A1(G384), .A2(G381), .A3(new_n1206), .A4(G390), .ZN(new_n1207));
  OR4_X1    g1007(.A1(G387), .A2(new_n1207), .A3(G375), .A4(G378), .ZN(G407));
  NOR2_X1   g1008(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n622), .A2(G213), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT124), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(G407), .B(G213), .C1(G375), .C2(new_n1212), .ZN(G409));
  OAI211_X1 g1013(.A(G378), .B(new_n1157), .C1(new_n1173), .C2(new_n1176), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1165), .A2(new_n941), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1209), .B1(new_n1215), .B2(new_n1156), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1210), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1098), .A2(KEYINPUT60), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1203), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1202), .A2(KEYINPUT60), .A3(new_n1158), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(new_n644), .A3(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1222), .A2(new_n1201), .A3(G384), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G384), .B1(new_n1222), .B2(new_n1201), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n622), .A2(G213), .A3(G2897), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT125), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1222), .A2(new_n1201), .ZN(new_n1228));
  INV_X1    g1028(.A(G384), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1222), .A2(new_n1201), .A3(G384), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(G2897), .A3(new_n1211), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1227), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT125), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1211), .A2(G2897), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1218), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT126), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G387), .B2(new_n1041), .ZN(new_n1240));
  XOR2_X1   g1040(.A(G393), .B(G396), .Z(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n975), .A2(new_n976), .A3(new_n944), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n944), .B1(new_n975), .B2(new_n976), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n686), .B1(new_n936), .B2(new_n938), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n690), .B1(new_n1246), .B2(new_n941), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n911), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(G390), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n911), .B(new_n1041), .C1(new_n1245), .C2(new_n1247), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n1240), .A2(new_n1242), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G387), .A2(new_n1041), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(G390), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1239), .A4(new_n1241), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1251), .A2(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(KEYINPUT61), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1217), .A2(new_n1210), .A3(new_n1225), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT63), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1211), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1225), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1238), .A2(new_n1256), .A3(new_n1259), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1237), .B1(new_n1227), .B2(new_n1233), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n1260), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT62), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1257), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1260), .A2(KEYINPUT62), .A3(new_n1225), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1265), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1255), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1262), .B1(new_n1269), .B2(new_n1270), .ZN(G405));
  INV_X1    g1071(.A(new_n1214), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n644), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT120), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1167), .A3(new_n1172), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G378), .B1(new_n1276), .B2(new_n1157), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1225), .B1(new_n1272), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G375), .A2(new_n1209), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(new_n1232), .A3(new_n1214), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1255), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1255), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  AOI211_X1 g1084(.A(KEYINPUT127), .B(new_n1255), .C1(new_n1278), .C2(new_n1280), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(G402));
endmodule


