//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1223, new_n1224, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n462), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n466), .A2(new_n474), .ZN(G160));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n471), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n477), .B2(new_n467), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n462), .B1(new_n477), .B2(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G138), .B(new_n462), .C1(new_n468), .C2(new_n469), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n463), .A2(new_n488), .A3(G138), .A4(new_n462), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n462), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT68), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n494), .A2(new_n496), .A3(new_n497), .A4(G2104), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n493), .A2(new_n498), .B1(new_n480), .B2(G126), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n490), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n503), .A2(KEYINPUT69), .A3(G50), .A4(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT70), .B1(new_n509), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT71), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(new_n509), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n514), .A2(new_n518), .A3(new_n503), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G88), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n514), .A2(new_n518), .A3(G62), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n508), .B(new_n520), .C1(new_n524), .C2(KEYINPUT72), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(KEYINPUT72), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(G166));
  AND2_X1   g102(.A1(new_n514), .A2(new_n518), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(new_n504), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n530), .A2(G51), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n519), .A2(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n540));
  OAI21_X1  g115(.A(G651), .B1(new_n539), .B2(KEYINPUT73), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n530), .A2(G52), .ZN(new_n543));
  INV_X1    g118(.A(new_n519), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT74), .B(G90), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n530), .A2(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n528), .A2(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n521), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n530), .A2(new_n561), .A3(KEYINPUT9), .A4(G53), .ZN(new_n562));
  XNOR2_X1  g137(.A(KEYINPUT76), .B(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n504), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n514), .A2(new_n518), .ZN(new_n568));
  XOR2_X1   g143(.A(KEYINPUT78), .B(G65), .Z(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n566), .B1(new_n570), .B2(G651), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n544), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n519), .A2(KEYINPUT77), .A3(G91), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n571), .A2(new_n576), .ZN(G299));
  OR2_X1    g152(.A1(new_n542), .A2(new_n546), .ZN(G301));
  OR2_X1    g153(.A1(new_n524), .A2(KEYINPUT72), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n524), .A2(KEYINPUT72), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n506), .A2(new_n507), .B1(new_n519), .B2(G88), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G303));
  NAND2_X1  g157(.A1(new_n530), .A2(G49), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n514), .A2(new_n518), .A3(G87), .A4(new_n503), .ZN(new_n584));
  AOI21_X1  g159(.A(G74), .B1(new_n514), .B2(new_n518), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n521), .C2(new_n585), .ZN(G288));
  NAND3_X1  g161(.A1(new_n514), .A2(new_n518), .A3(G61), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n521), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n514), .A2(new_n518), .A3(G86), .A4(new_n503), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n503), .A2(G48), .A3(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n590), .A2(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n521), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n530), .A2(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n544), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(new_n519), .A2(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n568), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G171), .B2(new_n611), .ZN(G284));
  OAI21_X1  g188(.A(new_n612), .B1(G171), .B2(new_n611), .ZN(G321));
  NAND2_X1  g189(.A1(G299), .A2(new_n611), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n611), .B2(G168), .ZN(G280));
  XOR2_X1   g191(.A(G280), .B(KEYINPUT79), .Z(G297));
  INV_X1    g192(.A(new_n610), .ZN(new_n618));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n463), .A2(new_n472), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT13), .Z(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n478), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n480), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n462), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(G2096), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n629), .A2(new_n630), .A3(new_n637), .ZN(G156));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT80), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n643), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT81), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(G401));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT82), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n636), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n676), .A2(new_n679), .A3(new_n683), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1991), .B(G1996), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n686), .B(new_n687), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(new_n690), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n674), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n690), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n689), .A2(new_n691), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n696), .A2(new_n697), .A3(new_n673), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  MUX2_X1   g275(.A(G23), .B(G288), .S(G16), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT87), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT33), .B(G1976), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(G166), .A2(G16), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G16), .B2(G22), .ZN(new_n706));
  INV_X1    g281(.A(G1971), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(G6), .B(G305), .S(G16), .Z(new_n709));
  XOR2_X1   g284(.A(KEYINPUT32), .B(G1981), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n706), .A2(new_n707), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n704), .A2(new_n708), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT86), .B(KEYINPUT34), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n713), .A2(new_n715), .ZN(new_n717));
  NOR2_X1   g292(.A1(G16), .A2(G24), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n601), .B2(G16), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1986), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n721), .A2(G25), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n480), .A2(G119), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n726));
  INV_X1    g301(.A(G107), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(G2105), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n478), .B2(G131), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n722), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT85), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n731), .A2(new_n733), .B1(KEYINPUT89), .B2(KEYINPUT36), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n731), .B2(new_n733), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n720), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n716), .A2(new_n717), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(KEYINPUT89), .B1(KEYINPUT88), .B2(KEYINPUT36), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G16), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n740), .A2(G21), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G286), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1966), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT97), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT30), .B(G28), .ZN(new_n746));
  OR2_X1    g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  NAND2_X1  g322(.A1(KEYINPUT31), .A2(G11), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n746), .A2(new_n721), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n635), .B2(new_n721), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n742), .B2(new_n743), .ZN(new_n751));
  INV_X1    g326(.A(G1961), .ZN(new_n752));
  NOR2_X1   g327(.A1(G171), .A2(new_n740), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G5), .B2(new_n740), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n745), .B(new_n751), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT98), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n721), .A2(G32), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n472), .A2(G105), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT95), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n480), .A2(G129), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n478), .A2(G141), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n759), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT96), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n757), .B1(new_n769), .B2(new_n721), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT27), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1996), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT25), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n463), .A2(G127), .ZN(new_n775));
  NAND2_X1  g350(.A1(G115), .A2(G2104), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n462), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n774), .B(new_n777), .C1(G139), .C2(new_n478), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(new_n721), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n721), .B2(G33), .ZN(new_n780));
  INV_X1    g355(.A(G2072), .ZN(new_n781));
  INV_X1    g356(.A(G2084), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n721), .B1(KEYINPUT24), .B2(G34), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(KEYINPUT24), .B2(G34), .ZN(new_n784));
  INV_X1    g359(.A(G160), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(G29), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n780), .A2(new_n781), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n721), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n721), .ZN(new_n789));
  INV_X1    g364(.A(G2078), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n787), .B(new_n791), .C1(new_n781), .C2(new_n780), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n721), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n721), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT29), .B(G2090), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n786), .A2(new_n782), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT94), .Z(new_n798));
  NOR3_X1   g373(.A1(new_n792), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n754), .A2(new_n752), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT99), .B(KEYINPUT23), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n740), .A2(G20), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G299), .B2(G16), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT100), .B(G1956), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n772), .A2(new_n799), .A3(new_n800), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n740), .A2(G4), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n618), .B2(new_n740), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT90), .B(G1348), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n721), .A2(G26), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT28), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n478), .A2(G140), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n480), .A2(G128), .ZN(new_n815));
  OR2_X1    g390(.A1(G104), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(new_n721), .ZN(new_n820));
  INV_X1    g395(.A(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n740), .A2(G19), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT91), .Z(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n554), .B2(new_n740), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT92), .B(G1341), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n811), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT93), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n756), .A2(new_n807), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n737), .A2(new_n738), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n739), .A2(new_n830), .A3(new_n831), .ZN(G150));
  INV_X1    g407(.A(G150), .ZN(G311));
  AOI22_X1  g408(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(new_n521), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n530), .A2(G55), .ZN(new_n836));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n544), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G860), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n610), .A2(new_n619), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT102), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n843), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n839), .A2(new_n554), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n835), .A2(new_n838), .B1(new_n550), .B2(new_n553), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n846), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT103), .B1(new_n850), .B2(new_n851), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n850), .B2(new_n851), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n842), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT104), .Z(G145));
  XOR2_X1   g434(.A(G160), .B(new_n635), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n484), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n730), .B(KEYINPUT106), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n626), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n730), .B(KEYINPUT106), .ZN(new_n864));
  INV_X1    g439(.A(new_n626), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n493), .A2(new_n498), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n463), .A2(G126), .A3(G2105), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n492), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n497), .B1(new_n873), .B2(new_n496), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT68), .ZN(new_n875));
  OAI211_X1 g450(.A(KEYINPUT105), .B(new_n869), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n490), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n778), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n867), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n769), .A2(new_n819), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n768), .A2(new_n818), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n478), .A2(G142), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n480), .A2(G130), .ZN(new_n884));
  OR2_X1    g459(.A1(G106), .A2(G2105), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n885), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n880), .A2(new_n887), .A3(new_n881), .ZN(new_n890));
  INV_X1    g465(.A(new_n878), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n863), .A2(new_n866), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n879), .A2(new_n889), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n879), .A2(new_n892), .B1(new_n889), .B2(new_n890), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n861), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  INV_X1    g472(.A(new_n861), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n893), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(G395));
  INV_X1    g478(.A(KEYINPUT110), .ZN(new_n904));
  XNOR2_X1  g479(.A(G166), .B(new_n601), .ZN(new_n905));
  XNOR2_X1  g480(.A(G305), .B(G288), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT42), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n621), .B(new_n849), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(G299), .A2(KEYINPUT108), .ZN(new_n912));
  NAND2_X1  g487(.A1(G299), .A2(KEYINPUT108), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n618), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n610), .A2(G299), .A3(KEYINPUT108), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n914), .B2(new_n916), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n911), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n914), .A2(new_n916), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n911), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n909), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n920), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n908), .B1(new_n925), .B2(new_n922), .ZN(new_n926));
  AND4_X1   g501(.A1(new_n904), .A2(new_n924), .A3(G868), .A4(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n904), .B1(new_n840), .B2(new_n611), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n925), .A2(new_n922), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n611), .B1(new_n930), .B2(new_n909), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n929), .B1(new_n931), .B2(new_n926), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT111), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n924), .A2(G868), .ZN(new_n934));
  INV_X1    g509(.A(new_n926), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n928), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n931), .A2(new_n904), .A3(new_n926), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n933), .A2(new_n939), .ZN(G295));
  NOR2_X1   g515(.A1(new_n927), .A2(new_n932), .ZN(G331));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n943));
  NAND3_X1  g518(.A1(G301), .A2(new_n848), .A3(new_n847), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n849), .A2(G171), .ZN(new_n945));
  AOI21_X1  g520(.A(G168), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(G168), .A3(new_n945), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n947), .B(new_n948), .C1(new_n917), .C2(new_n919), .ZN(new_n949));
  INV_X1    g524(.A(new_n921), .ZN(new_n950));
  INV_X1    g525(.A(new_n948), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(new_n951), .B2(new_n946), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n952), .A3(new_n907), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n900), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n921), .A2(new_n915), .ZN(new_n955));
  INV_X1    g530(.A(new_n918), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n914), .A2(new_n956), .A3(new_n916), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n955), .A2(new_n947), .A3(new_n948), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n907), .B1(new_n958), .B2(new_n952), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n943), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n952), .ZN(new_n961));
  INV_X1    g536(.A(new_n907), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n963), .A2(KEYINPUT112), .A3(new_n900), .A4(new_n953), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n942), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n907), .B1(new_n949), .B2(new_n952), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n954), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT44), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n954), .B2(new_n966), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n963), .A2(new_n942), .A3(new_n900), .A4(new_n953), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(G397));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n876), .A2(new_n490), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT105), .B1(new_n868), .B2(new_n869), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G40), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n466), .A2(new_n982), .A3(new_n474), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n768), .B(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n818), .B(new_n821), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n730), .B(new_n732), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n601), .B(G1986), .Z(new_n991));
  OAI21_X1  g566(.A(new_n985), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(KEYINPUT55), .B(G8), .C1(new_n525), .C2(new_n526), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(G166), .B2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(G303), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(G8), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n995), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n877), .B2(new_n976), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT117), .B1(new_n1002), .B2(new_n984), .ZN(new_n1003));
  INV_X1    g578(.A(G2090), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n500), .A2(new_n976), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n499), .A2(KEYINPUT105), .B1(new_n487), .B2(new_n489), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1384), .B1(new_n1009), .B2(new_n872), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1008), .B(new_n983), .C1(new_n1010), .C2(new_n1001), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1003), .A2(new_n1004), .A3(new_n1007), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1005), .A2(new_n980), .ZN(new_n1013));
  OAI211_X1 g588(.A(KEYINPUT45), .B(new_n976), .C1(new_n977), .C2(new_n978), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n983), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n707), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1000), .B1(new_n1017), .B2(G8), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT50), .B1(new_n877), .B2(new_n976), .ZN(new_n1019));
  AOI211_X1 g594(.A(new_n1001), .B(G1384), .C1(new_n490), .C2(new_n499), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n983), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1016), .B1(new_n1021), .B2(G2090), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(new_n1000), .A3(G8), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n997), .B1(new_n1010), .B2(new_n983), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n583), .A2(new_n584), .ZN(new_n1025));
  OAI21_X1  g600(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(KEYINPUT115), .A3(G1976), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(G288), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1024), .A2(new_n1027), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n589), .A2(new_n593), .A3(G1981), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(G1981), .B1(new_n589), .B2(new_n593), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(KEYINPUT49), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1035), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(new_n1033), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1024), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n983), .B(new_n976), .C1(new_n977), .C2(new_n978), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1030), .A2(new_n1041), .A3(new_n1027), .A4(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1032), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1023), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1018), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT45), .B1(new_n877), .B2(new_n976), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n983), .B1(new_n1005), .B2(new_n980), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(G2078), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1021), .A2(new_n752), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1013), .A2(new_n1014), .A3(new_n790), .A4(new_n983), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT124), .B1(new_n1053), .B2(new_n1050), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(KEYINPUT124), .A3(new_n1050), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1052), .B(G301), .C1(new_n1054), .C2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1020), .B1(new_n979), .B2(new_n1001), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n752), .B1(new_n1058), .B2(new_n984), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n474), .A2(KEYINPUT126), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n474), .A2(KEYINPUT126), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1051), .A2(G40), .ZN(new_n1062));
  NOR4_X1   g637(.A1(new_n1060), .A2(new_n1061), .A3(new_n466), .A4(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n981), .A2(new_n1014), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1054), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(new_n1055), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1057), .B(KEYINPUT54), .C1(new_n1067), .C2(G301), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1046), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT125), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n1059), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n1066), .B2(new_n1055), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1071), .B1(new_n1074), .B2(G301), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1052), .B1(new_n1056), .B2(new_n1054), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1067), .A2(G301), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1069), .B1(new_n1070), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(G168), .A2(new_n997), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(G1384), .B1(new_n490), .B2(new_n499), .ZN(new_n1083));
  INV_X1    g658(.A(new_n980), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n984), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT45), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n979), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1966), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n983), .A2(new_n782), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n979), .A2(new_n1001), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1020), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT122), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n743), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1089), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1082), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1088), .A2(new_n1092), .A3(KEYINPUT122), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1097), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1103));
  OAI21_X1  g678(.A(G8), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1081), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1105), .B(new_n997), .C1(new_n1093), .C2(new_n1098), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1101), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(G8), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(new_n1101), .A3(new_n1082), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1100), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1956), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1011), .A2(new_n1007), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n984), .B1(new_n979), .B2(KEYINPUT50), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n1008), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1114), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1121), .B(new_n1122), .C1(new_n571), .C2(new_n576), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n571), .A2(new_n1119), .A3(new_n576), .A4(new_n1120), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1015), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT56), .B(G2072), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1118), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT119), .B1(new_n1041), .B2(G2067), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1010), .A2(new_n1132), .A3(new_n821), .A4(new_n983), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n810), .B1(new_n1058), .B2(new_n984), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n610), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1130), .A2(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1006), .B1(new_n1116), .B2(new_n1008), .ZN(new_n1139));
  AOI21_X1  g714(.A(G1956), .B1(new_n1139), .B2(new_n1003), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1129), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1138), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n810), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1091), .B1(new_n1010), .B2(KEYINPUT50), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(new_n983), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1146), .A2(new_n1147), .A3(new_n618), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT60), .B1(new_n1148), .B2(new_n1136), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1013), .A2(new_n1014), .A3(new_n986), .A4(new_n983), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT58), .B(G1341), .Z(new_n1151));
  NAND2_X1  g726(.A1(new_n1041), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n554), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1153), .A2(new_n1156), .A3(new_n554), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n610), .A2(KEYINPUT60), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1155), .A2(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1149), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT61), .B1(new_n1142), .B2(new_n1130), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1126), .B1(new_n1118), .B2(new_n1129), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1130), .B1(new_n1164), .B2(KEYINPUT120), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1118), .A2(new_n1166), .A3(new_n1126), .A4(new_n1129), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1165), .A2(KEYINPUT61), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1143), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1080), .B(new_n1113), .C1(new_n1169), .C2(KEYINPUT121), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1169), .A2(KEYINPUT121), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1044), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1024), .ZN(new_n1174));
  NOR2_X1   g749(.A1(G288), .A2(G1976), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT116), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1033), .B1(new_n1040), .B2(new_n1176), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1173), .A2(new_n1023), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1046), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1110), .A2(G286), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1000), .B1(new_n1022), .B2(G8), .ZN(new_n1183));
  OR4_X1    g758(.A1(new_n1179), .A2(new_n1045), .A3(new_n1181), .A4(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1178), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1180), .B1(new_n1077), .B2(new_n1075), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n997), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1082), .B1(new_n1187), .B2(KEYINPUT123), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT51), .B1(new_n1188), .B2(new_n1107), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1099), .B1(new_n1189), .B2(new_n1111), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1186), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI211_X1 g767(.A(KEYINPUT62), .B(new_n1099), .C1(new_n1189), .C2(new_n1111), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1185), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n992), .B1(new_n1172), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n987), .A2(new_n988), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n725), .A2(new_n729), .A3(new_n732), .ZN(new_n1197));
  OAI22_X1  g772(.A1(new_n1196), .A2(new_n1197), .B1(G2067), .B2(new_n818), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1198), .A2(new_n985), .ZN(new_n1199));
  INV_X1    g774(.A(new_n988), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n985), .B1(new_n768), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n985), .A2(new_n986), .ZN(new_n1202));
  AND2_X1   g777(.A1(new_n1202), .A2(KEYINPUT46), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1202), .A2(KEYINPUT46), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  XOR2_X1   g780(.A(new_n1205), .B(KEYINPUT47), .Z(new_n1206));
  INV_X1    g781(.A(G1986), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n985), .A2(new_n1207), .A3(new_n601), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT48), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1211), .B1(new_n990), .B2(new_n985), .ZN(new_n1212));
  AOI211_X1 g787(.A(new_n1199), .B(new_n1206), .C1(new_n1210), .C2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1195), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n1216));
  OR2_X1    g790(.A1(G227), .A2(new_n460), .ZN(new_n1217));
  AOI21_X1  g791(.A(new_n1217), .B1(new_n657), .B2(new_n658), .ZN(new_n1218));
  AND3_X1   g792(.A1(new_n901), .A2(new_n699), .A3(new_n1218), .ZN(new_n1219));
  AND3_X1   g793(.A1(new_n972), .A2(new_n1216), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g794(.A(new_n1216), .B1(new_n972), .B2(new_n1219), .ZN(new_n1221));
  NOR2_X1   g795(.A1(new_n1220), .A2(new_n1221), .ZN(G308));
  NAND2_X1  g796(.A1(new_n972), .A2(new_n1219), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n1223), .A2(KEYINPUT127), .ZN(new_n1224));
  NAND3_X1  g798(.A1(new_n972), .A2(new_n1219), .A3(new_n1216), .ZN(new_n1225));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n1225), .ZN(G225));
endmodule


