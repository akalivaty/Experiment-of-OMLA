//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G952), .ZN(new_n189));
  AOI211_X1 g003(.A(G953), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT21), .B(G898), .Z(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT96), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G902), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  AOI211_X1 g009(.A(new_n194), .B(new_n195), .C1(G234), .C2(G237), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n190), .B1(new_n193), .B2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G110), .B(G122), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(new_n200), .B2(G107), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT80), .A3(G101), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n201), .A2(new_n204), .A3(new_n208), .A4(new_n205), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n206), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(G101), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT71), .A2(G119), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT71), .A2(G119), .ZN(new_n214));
  OAI21_X1  g028(.A(G116), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G116), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g032(.A(KEYINPUT2), .B(G113), .Z(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n215), .A3(new_n217), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n211), .A2(new_n212), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n215), .A2(KEYINPUT5), .A3(new_n217), .ZN(new_n224));
  OR2_X1    g038(.A1(KEYINPUT71), .A2(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT71), .A2(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT5), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G116), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n224), .A2(G113), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n203), .A2(G104), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n200), .A2(G107), .ZN(new_n232));
  OAI21_X1  g046(.A(G101), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n209), .A2(new_n233), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n230), .A2(new_n234), .A3(new_n222), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n199), .B1(new_n223), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n211), .A2(new_n212), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n221), .A2(new_n222), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n230), .A2(new_n234), .A3(new_n222), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(new_n198), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n241), .A3(KEYINPUT6), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT0), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT64), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(KEYINPUT0), .B2(G128), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G146), .ZN(new_n249));
  INV_X1    g063(.A(G146), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n245), .B(new_n247), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n250), .A2(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n248), .A2(G146), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G125), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n248), .B(G146), .C1(new_n244), .C2(KEYINPUT1), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n244), .A2(new_n250), .A3(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n255), .A2(new_n256), .A3(new_n266), .A4(G128), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n261), .A2(KEYINPUT69), .A3(new_n262), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G125), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n260), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n195), .A2(G224), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n260), .A2(new_n271), .A3(G224), .A4(new_n195), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n277), .B(new_n199), .C1(new_n223), .C2(new_n235), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n242), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n273), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(KEYINPUT7), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n260), .A2(new_n271), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n198), .B(KEYINPUT8), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n234), .B1(new_n230), .B2(new_n222), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n235), .B2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n280), .A2(new_n241), .A3(new_n282), .A4(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n279), .A2(new_n194), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G210), .B1(G237), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n279), .A2(new_n194), .A3(new_n288), .A4(new_n286), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n188), .B(new_n197), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n267), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n209), .B(new_n233), .C1(new_n293), .C2(new_n263), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n294), .B1(new_n269), .B2(new_n234), .ZN(new_n295));
  AND2_X1   g109(.A1(KEYINPUT67), .A2(G137), .ZN(new_n296));
  NOR2_X1   g110(.A1(KEYINPUT67), .A2(G137), .ZN(new_n297));
  OAI211_X1 g111(.A(KEYINPUT11), .B(G134), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G137), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G134), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT11), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT66), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT11), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G134), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G137), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n298), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G131), .ZN(new_n309));
  INV_X1    g123(.A(G131), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n298), .A2(new_n305), .A3(new_n310), .A4(new_n307), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n295), .A2(new_n312), .A3(KEYINPUT12), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT81), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n295), .A2(new_n312), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT12), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT81), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n295), .A2(new_n312), .A3(new_n318), .A4(KEYINPUT12), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n314), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n237), .A2(new_n259), .ZN(new_n321));
  INV_X1    g135(.A(new_n312), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT10), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n294), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n269), .A2(KEYINPUT10), .A3(new_n234), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n321), .A2(new_n322), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n195), .A2(G227), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT79), .ZN(new_n329));
  INV_X1    g143(.A(G110), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(G140), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n332), .A2(new_n326), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n321), .A2(new_n324), .A3(new_n325), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n312), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n332), .B1(new_n320), .B2(new_n326), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n338), .A2(new_n326), .A3(new_n332), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT82), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(G469), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G469), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(new_n194), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n336), .A2(new_n320), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n269), .A2(new_n234), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n348), .A2(KEYINPUT10), .B1(new_n237), .B2(new_n259), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n322), .B1(new_n349), .B2(new_n324), .ZN(new_n350));
  INV_X1    g164(.A(new_n326), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n333), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(G902), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n346), .B1(new_n353), .B2(new_n345), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n344), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT84), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n248), .ZN(new_n357));
  NOR2_X1   g171(.A1(G237), .A2(G953), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(G214), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G237), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n195), .A3(G214), .ZN(new_n361));
  NOR2_X1   g175(.A1(KEYINPUT84), .A2(G143), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G131), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT17), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n362), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n357), .A2(G214), .A3(new_n358), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(new_n310), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n364), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n270), .A2(G140), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT16), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n374));
  INV_X1    g188(.A(G140), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n374), .B1(new_n375), .B2(G125), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n270), .A2(KEYINPUT74), .A3(G140), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n370), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n373), .B1(new_n378), .B2(new_n372), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G146), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n250), .B(new_n373), .C1(new_n378), .C2(new_n372), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n310), .B1(new_n366), .B2(new_n367), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT17), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n369), .A2(new_n380), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n270), .A2(G140), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n371), .A2(new_n385), .A3(new_n250), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n378), .B2(new_n250), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT18), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n366), .B(new_n367), .C1(new_n388), .C2(new_n310), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n387), .B(new_n389), .C1(new_n364), .C2(new_n388), .ZN(new_n390));
  OR2_X1    g204(.A1(G113), .A2(G122), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT86), .ZN(new_n392));
  NAND2_X1  g206(.A1(G113), .A2(G122), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(G113), .A2(G122), .ZN(new_n395));
  NOR2_X1   g209(.A1(G113), .A2(G122), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT86), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n394), .A2(new_n397), .A3(G104), .ZN(new_n398));
  AOI21_X1  g212(.A(G104), .B1(new_n394), .B2(new_n397), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT87), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n394), .A2(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n200), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT87), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n394), .A2(new_n397), .A3(G104), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n384), .A2(new_n390), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n398), .A2(new_n399), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n384), .B2(new_n390), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n194), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT90), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT89), .B(G475), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n413), .B(new_n194), .C1(new_n407), .C2(new_n409), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(G475), .A2(G902), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT85), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n366), .A2(new_n367), .A3(new_n310), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n418), .B2(new_n382), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n364), .A2(KEYINPUT85), .A3(new_n368), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT19), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n371), .A2(new_n385), .A3(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n422), .B(new_n250), .C1(new_n378), .C2(new_n421), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n419), .A2(new_n420), .A3(new_n380), .A4(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n408), .B1(new_n424), .B2(new_n390), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n416), .B1(new_n407), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n416), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT20), .B1(new_n429), .B2(KEYINPUT88), .ZN(new_n430));
  OAI221_X1 g244(.A(new_n430), .B1(KEYINPUT88), .B2(new_n429), .C1(new_n407), .C2(new_n425), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n415), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n248), .A2(G128), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n244), .A2(G143), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT91), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT91), .B1(new_n434), .B2(new_n435), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n436), .A2(new_n437), .A3(new_n306), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n244), .A2(G143), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n248), .A2(G128), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT91), .ZN(new_n443));
  AOI21_X1  g257(.A(G134), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT92), .B1(new_n438), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n306), .B1(new_n436), .B2(new_n437), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n442), .A2(G134), .A3(new_n443), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n216), .A2(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT14), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT94), .ZN(new_n452));
  INV_X1    g266(.A(G122), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G116), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT94), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(new_n455), .A3(KEYINPUT14), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n450), .A2(KEYINPUT14), .ZN(new_n458));
  OAI21_X1  g272(.A(G107), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n454), .A2(new_n450), .A3(new_n203), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT93), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n445), .A2(new_n449), .A3(new_n459), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n203), .B1(new_n454), .B2(new_n450), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n454), .A2(new_n450), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G107), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n440), .A2(KEYINPUT13), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n440), .A2(KEYINPUT13), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n466), .A2(new_n467), .A3(new_n441), .ZN(new_n468));
  OAI221_X1 g282(.A(new_n446), .B1(new_n463), .B2(new_n465), .C1(new_n468), .C2(new_n306), .ZN(new_n469));
  XOR2_X1   g283(.A(KEYINPUT9), .B(G234), .Z(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G217), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n471), .A2(new_n472), .A3(G953), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n462), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n462), .B2(new_n469), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n194), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G478), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(KEYINPUT15), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n478), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n194), .B(new_n480), .C1(new_n474), .C2(new_n475), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(KEYINPUT95), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT95), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n462), .A2(new_n469), .ZN(new_n484));
  INV_X1    g298(.A(new_n473), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n462), .A2(new_n469), .A3(new_n473), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n480), .B1(new_n488), .B2(new_n194), .ZN(new_n489));
  INV_X1    g303(.A(new_n481), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n483), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n433), .B1(new_n482), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G221), .B1(new_n471), .B2(G902), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n292), .A2(new_n355), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT97), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT32), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n358), .A2(G210), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n498), .B(KEYINPUT27), .Z(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT26), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(new_n208), .ZN(new_n501));
  OR3_X1    g315(.A1(new_n306), .A2(KEYINPUT68), .A3(G137), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n300), .A2(KEYINPUT68), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n296), .A2(new_n297), .A3(G134), .ZN(new_n505));
  OAI21_X1  g319(.A(G131), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n269), .A2(new_n311), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n309), .A2(new_n311), .B1(new_n254), .B2(new_n258), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n507), .A2(new_n508), .A3(new_n238), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n269), .A2(new_n311), .A3(new_n506), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n269), .A2(new_n506), .A3(new_n514), .A4(new_n311), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT65), .B1(new_n254), .B2(new_n258), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT65), .ZN(new_n518));
  AOI211_X1 g332(.A(new_n518), .B(new_n257), .C1(new_n252), .C2(new_n253), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n312), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n238), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n501), .B1(new_n511), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n507), .A2(new_n508), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n522), .B2(new_n525), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n509), .B1(new_n527), .B2(new_n238), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n528), .A2(KEYINPUT72), .A3(KEYINPUT31), .A4(new_n501), .ZN(new_n529));
  OR3_X1    g343(.A1(new_n507), .A2(new_n508), .A3(new_n525), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n513), .A2(new_n515), .B1(new_n520), .B2(new_n312), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n238), .B(new_n530), .C1(new_n531), .C2(KEYINPUT30), .ZN(new_n532));
  INV_X1    g346(.A(new_n509), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n532), .A2(KEYINPUT72), .A3(new_n533), .A4(new_n501), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n524), .B1(new_n529), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT73), .ZN(new_n538));
  OR3_X1    g352(.A1(new_n538), .A2(G472), .A3(G902), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n538), .B1(G472), .B2(G902), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n497), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n524), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n534), .A2(new_n535), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n534), .A2(new_n535), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(KEYINPUT32), .A3(new_n541), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n511), .A2(new_n523), .A3(new_n501), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n501), .B1(new_n532), .B2(new_n533), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT29), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n238), .B1(new_n507), .B2(new_n508), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n511), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n501), .A2(KEYINPUT29), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n194), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G472), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n543), .A2(new_n548), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n493), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(new_n344), .B2(new_n354), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n559), .A2(new_n292), .A3(KEYINPUT97), .A4(new_n492), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT78), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT22), .B(G137), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n244), .B1(new_n225), .B2(new_n226), .ZN(new_n568));
  INV_X1    g382(.A(G119), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(G128), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT24), .B(G110), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT23), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n573), .A2(new_n569), .A3(G128), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n244), .A2(KEYINPUT23), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n227), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n573), .A2(G128), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n330), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n572), .B(new_n578), .C1(new_n380), .C2(new_n381), .ZN(new_n579));
  INV_X1    g393(.A(new_n386), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n576), .A2(new_n330), .A3(new_n577), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n571), .B1(new_n568), .B2(new_n570), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n583), .A2(new_n380), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n567), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n572), .B1(new_n380), .B2(new_n381), .ZN(new_n586));
  INV_X1    g400(.A(new_n578), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n583), .A2(new_n380), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(new_n566), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n585), .A2(new_n590), .A3(new_n194), .ZN(new_n591));
  NOR2_X1   g405(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n592), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n585), .A2(new_n590), .A3(new_n194), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n472), .B1(G234), .B2(new_n194), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n561), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n597), .ZN(new_n599));
  AOI211_X1 g413(.A(KEYINPUT78), .B(new_n599), .C1(new_n593), .C2(new_n595), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n585), .A2(new_n590), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n601), .A2(G902), .A3(new_n597), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n598), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n496), .A2(new_n557), .A3(new_n560), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  NAND2_X1  g419(.A1(new_n547), .A2(new_n194), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n606), .A2(G472), .B1(new_n541), .B2(new_n547), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n559), .A2(new_n292), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n607), .A2(new_n608), .A3(new_n603), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n476), .A2(new_n477), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n488), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n486), .A2(KEYINPUT33), .A3(new_n487), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n194), .A2(G478), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n433), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT98), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT34), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(new_n200), .ZN(G6));
  AND2_X1   g436(.A1(new_n491), .A2(new_n482), .ZN(new_n623));
  INV_X1    g437(.A(new_n425), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n384), .A2(new_n390), .A3(new_n406), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n427), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n416), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n628), .A2(KEYINPUT99), .A3(new_n428), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT99), .B1(new_n628), .B2(new_n428), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n623), .A2(new_n415), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n609), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  OAI22_X1  g449(.A1(new_n579), .A2(new_n584), .B1(KEYINPUT36), .B2(new_n567), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT36), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n588), .A2(new_n637), .A3(new_n589), .A4(new_n566), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n636), .A2(new_n194), .A3(new_n599), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT100), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n598), .A2(new_n600), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(G472), .B1(new_n537), .B2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n547), .A2(new_n541), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT101), .A4(new_n644), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n647), .A2(new_n496), .A3(new_n560), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT37), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n330), .ZN(G12));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n190), .B1(new_n196), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n623), .A2(new_n631), .A3(new_n415), .A4(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n641), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n290), .A2(new_n291), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n187), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n557), .A2(new_n656), .A3(new_n559), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XNOR2_X1  g475(.A(new_n653), .B(KEYINPUT39), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n559), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT40), .ZN(new_n665));
  INV_X1    g479(.A(new_n501), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n528), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n501), .A2(new_n509), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n552), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n194), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n543), .A2(new_n548), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n623), .A2(new_n433), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n672), .A2(new_n187), .A3(new_n641), .A4(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n657), .A2(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n657), .A2(KEYINPUT102), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT38), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n676), .A2(KEYINPUT38), .A3(new_n677), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n665), .A2(new_n675), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n248), .ZN(G45));
  NAND3_X1  g497(.A1(new_n616), .A2(new_n433), .A3(new_n654), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n641), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n557), .A2(new_n559), .A3(new_n685), .A4(new_n659), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  AND2_X1   g501(.A1(new_n557), .A2(new_n603), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n353), .A2(new_n345), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n353), .A2(new_n345), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n493), .A3(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n691), .A2(new_n658), .A3(new_n197), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n618), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT103), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n694), .B(new_n696), .ZN(G15));
  NAND2_X1  g511(.A1(new_n693), .A2(new_n632), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  NOR4_X1   g513(.A1(new_n641), .A2(new_n433), .A3(new_n623), .A4(new_n197), .ZN(new_n700));
  INV_X1    g514(.A(new_n691), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(new_n659), .A3(new_n557), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  NAND2_X1  g517(.A1(new_n553), .A2(new_n666), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n704), .B1(new_n545), .B2(new_n546), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n541), .B(KEYINPUT104), .Z(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n643), .A2(new_n603), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n674), .A3(new_n692), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G122), .ZN(G24));
  NOR2_X1   g524(.A1(new_n691), .A2(new_n658), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n685), .A2(new_n643), .A3(new_n711), .A4(new_n707), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  NOR2_X1   g527(.A1(new_n657), .A2(new_n188), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n341), .A2(new_n342), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G469), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n354), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n493), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n684), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n557), .A2(new_n603), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(KEYINPUT105), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n557), .B2(new_n603), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n722), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n723), .A2(new_n721), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n684), .A2(KEYINPUT42), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n727), .A2(KEYINPUT42), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G131), .ZN(G33));
  NOR3_X1   g545(.A1(new_n723), .A2(new_n721), .A3(new_n655), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n306), .ZN(G36));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n335), .B1(new_n334), .B2(new_n339), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT82), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(KEYINPUT106), .A3(G469), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT45), .B1(new_n340), .B2(new_n343), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n739), .B1(new_n740), .B2(new_n345), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n716), .A2(KEYINPUT45), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n738), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n346), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n744), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n690), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n493), .ZN(new_n750));
  INV_X1    g564(.A(new_n607), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n616), .A2(new_n432), .A3(new_n415), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT108), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n616), .A2(KEYINPUT43), .A3(new_n432), .A4(new_n415), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n752), .A2(new_n757), .A3(new_n753), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n751), .A2(new_n759), .A3(new_n642), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n714), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  OR4_X1    g577(.A1(new_n662), .A2(new_n750), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT109), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n299), .ZN(G39));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n749), .B2(new_n493), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n767), .A2(new_n768), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n750), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n771), .B1(new_n773), .B2(new_n770), .ZN(new_n774));
  INV_X1    g588(.A(new_n684), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n557), .A2(new_n603), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n774), .A2(new_n775), .A3(new_n714), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  NOR2_X1   g592(.A1(new_n752), .A2(new_n188), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n493), .A2(new_n681), .A3(new_n603), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n672), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n689), .A2(new_n690), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT49), .Z(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT111), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n782), .A2(new_n493), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n769), .B1(new_n750), .B2(new_n772), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n788), .B2(new_n771), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n759), .A2(new_n708), .A3(new_n190), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n789), .A2(new_n790), .A3(new_n714), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n715), .A2(new_n691), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n603), .A2(new_n190), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n616), .A2(new_n433), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n781), .A2(new_n793), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n759), .A2(new_n190), .A3(new_n642), .A4(new_n793), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n643), .A2(new_n707), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n691), .A2(new_n187), .ZN(new_n803));
  INV_X1    g617(.A(new_n677), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n657), .A2(KEYINPUT102), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT38), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n802), .B(new_n803), .C1(new_n807), .C2(new_n678), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(new_n190), .A3(new_n708), .A4(new_n759), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n802), .B1(new_n681), .B2(new_n803), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n801), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n803), .B1(new_n807), .B2(new_n678), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT117), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n791), .A2(new_n813), .A3(KEYINPUT50), .A4(new_n808), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n792), .A2(new_n800), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n791), .A2(new_n711), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n781), .A2(new_n793), .A3(new_n794), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n189), .B(G953), .C1(new_n820), .C2(new_n618), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n724), .A2(new_n726), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT48), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n759), .A2(new_n190), .A3(new_n793), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n823), .B1(new_n822), .B2(new_n824), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n821), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n789), .A2(new_n714), .A3(new_n791), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n800), .A2(KEYINPUT118), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n799), .B2(new_n817), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n815), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n817), .A2(KEYINPUT116), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n819), .B(new_n828), .C1(new_n829), .C2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n818), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n837), .B1(new_n818), .B2(new_n836), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n694), .A2(new_n698), .A3(new_n702), .A4(new_n709), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n617), .A2(KEYINPUT112), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n616), .A2(new_n843), .A3(new_n433), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n607), .A2(new_n608), .A3(new_n603), .A4(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n604), .A2(KEYINPUT113), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT113), .B1(new_n604), .B2(new_n846), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n479), .A2(new_n481), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n433), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n609), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n649), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n841), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n604), .A2(new_n846), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n604), .A2(new_n846), .A3(KEYINPUT113), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n649), .A2(new_n853), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT114), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n840), .B1(new_n855), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n660), .A2(new_n686), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n719), .A2(new_n673), .A3(new_n658), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n672), .A3(new_n641), .A4(new_n654), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n864), .A2(KEYINPUT52), .A3(new_n712), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n660), .A3(new_n686), .A4(new_n712), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n629), .A2(new_n630), .A3(new_n653), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n415), .A2(new_n714), .A3(new_n851), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n557), .A2(new_n873), .A3(new_n559), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n720), .A2(new_n643), .A3(new_n775), .A4(new_n707), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n642), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n688), .A2(new_n632), .A3(new_n654), .A4(new_n720), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n641), .B1(new_n874), .B2(new_n875), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT115), .B1(new_n881), .B2(new_n732), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n871), .A2(new_n883), .A3(new_n730), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n863), .A2(KEYINPUT53), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT53), .B1(new_n863), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT54), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n888));
  INV_X1    g702(.A(new_n840), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n849), .A2(new_n841), .A3(new_n854), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT114), .B1(new_n860), .B2(new_n861), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n871), .A2(new_n883), .A3(new_n730), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n863), .A2(new_n884), .A3(KEYINPUT53), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n887), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n838), .A2(new_n839), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(G952), .A2(G953), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n785), .B1(new_n899), .B2(new_n900), .ZN(G75));
  AOI21_X1  g715(.A(new_n194), .B1(new_n894), .B2(new_n896), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(G210), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n242), .A2(new_n278), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n276), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  XOR2_X1   g720(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n907));
  AND3_X1   g721(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n906), .B1(new_n903), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n195), .A2(G952), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(G51));
  XNOR2_X1  g726(.A(new_n346), .B(KEYINPUT57), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n898), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n347), .A2(new_n352), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n743), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n902), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n911), .B1(new_n916), .B2(new_n918), .ZN(G54));
  NAND3_X1  g733(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n624), .A3(new_n625), .ZN(new_n921));
  INV_X1    g735(.A(new_n911), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .A4(new_n626), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G60));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n898), .A2(new_n927), .B1(new_n612), .B2(new_n613), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n614), .B(new_n926), .C1(new_n887), .C2(new_n897), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n911), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT60), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n636), .A2(new_n638), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT121), .Z(new_n935));
  OAI211_X1 g749(.A(new_n933), .B(new_n935), .C1(new_n885), .C2(new_n886), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n932), .B1(new_n894), .B2(new_n896), .ZN(new_n937));
  INV_X1    g751(.A(new_n601), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n936), .B(new_n922), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  OAI211_X1 g754(.A(KEYINPUT122), .B(new_n922), .C1(new_n937), .C2(new_n938), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n933), .B1(new_n885), .B2(new_n886), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n911), .B1(new_n943), .B2(new_n601), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n944), .B(new_n936), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n945), .ZN(G66));
  NOR2_X1   g760(.A1(new_n863), .A2(G953), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT123), .ZN(new_n948));
  INV_X1    g762(.A(G224), .ZN(new_n949));
  OAI21_X1  g763(.A(G953), .B1(new_n193), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n904), .B1(G898), .B2(new_n195), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G69));
  OAI21_X1  g767(.A(new_n422), .B1(new_n378), .B2(new_n421), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n527), .B(new_n954), .Z(new_n955));
  NAND2_X1  g769(.A1(G900), .A2(G953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n724), .A2(new_n726), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n673), .A2(new_n658), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NOR4_X1   g773(.A1(new_n750), .A2(new_n957), .A3(new_n662), .A4(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n660), .A2(new_n686), .A3(new_n712), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n732), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n730), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n960), .B2(KEYINPUT126), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(new_n764), .A3(new_n777), .A4(new_n965), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n955), .B(new_n956), .C1(new_n966), .C2(G953), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT124), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT62), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n682), .A2(new_n962), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n968), .A2(new_n969), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n845), .A2(new_n852), .ZN(new_n974));
  OR4_X1    g788(.A1(new_n723), .A2(new_n974), .A3(new_n664), .A4(new_n715), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n777), .A2(new_n973), .A3(new_n764), .A4(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n955), .B1(new_n976), .B2(new_n195), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n967), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n981), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n967), .A2(new_n979), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n976), .B2(new_n892), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n667), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n528), .A2(new_n501), .ZN(new_n990));
  OAI221_X1 g804(.A(new_n987), .B1(new_n990), .B2(new_n550), .C1(new_n885), .C2(new_n886), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n989), .A2(new_n991), .A3(new_n922), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n993), .B(new_n987), .C1(new_n966), .C2(new_n892), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n994), .A2(new_n668), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n987), .B1(new_n966), .B2(new_n892), .ZN(new_n996));
  AOI22_X1  g810(.A1(new_n996), .A2(KEYINPUT127), .B1(new_n238), .B2(new_n527), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n992), .B1(new_n995), .B2(new_n997), .ZN(G57));
endmodule


