//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n450, new_n453, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n550, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n591, new_n594, new_n596, new_n597, new_n598,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g029(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT69), .Z(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(G137), .A3(new_n464), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n464), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G112), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT70), .Z(new_n481));
  AOI21_X1  g056(.A(new_n464), .B1(new_n477), .B2(new_n478), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n476), .B(new_n481), .C1(G124), .C2(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  OAI211_X1 g060(.A(G138), .B(new_n464), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n465), .A2(new_n488), .A3(G138), .A4(new_n464), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n464), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n482), .A2(G126), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(G62), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(G75), .A2(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(G651), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT71), .B1(new_n503), .B2(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(G651), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n508), .A2(G50), .A3(G543), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n498), .A2(new_n499), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n502), .B(new_n510), .C1(new_n512), .C2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  INV_X1    g092(.A(G89), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n508), .A2(G543), .A3(new_n509), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n511), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n506), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n524), .A2(G51), .B1(new_n526), .B2(G63), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n521), .A2(new_n522), .A3(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  INV_X1    g104(.A(new_n512), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n524), .A2(G52), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n506), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  NAND2_X1  g111(.A1(G68), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G56), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n525), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(new_n540), .A3(G651), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n508), .A2(G81), .A3(new_n509), .A4(new_n511), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n508), .A2(G43), .A3(G543), .A4(new_n509), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT73), .B1(new_n545), .B2(new_n506), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n541), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT74), .ZN(G176));
  XOR2_X1   g126(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n552));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND4_X1  g130(.A1(new_n508), .A2(G53), .A3(G543), .A4(new_n509), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n525), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n530), .A2(G91), .B1(new_n560), .B2(G651), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G299));
  OAI21_X1  g137(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT76), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n524), .A2(G49), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n530), .A2(G87), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  INV_X1    g142(.A(G61), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n498), .B2(new_n499), .ZN(new_n569));
  AND2_X1   g144(.A1(G73), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n508), .A2(G48), .A3(G543), .A4(new_n509), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n508), .A2(G86), .A3(new_n509), .A4(new_n511), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G305));
  NAND2_X1  g149(.A1(new_n530), .A2(G85), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n524), .A2(G47), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n506), .C2(new_n577), .ZN(G290));
  NAND2_X1  g153(.A1(G301), .A2(G868), .ZN(new_n579));
  INV_X1    g154(.A(G54), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n580), .A2(new_n523), .B1(new_n581), .B2(new_n506), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n530), .A2(KEYINPUT10), .A3(G92), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT10), .ZN(new_n584));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n512), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n582), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n579), .B1(G868), .B2(new_n587), .ZN(G284));
  OAI21_X1  g163(.A(new_n579), .B1(G868), .B2(new_n587), .ZN(G321));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NAND2_X1  g165(.A1(G299), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n591), .B1(G168), .B2(new_n590), .ZN(G297));
  OAI21_X1  g167(.A(new_n591), .B1(G168), .B2(new_n590), .ZN(G280));
  INV_X1    g168(.A(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n587), .B1(new_n594), .B2(G860), .ZN(G148));
  NOR2_X1   g170(.A1(new_n548), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n587), .A2(new_n594), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT77), .ZN(G323));
  XNOR2_X1  g174(.A(KEYINPUT78), .B(KEYINPUT11), .ZN(new_n600));
  XNOR2_X1  g175(.A(G323), .B(new_n600), .ZN(G282));
  NAND2_X1  g176(.A1(new_n465), .A2(new_n470), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT13), .ZN(new_n604));
  INV_X1    g179(.A(G2100), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n479), .A2(G135), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n482), .A2(G123), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n464), .A2(G111), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(G2096), .Z(new_n613));
  NAND3_X1  g188(.A1(new_n606), .A2(new_n607), .A3(new_n613), .ZN(G156));
  XNOR2_X1  g189(.A(G2427), .B(G2438), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2430), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT15), .B(G2435), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n618), .A2(KEYINPUT14), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2451), .B(G2454), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT16), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n620), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G2443), .B(G2446), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G1341), .B(G1348), .Z(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT79), .Z(new_n628));
  OAI21_X1  g203(.A(G14), .B1(new_n625), .B2(new_n626), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n628), .A2(new_n629), .ZN(G401));
  XNOR2_X1  g205(.A(G2067), .B(G2678), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT80), .ZN(new_n632));
  XOR2_X1   g207(.A(G2084), .B(G2090), .Z(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2072), .B(G2078), .Z(new_n635));
  NOR3_X1   g210(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT18), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(KEYINPUT17), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n638), .A2(new_n633), .A3(new_n632), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n633), .B1(new_n632), .B2(new_n635), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n640), .A2(KEYINPUT81), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(KEYINPUT81), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n632), .B2(new_n638), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n637), .B(new_n639), .C1(new_n641), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2096), .B(G2100), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(G227));
  XOR2_X1   g221(.A(G1971), .B(G1976), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT19), .ZN(new_n648));
  XOR2_X1   g223(.A(G1956), .B(G2474), .Z(new_n649));
  XOR2_X1   g224(.A(G1961), .B(G1966), .Z(new_n650));
  AND2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n649), .A2(new_n650), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  MUX2_X1   g231(.A(new_n656), .B(new_n655), .S(new_n648), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1991), .B(G1996), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1981), .B(G1986), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G229));
  INV_X1    g239(.A(G29), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G35), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(G162), .B2(new_n665), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT29), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n668), .A2(G2090), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(G2090), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT83), .B(G16), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G20), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT23), .Z(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(G299), .B2(G16), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT95), .B(G1956), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n669), .A2(new_n670), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n665), .A2(G33), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n465), .A2(G127), .ZN(new_n679));
  NAND2_X1  g254(.A1(G115), .A2(G2104), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n464), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT25), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI211_X1 g261(.A(new_n681), .B(new_n686), .C1(G139), .C2(new_n479), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT92), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n678), .B1(new_n688), .B2(new_n665), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G2072), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G4), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n587), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1348), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(G5), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G171), .B2(new_n691), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1961), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n690), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n691), .A2(G21), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G168), .B2(new_n691), .ZN(new_n700));
  INV_X1    g275(.A(G1966), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n470), .A2(G105), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT26), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n479), .A2(G141), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n482), .A2(G129), .ZN(new_n707));
  AND4_X1   g282(.A1(new_n703), .A2(new_n705), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G29), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G29), .B2(G32), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT27), .B(G1996), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT93), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n612), .A2(new_n665), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT31), .B(G11), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT94), .ZN(new_n716));
  INV_X1    g291(.A(G28), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT30), .ZN(new_n718));
  AOI21_X1  g293(.A(G29), .B1(new_n717), .B2(KEYINPUT30), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND3_X1   g295(.A1(new_n713), .A2(new_n714), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n674), .A2(new_n675), .ZN(new_n722));
  NOR2_X1   g297(.A1(G164), .A2(new_n665), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G27), .B2(new_n665), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(new_n443), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n443), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n721), .A2(new_n722), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n671), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n728), .A2(G19), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n548), .B2(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G1341), .ZN(new_n731));
  INV_X1    g306(.A(G34), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n732), .A2(KEYINPUT24), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(KEYINPUT24), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n665), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G160), .B2(new_n665), .ZN(new_n736));
  INV_X1    g311(.A(G2084), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n710), .A2(new_n712), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n731), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n665), .A2(G26), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT28), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n479), .A2(G140), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT91), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n746));
  INV_X1    g321(.A(G116), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(G2105), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G128), .B2(new_n482), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n742), .B1(new_n750), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2067), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G1341), .B2(new_n730), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n727), .A2(new_n740), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n677), .A2(new_n698), .A3(new_n702), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT90), .B(KEYINPUT36), .ZN(new_n756));
  MUX2_X1   g331(.A(G6), .B(G305), .S(G16), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT85), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT32), .B(G1981), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n691), .A2(G23), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G288), .B2(G16), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT87), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT33), .B(G1976), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT86), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n760), .B(new_n761), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n764), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n671), .A2(G22), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT88), .Z(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G166), .B2(new_n671), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1971), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT84), .B(KEYINPUT34), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n767), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n665), .A2(G25), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n479), .A2(G131), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n482), .A2(G119), .ZN(new_n779));
  OR2_X1    g354(.A1(G95), .A2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n780), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n777), .B1(new_n783), .B2(new_n665), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT82), .Z(new_n785));
  XOR2_X1   g360(.A(KEYINPUT35), .B(G1991), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G24), .B(G290), .S(new_n728), .Z(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1986), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n776), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT89), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n775), .B1(new_n767), .B2(new_n773), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n756), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n792), .A2(new_n793), .A3(new_n756), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n755), .B1(new_n795), .B2(new_n796), .ZN(G311));
  INV_X1    g372(.A(new_n755), .ZN(new_n798));
  INV_X1    g373(.A(new_n796), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n794), .ZN(G150));
  INV_X1    g375(.A(G55), .ZN(new_n801));
  INV_X1    g376(.A(G93), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n801), .A2(new_n523), .B1(new_n512), .B2(new_n802), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n804), .A2(KEYINPUT97), .A3(new_n506), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT97), .B1(new_n804), .B2(new_n506), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n541), .A2(new_n544), .A3(KEYINPUT98), .A4(new_n546), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT99), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n547), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n812), .B1(new_n547), .B2(new_n811), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n810), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n547), .A2(new_n811), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT99), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n818), .A2(new_n809), .A3(new_n808), .A4(new_n813), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n587), .A2(G559), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n820), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n825));
  AOI21_X1  g400(.A(G860), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n825), .B2(new_n824), .ZN(new_n827));
  INV_X1    g402(.A(new_n808), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G860), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(new_n831), .ZN(G145));
  XNOR2_X1  g407(.A(new_n750), .B(KEYINPUT102), .ZN(new_n833));
  INV_X1    g408(.A(new_n708), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT102), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n750), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n708), .ZN(new_n838));
  INV_X1    g413(.A(new_n494), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT101), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n488), .B1(new_n479), .B2(G138), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT101), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n839), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n835), .A2(new_n838), .A3(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n845), .B1(new_n835), .B2(new_n838), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n687), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n835), .A2(new_n838), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT101), .ZN(new_n851));
  AOI21_X1  g426(.A(KEYINPUT101), .B1(new_n487), .B2(new_n489), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n494), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n688), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(new_n855), .A3(new_n846), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n482), .A2(G130), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n464), .A2(G118), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(G142), .B2(new_n479), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n603), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n783), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n849), .A2(new_n856), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n864), .B1(new_n849), .B2(new_n856), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(G160), .B(new_n612), .Z(new_n869));
  XOR2_X1   g444(.A(G162), .B(new_n869), .Z(new_n870));
  AOI21_X1  g445(.A(G37), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n872));
  INV_X1    g447(.A(new_n867), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n865), .ZN(new_n874));
  INV_X1    g449(.A(new_n870), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI211_X1 g451(.A(KEYINPUT103), .B(new_n870), .C1(new_n873), .C2(new_n865), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n871), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g454(.A(KEYINPUT106), .B1(new_n808), .B2(G868), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n820), .B(new_n597), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n557), .A2(new_n561), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n583), .A2(new_n586), .ZN(new_n883));
  INV_X1    g458(.A(new_n582), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT104), .B1(G299), .B2(new_n587), .ZN(new_n888));
  NAND2_X1  g463(.A1(G299), .A2(new_n587), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT41), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n881), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n890), .B2(new_n881), .ZN(new_n896));
  XOR2_X1   g471(.A(G288), .B(G305), .Z(new_n897));
  XNOR2_X1  g472(.A(G290), .B(G166), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n897), .B(new_n898), .Z(new_n899));
  XOR2_X1   g474(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n590), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n901), .B2(new_n896), .ZN(new_n903));
  MUX2_X1   g478(.A(KEYINPUT106), .B(new_n880), .S(new_n903), .Z(G295));
  MUX2_X1   g479(.A(KEYINPUT106), .B(new_n880), .S(new_n903), .Z(G331));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n906));
  NAND2_X1  g481(.A1(G286), .A2(G301), .ZN(new_n907));
  NAND4_X1  g482(.A1(G171), .A2(new_n522), .A3(new_n521), .A4(new_n527), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n814), .A2(new_n810), .A3(new_n815), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n818), .A2(new_n813), .B1(new_n809), .B2(new_n808), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n816), .A2(new_n819), .A3(new_n909), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n894), .A2(new_n892), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n820), .A2(KEYINPUT107), .A3(new_n910), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n899), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n913), .A2(new_n890), .A3(new_n915), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n916), .A2(new_n918), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n890), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n892), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n890), .A2(KEYINPUT109), .A3(new_n891), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n894), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n913), .A2(new_n915), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n920), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT43), .B1(new_n924), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n924), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n934), .A2(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n924), .C2(new_n933), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n906), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n924), .B2(new_n936), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n930), .A2(new_n931), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n893), .B1(new_n916), .B2(new_n918), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n899), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(new_n938), .A3(new_n923), .A4(new_n922), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n942), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n919), .A2(new_n921), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n899), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n923), .A3(new_n922), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT108), .B1(new_n951), .B2(KEYINPUT43), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n948), .A2(KEYINPUT44), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n941), .A2(new_n953), .ZN(G397));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n845), .B2(G1384), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n466), .A2(new_n467), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(G2105), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n469), .A2(new_n471), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(G40), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(G290), .A2(G1986), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT48), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n961), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n965));
  INV_X1    g540(.A(new_n962), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n750), .A2(G2067), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n750), .A2(G2067), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n708), .B(G1996), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n783), .A2(new_n786), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n783), .A2(new_n786), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n963), .B(new_n967), .C1(new_n961), .C2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n970), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n961), .B1(new_n976), .B2(new_n834), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n964), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n979));
  INV_X1    g554(.A(G1996), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n961), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT47), .Z(new_n983));
  NAND2_X1  g558(.A1(new_n970), .A2(new_n971), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n968), .B1(new_n984), .B2(new_n973), .ZN(new_n985));
  AOI211_X1 g560(.A(new_n975), .B(new_n983), .C1(new_n961), .C2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n495), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n960), .B1(new_n988), .B2(new_n955), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n955), .A2(G1384), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n853), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(new_n442), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT50), .B1(new_n845), .B2(G1384), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n490), .B2(new_n494), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n960), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(G1956), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT119), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(G299), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  OR2_X1    g578(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1004));
  NAND2_X1  g579(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1005));
  AND4_X1   g580(.A1(new_n557), .A2(new_n561), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT120), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1006), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n1002), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT120), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1001), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n995), .A2(new_n1000), .A3(KEYINPUT119), .ZN(new_n1014));
  INV_X1    g589(.A(G40), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n468), .A2(new_n472), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n853), .A2(new_n987), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G2067), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT50), .B1(new_n853), .B2(new_n987), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n988), .A2(new_n997), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1016), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1348), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1018), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1013), .A2(new_n1014), .B1(new_n885), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n996), .A2(new_n999), .ZN(new_n1025));
  INV_X1    g600(.A(G1956), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1007), .A2(new_n1027), .A3(new_n994), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g604(.A(KEYINPUT58), .B(G1341), .Z(new_n1030));
  NAND2_X1  g605(.A1(new_n1017), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n989), .A2(new_n991), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1031), .B1(new_n1032), .B2(G1996), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT122), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n548), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n990), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n843), .A2(new_n844), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(new_n494), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1016), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1039), .A2(new_n1040), .A3(G1996), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1030), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1384), .B1(new_n1038), .B2(new_n494), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1042), .B1(new_n1043), .B2(new_n1016), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n548), .B(new_n1035), .C1(new_n1041), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT122), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1033), .B2(new_n548), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1036), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT123), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(KEYINPUT123), .B(new_n1036), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1020), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n997), .B1(new_n845), .B2(G1384), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n960), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g631(.A1(new_n1056), .A2(G1348), .B1(G2067), .B2(new_n1017), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT60), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1023), .A2(KEYINPUT60), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n587), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1023), .A2(KEYINPUT60), .A3(new_n885), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT61), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1010), .B1(new_n995), .B2(new_n1000), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1028), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1028), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1061), .B(new_n1062), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1029), .B1(new_n1053), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT45), .B1(new_n853), .B2(new_n987), .ZN(new_n1070));
  NOR2_X1   g645(.A1(G164), .A2(new_n1037), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1070), .A2(new_n960), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(G2078), .ZN(new_n1074));
  INV_X1    g649(.A(G1961), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1072), .A2(new_n1074), .B1(new_n1021), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n989), .A2(new_n991), .A3(new_n443), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1073), .ZN(new_n1078));
  AOI21_X1  g653(.A(G301), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1021), .A2(new_n1075), .ZN(new_n1080));
  AOI21_X1  g655(.A(G171), .B1(new_n1077), .B2(new_n1073), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1074), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n853), .B2(new_n990), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n956), .A2(new_n1083), .A3(new_n1016), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT126), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n956), .A2(new_n1083), .A3(KEYINPUT126), .A4(new_n1016), .ZN(new_n1087));
  AND4_X1   g662(.A1(new_n1080), .A2(new_n1081), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1069), .B1(new_n1079), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G303), .A2(G8), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(G303), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G2090), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1016), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT112), .B(G1971), .Z(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n989), .B2(new_n991), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1097), .B(G8), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G8), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1043), .B2(new_n1016), .ZN(new_n1105));
  INV_X1    g680(.A(G1976), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT52), .B1(G288), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1105), .B(new_n1107), .C1(new_n1106), .C2(G288), .ZN(new_n1108));
  NAND2_X1  g683(.A1(G305), .A2(G1981), .ZN(new_n1109));
  INV_X1    g684(.A(G1981), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT49), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT114), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1109), .A2(new_n1115), .A3(KEYINPUT49), .A4(new_n1111), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(new_n1105), .A3(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1017), .B(G8), .C1(new_n1106), .C2(G288), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT52), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1103), .A2(new_n1108), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1101), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1032), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n996), .A2(new_n1098), .A3(new_n999), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1097), .B1(new_n1126), .B2(G8), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1080), .A2(new_n1086), .A3(new_n1087), .A4(new_n1078), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G171), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1069), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1089), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1071), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n956), .A2(new_n1016), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n701), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n737), .B(new_n1016), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1138), .A2(G8), .A3(G286), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT124), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1138), .A2(new_n1141), .A3(G8), .A4(G286), .ZN(new_n1142));
  NAND2_X1  g717(.A1(G286), .A2(G8), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT51), .B1(new_n1143), .B2(KEYINPUT125), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1056), .A2(new_n737), .B1(new_n1135), .B2(new_n701), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1143), .B(new_n1144), .C1(new_n1145), .C2(new_n1104), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1144), .ZN(new_n1147));
  OAI211_X1 g722(.A(G8), .B(new_n1147), .C1(new_n1138), .C2(G286), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1140), .A2(new_n1142), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1133), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1068), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT62), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1149), .A2(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1128), .A2(new_n1079), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1108), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1127), .ZN(new_n1162));
  AOI211_X1 g737(.A(new_n1104), .B(G286), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1103), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1098), .B(new_n1016), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1104), .B1(new_n1166), .B2(new_n1124), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT63), .B1(new_n1167), .B2(new_n1097), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1122), .A2(new_n1168), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1164), .A2(new_n1165), .B1(new_n1169), .B2(new_n1163), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1111), .B(KEYINPUT115), .Z(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(G288), .A2(G1976), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1172), .B1(new_n1119), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1105), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1160), .A2(new_n1103), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT116), .B1(new_n1170), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT116), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n1128), .B2(new_n1163), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1163), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1183), .A2(new_n1122), .A3(new_n1168), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1178), .B(new_n1181), .C1(new_n1182), .C2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1151), .A2(new_n1159), .A3(new_n1180), .A4(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n962), .A2(KEYINPUT111), .ZN(new_n1188));
  NAND2_X1  g763(.A1(G290), .A2(G1986), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1188), .B(new_n1189), .Z(new_n1190));
  OAI21_X1  g765(.A(new_n961), .B1(new_n1190), .B2(new_n974), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1186), .A2(new_n1187), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1187), .B1(new_n1186), .B2(new_n1191), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n986), .B1(new_n1192), .B2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g769(.A1(G401), .A2(G229), .A3(new_n462), .A4(G227), .ZN(new_n1196));
  OAI211_X1 g770(.A(new_n878), .B(new_n1196), .C1(new_n948), .C2(new_n952), .ZN(G225));
  INV_X1    g771(.A(G225), .ZN(G308));
endmodule


