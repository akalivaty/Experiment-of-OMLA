//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT81), .ZN(new_n203));
  INV_X1    g002(.A(G204gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G197gat), .ZN(new_n205));
  INV_X1    g004(.A(G197gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G204gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT22), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT72), .ZN(new_n209));
  AND2_X1   g008(.A1(G211gat), .A2(G218gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(G211gat), .A2(G218gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G211gat), .A2(G218gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT22), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n214), .A2(new_n205), .A3(new_n217), .A4(new_n207), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n209), .B1(new_n208), .B2(new_n212), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G155gat), .B(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(G155gat), .ZN(new_n226));
  INV_X1    g025(.A(G162gat), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT2), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(G141gat), .A2(G148gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n231));
  NAND2_X1  g030(.A1(G141gat), .A2(G148gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n229), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G228gat), .A2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n229), .A2(new_n237), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n240), .B1(new_n219), .B2(new_n220), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n243), .B(KEYINPUT80), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n229), .A2(new_n237), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n208), .A2(new_n212), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT29), .B1(new_n218), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n238), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n251), .B1(new_n242), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(G22gat), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n256), .ZN(new_n259));
  INV_X1    g058(.A(new_n251), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n243), .B1(new_n221), .B2(new_n241), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n253), .A2(KEYINPUT72), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(new_n213), .A3(new_n218), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT3), .B1(new_n264), .B2(new_n240), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n262), .B1(new_n265), .B2(new_n246), .ZN(new_n266));
  INV_X1    g065(.A(G22gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n261), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n203), .B1(new_n258), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G78gat), .B(G106gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT31), .B(G50gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT82), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n261), .A2(new_n266), .A3(new_n267), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n267), .B1(new_n261), .B2(new_n266), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT81), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT82), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n272), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT81), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n274), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n280), .B1(new_n274), .B2(new_n279), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(KEYINPUT27), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n292), .B1(KEYINPUT66), .B2(G183gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n288), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT68), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n289), .A2(KEYINPUT28), .ZN(new_n296));
  INV_X1    g095(.A(G183gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT27), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n292), .A2(G183gat), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT69), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT69), .B1(new_n298), .B2(new_n299), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n296), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n288), .B(new_n303), .C1(new_n291), .C2(new_n293), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n295), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT26), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n307), .A2(new_n311), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT64), .B1(new_n306), .B2(KEYINPUT23), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT64), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n315), .B(new_n316), .C1(G169gat), .C2(G176gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  OR2_X1    g117(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(G190gat), .A3(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n289), .A2(new_n322), .B1(new_n306), .B2(KEYINPUT23), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n318), .A2(new_n321), .A3(new_n311), .A4(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G169gat), .ZN(new_n327));
  INV_X1    g126(.A(G176gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT23), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n289), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n310), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n329), .B(new_n330), .C1(new_n331), .C2(new_n308), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n333), .A2(KEYINPUT25), .A3(new_n318), .A4(new_n321), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n285), .B1(new_n336), .B2(new_n240), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n305), .A2(new_n312), .B1(new_n326), .B2(new_n334), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(new_n284), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n221), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n284), .B1(new_n338), .B2(KEYINPUT29), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(new_n285), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n264), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT73), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(new_n344), .A3(new_n264), .ZN(new_n347));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n342), .A2(new_n346), .A3(new_n347), .A4(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n342), .A2(new_n346), .A3(new_n347), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n350), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n354), .B1(new_n352), .B2(new_n353), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT1), .ZN(new_n361));
  AND2_X1   g160(.A1(G113gat), .A2(G120gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(G113gat), .A2(G120gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G134gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G127gat), .ZN(new_n366));
  INV_X1    g165(.A(G127gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G134gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT70), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n361), .B(new_n364), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G113gat), .ZN(new_n372));
  INV_X1    g171(.A(G120gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G113gat), .A2(G120gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n361), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n370), .A3(new_n375), .ZN(new_n377));
  XNOR2_X1  g176(.A(G127gat), .B(G134gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n380), .B(new_n239), .C1(new_n248), .C2(new_n246), .ZN(new_n381));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(KEYINPUT5), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n252), .B1(new_n371), .B2(new_n379), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT78), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n379), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT76), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n246), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n246), .B2(new_n388), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n387), .B1(new_n392), .B2(KEYINPUT4), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT76), .B1(new_n380), .B2(new_n252), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n246), .A2(new_n388), .A3(new_n389), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT4), .A4(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n381), .B(new_n384), .C1(new_n393), .C2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n246), .A2(new_n388), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n390), .A2(new_n391), .A3(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n400), .B(KEYINPUT5), .C1(new_n402), .C2(new_n382), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n394), .A2(new_n386), .A3(new_n396), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n246), .A2(new_n388), .A3(KEYINPUT4), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n404), .A2(new_n382), .A3(new_n405), .A4(new_n381), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n380), .A2(new_n252), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n394), .A2(new_n408), .A3(new_n396), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n383), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n400), .B1(new_n410), .B2(KEYINPUT5), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n399), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  XOR2_X1   g216(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n412), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n416), .B(new_n399), .C1(new_n407), .C2(new_n411), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n418), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT5), .B1(new_n402), .B2(new_n382), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT77), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(new_n403), .A3(new_n406), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n416), .B1(new_n425), .B2(new_n399), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n420), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n283), .B1(new_n360), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n313), .A2(new_n388), .A3(new_n335), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n388), .B1(new_n313), .B2(new_n335), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(KEYINPUT32), .ZN(new_n436));
  XOR2_X1   g235(.A(G15gat), .B(G43gat), .Z(new_n437));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n439), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n433), .B(KEYINPUT32), .C1(new_n434), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n431), .A2(new_n432), .A3(new_n430), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT34), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT71), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n336), .A2(new_n380), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n338), .A2(new_n388), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n429), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT71), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT34), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(new_n445), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n446), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n443), .A2(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n451), .A2(new_n452), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n455), .A2(new_n446), .A3(new_n442), .A4(new_n440), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT36), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(new_n456), .A3(KEYINPUT36), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n202), .B1(new_n428), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n274), .A2(new_n279), .ZN(new_n463));
  INV_X1    g262(.A(new_n280), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n274), .A2(new_n279), .A3(new_n280), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT40), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n396), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n246), .A2(new_n388), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n395), .B1(new_n470), .B2(KEYINPUT4), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n397), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n382), .B1(new_n473), .B2(new_n381), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n402), .A2(new_n382), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT39), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n416), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n381), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n472), .B2(new_n397), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n479), .A2(KEYINPUT39), .A3(new_n382), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n468), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n480), .ZN(new_n482));
  OAI211_X1 g281(.A(KEYINPUT39), .B(new_n475), .C1(new_n479), .C2(new_n382), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT40), .A4(new_n416), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n412), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT84), .B(new_n399), .C1(new_n407), .C2(new_n411), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n416), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n352), .A2(new_n353), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT30), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(new_n355), .A3(new_n357), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n467), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT86), .B(KEYINPUT37), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n342), .A2(new_n346), .A3(new_n347), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT87), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n337), .A2(new_n339), .A3(new_n221), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n341), .B2(new_n340), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n346), .A4(new_n495), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(KEYINPUT85), .B(KEYINPUT37), .C1(new_n498), .C2(new_n345), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT37), .B1(new_n498), .B2(new_n345), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n351), .A2(KEYINPUT38), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n502), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n488), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT84), .B1(new_n425), .B2(new_n399), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n417), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n422), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n509), .A2(new_n514), .A3(new_n420), .A4(new_n352), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT38), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n351), .B1(new_n356), .B2(KEYINPUT37), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n516), .B1(new_n502), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n494), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n427), .A2(new_n492), .A3(new_n355), .A4(new_n357), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n520), .A2(new_n467), .B1(new_n459), .B2(new_n460), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT83), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n462), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n467), .A2(new_n457), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n514), .A2(new_n420), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT35), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n360), .ZN(new_n527));
  INV_X1    g326(.A(new_n457), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n283), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT35), .B1(new_n529), .B2(new_n520), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n523), .A2(KEYINPUT88), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT88), .B1(new_n523), .B2(new_n531), .ZN(new_n533));
  NOR2_X1   g332(.A1(G29gat), .A2(G36gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT14), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT91), .B(G36gat), .Z(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT90), .B(G29gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n536), .A2(KEYINPUT89), .A3(new_n537), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(G43gat), .B(G50gat), .Z(new_n546));
  INV_X1    g345(.A(KEYINPUT15), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n546), .A2(new_n547), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n547), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n550), .A2(new_n538), .A3(new_n543), .A4(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT92), .B1(new_n553), .B2(KEYINPUT17), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n552), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT92), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n553), .A2(KEYINPUT93), .A3(KEYINPUT17), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n555), .B2(new_n557), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G15gat), .B(G22gat), .ZN(new_n564));
  INV_X1    g363(.A(G1gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(KEYINPUT16), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n565), .B2(new_n564), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G8gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n559), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n553), .A2(new_n568), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n569), .A2(KEYINPUT18), .A3(new_n570), .A4(new_n571), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n553), .B(new_n568), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n570), .B(KEYINPUT13), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G113gat), .B(G141gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT11), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(new_n327), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G197gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT12), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n574), .A2(new_n575), .A3(new_n578), .A4(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT95), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT94), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n587));
  INV_X1    g386(.A(new_n583), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n586), .A3(new_n588), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n585), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n532), .A2(new_n533), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  INV_X1    g397(.A(G85gat), .ZN(new_n599));
  INV_X1    g398(.A(G92gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G99gat), .B(G106gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT102), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n602), .B(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n605), .A2(new_n555), .B1(KEYINPUT41), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n559), .A2(new_n563), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n607), .B1(new_n608), .B2(new_n605), .ZN(new_n609));
  XOR2_X1   g408(.A(G190gat), .B(G218gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n606), .A2(KEYINPUT41), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n611), .A2(new_n613), .ZN(new_n615));
  XOR2_X1   g414(.A(G134gat), .B(G162gat), .Z(new_n616));
  OR3_X1    g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n616), .B1(new_n614), .B2(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G183gat), .B(G211gat), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G71gat), .B(G78gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT96), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G57gat), .B(G64gat), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n625), .A2(KEYINPUT97), .ZN(new_n627));
  INV_X1    g426(.A(new_n624), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(KEYINPUT97), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n622), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT98), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT99), .B(KEYINPUT19), .Z(new_n637));
  AND2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G127gat), .B(G155gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT20), .Z(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n636), .B(new_n637), .ZN(new_n644));
  INV_X1    g443(.A(new_n642), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n621), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n640), .A2(new_n642), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n645), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n649), .A3(new_n620), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n568), .B1(new_n631), .B2(new_n632), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT100), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n647), .A2(new_n653), .A3(new_n650), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT103), .B1(new_n619), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(new_n617), .A3(new_n660), .A4(new_n618), .ZN(new_n661));
  INV_X1    g460(.A(G230gat), .ZN(new_n662));
  INV_X1    g461(.A(G233gat), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n626), .A2(new_n630), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n605), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n602), .A2(new_n604), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n602), .A2(new_n604), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n631), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n667), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n667), .A2(KEYINPUT104), .A3(new_n671), .A4(new_n668), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n667), .A2(new_n668), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n665), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n667), .A2(new_n671), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n665), .ZN(new_n680));
  XNOR2_X1  g479(.A(G120gat), .B(G148gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n658), .A2(new_n661), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n594), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n427), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(new_n565), .ZN(G1324gat));
  NOR2_X1   g490(.A1(new_n689), .A2(new_n360), .ZN(new_n692));
  INV_X1    g491(.A(G8gat), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  AOI21_X1  g494(.A(KEYINPUT105), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n697), .B2(new_n696), .ZN(G1325gat));
  NAND3_X1  g498(.A1(new_n594), .A2(new_n461), .A3(new_n688), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G15gat), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n457), .A2(G15gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n689), .B2(new_n702), .ZN(G1326gat));
  NOR2_X1   g502(.A1(new_n689), .A2(new_n283), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT43), .B(G22gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  INV_X1    g505(.A(new_n427), .ZN(new_n707));
  INV_X1    g506(.A(new_n542), .ZN(new_n708));
  INV_X1    g507(.A(new_n619), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n659), .A3(new_n686), .ZN(new_n710));
  AND4_X1   g509(.A1(new_n707), .A2(new_n594), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT45), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n420), .B(new_n352), .C1(new_n489), .C2(new_n422), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n506), .A2(new_n503), .A3(new_n507), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n497), .B2(new_n501), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n713), .A2(new_n518), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n512), .A2(new_n484), .A3(new_n481), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n283), .B1(new_n717), .B2(new_n360), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n521), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n719), .A2(new_n531), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n719), .B2(new_n531), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n619), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  OAI22_X1  g524(.A1(new_n716), .A2(new_n718), .B1(new_n521), .B2(KEYINPUT83), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n428), .A2(new_n461), .A3(new_n202), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n531), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT88), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n523), .A2(KEYINPUT88), .A3(new_n531), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n731), .A3(new_n619), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n725), .B1(new_n732), .B2(KEYINPUT44), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n592), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n585), .B(KEYINPUT106), .C1(new_n589), .C2(new_n591), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n686), .B(KEYINPUT107), .Z(new_n738));
  NOR4_X1   g537(.A1(new_n733), .A2(new_n659), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n708), .B1(new_n739), .B2(new_n707), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n712), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT109), .ZN(G1328gat));
  NAND2_X1  g541(.A1(new_n594), .A2(new_n710), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n360), .A2(new_n541), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT46), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT110), .Z(new_n748));
  NAND2_X1  g547(.A1(new_n739), .A2(new_n493), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n541), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n748), .B(new_n750), .C1(KEYINPUT46), .C2(new_n746), .ZN(G1329gat));
  AOI21_X1  g550(.A(G43gat), .B1(new_n744), .B2(new_n528), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n461), .A2(G43gat), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n739), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756));
  INV_X1    g555(.A(G50gat), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n739), .B2(new_n467), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n743), .A2(G50gat), .A3(new_n283), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n739), .A2(new_n467), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n759), .A2(new_n756), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(G1331gat));
  AND2_X1   g565(.A1(new_n658), .A2(new_n661), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n767), .A2(new_n737), .A3(new_n738), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n768), .A2(new_n722), .A3(new_n721), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n707), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g570(.A1(new_n493), .A2(KEYINPUT112), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n493), .A2(KEYINPUT112), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  AND2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n776), .B2(new_n775), .ZN(G1333gat));
  INV_X1    g578(.A(G71gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n457), .B(KEYINPUT113), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n769), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n769), .A2(new_n461), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n780), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n467), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g586(.A1(new_n737), .A2(new_n657), .A3(new_n619), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n531), .B2(new_n719), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT51), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT115), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n792), .A3(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n789), .A2(KEYINPUT51), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(new_n599), .A3(new_n707), .A4(new_n686), .ZN(new_n797));
  INV_X1    g596(.A(new_n725), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n532), .A2(new_n533), .A3(new_n709), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n723), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n737), .A2(new_n657), .A3(new_n686), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(KEYINPUT114), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n733), .B2(new_n801), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(new_n707), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n797), .B1(new_n807), .B2(new_n599), .ZN(G1336gat));
  NAND3_X1  g607(.A1(new_n738), .A2(new_n600), .A3(new_n774), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n794), .B2(new_n795), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n800), .A2(new_n774), .A3(new_n802), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n811), .B(new_n812), .C1(new_n600), .C2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n803), .A2(new_n805), .A3(new_n493), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G92gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n811), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT116), .B1(new_n817), .B2(KEYINPUT52), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n810), .B1(new_n815), .B2(G92gat), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n819), .A2(new_n820), .A3(new_n812), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n814), .B1(new_n818), .B2(new_n821), .ZN(G1337gat));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n461), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G99gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n687), .A2(G99gat), .A3(new_n457), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n796), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(G1338gat));
  INV_X1    g626(.A(new_n738), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(G106gat), .A3(new_n283), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n796), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(KEYINPUT53), .ZN(new_n831));
  XNOR2_X1  g630(.A(KEYINPUT117), .B(G106gat), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n733), .A2(new_n283), .A3(new_n801), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n832), .B1(new_n806), .B2(new_n467), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT53), .B1(new_n835), .B2(new_n830), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(G1339gat));
  AOI21_X1  g636(.A(new_n677), .B1(new_n674), .B2(new_n675), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n664), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n678), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n683), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n838), .A2(new_n664), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n684), .ZN(new_n848));
  OR3_X1    g647(.A1(new_n845), .A2(KEYINPUT118), .A3(new_n846), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT118), .B1(new_n845), .B2(new_n846), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n735), .A2(new_n851), .A3(new_n736), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n576), .A2(new_n577), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n582), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT119), .Z(new_n856));
  AND2_X1   g655(.A1(new_n585), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n686), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n619), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n851), .A2(new_n619), .A3(new_n857), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n657), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n688), .A2(new_n737), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n774), .A2(new_n427), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n865), .A2(new_n529), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n372), .B1(new_n868), .B2(new_n592), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT120), .ZN(new_n870));
  INV_X1    g669(.A(new_n737), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n868), .A2(new_n372), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(G1340gat));
  AOI21_X1  g672(.A(G120gat), .B1(new_n868), .B2(new_n686), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n828), .A2(new_n373), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n868), .B2(new_n875), .ZN(G1341gat));
  NAND2_X1  g675(.A1(new_n868), .A2(new_n659), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(G127gat), .ZN(G1342gat));
  AOI21_X1  g677(.A(new_n365), .B1(new_n868), .B2(new_n619), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT121), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n709), .A2(new_n427), .A3(new_n493), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n864), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n524), .A2(new_n365), .ZN(new_n884));
  OR3_X1    g683(.A1(new_n883), .A2(KEYINPUT56), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT56), .B1(new_n883), .B2(new_n884), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n880), .B(new_n885), .C1(new_n888), .C2(new_n889), .ZN(G1343gat));
  NOR2_X1   g689(.A1(new_n867), .A2(new_n461), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n851), .A2(new_n592), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(KEYINPUT123), .A3(new_n858), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n709), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT123), .B1(new_n893), .B2(new_n858), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n860), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n657), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n892), .B(new_n283), .C1(new_n898), .C2(new_n863), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n283), .B1(new_n862), .B2(new_n863), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(KEYINPUT57), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n891), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G141gat), .B1(new_n902), .B2(new_n593), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n461), .A2(new_n283), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n864), .A2(new_n866), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n593), .A2(G141gat), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT58), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n871), .B(new_n891), .C1(new_n899), .C2(new_n901), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n909), .A2(G141gat), .B1(new_n905), .B2(new_n906), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1344gat));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n913), .B(G148gat), .C1(new_n902), .C2(new_n687), .ZN(new_n914));
  INV_X1    g713(.A(G148gat), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n897), .A2(new_n657), .B1(new_n593), .B2(new_n688), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n892), .B1(new_n916), .B2(new_n283), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n900), .A2(KEYINPUT124), .A3(KEYINPUT57), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT124), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n867), .A2(new_n461), .A3(new_n687), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n914), .B1(new_n913), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n915), .A3(new_n686), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1345gat));
  OAI21_X1  g724(.A(G155gat), .B1(new_n902), .B2(new_n657), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n905), .A2(new_n226), .A3(new_n659), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1346gat));
  OAI21_X1  g727(.A(G162gat), .B1(new_n902), .B2(new_n709), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n882), .A2(new_n227), .A3(new_n904), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n360), .A2(new_n707), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n781), .A2(new_n932), .A3(new_n283), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n865), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n327), .A3(new_n593), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n707), .B1(new_n862), .B2(new_n863), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(new_n524), .A3(new_n774), .ZN(new_n937));
  AOI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n871), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n935), .A2(new_n938), .ZN(G1348gat));
  OAI21_X1  g738(.A(G176gat), .B1(new_n934), .B2(new_n828), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n328), .A3(new_n686), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1349gat));
  OAI211_X1 g741(.A(new_n937), .B(new_n659), .C1(new_n300), .C2(new_n301), .ZN(new_n943));
  OAI21_X1  g742(.A(G183gat), .B1(new_n934), .B2(new_n657), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n937), .A2(new_n289), .A3(new_n619), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n948));
  OR3_X1    g747(.A1(new_n865), .A2(new_n709), .A3(new_n933), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(G190gat), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n949), .A2(new_n948), .A3(G190gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n952), .B1(new_n950), .B2(KEYINPUT125), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n947), .B1(new_n951), .B2(new_n953), .ZN(G1351gat));
  AND2_X1   g753(.A1(new_n904), .A2(new_n774), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(G197gat), .B1(new_n957), .B2(new_n871), .ZN(new_n958));
  INV_X1    g757(.A(new_n920), .ZN(new_n959));
  INV_X1    g758(.A(new_n932), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n960), .A2(new_n461), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n593), .A2(new_n206), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n958), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  NOR3_X1   g764(.A1(new_n956), .A2(G204gat), .A3(new_n687), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT62), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n959), .A2(new_n828), .A3(new_n962), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n204), .ZN(G1353gat));
  OR3_X1    g768(.A1(new_n956), .A2(G211gat), .A3(new_n657), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n920), .A2(new_n659), .A3(new_n961), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  AOI21_X1  g773(.A(G218gat), .B1(new_n957), .B2(new_n619), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n619), .A2(G218gat), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT126), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n975), .B1(new_n963), .B2(new_n977), .ZN(G1355gat));
endmodule


