//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(KEYINPUT22), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n203), .B1(new_n210), .B2(KEYINPUT29), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(KEYINPUT79), .A2(G155gat), .A3(G162gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G148gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G141gat), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G148gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT80), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G155gat), .B(G162gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n219), .A2(KEYINPUT80), .A3(G141gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  INV_X1    g027(.A(G162gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT81), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT81), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G162gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n228), .B1(new_n233), .B2(G155gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n218), .B1(new_n227), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n211), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n203), .B(new_n218), .C1(new_n227), .C2(new_n234), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n210), .B1(new_n238), .B2(KEYINPUT29), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G78gat), .B(G106gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G228gat), .A2(G233gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(G22gat), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT31), .B(G50gat), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n242), .B(new_n246), .Z(new_n247));
  XNOR2_X1  g046(.A(G8gat), .B(G36gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(G64gat), .B(G92gat), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n248), .B(new_n249), .Z(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G226gat), .ZN(new_n252));
  INV_X1    g051(.A(G233gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT70), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT26), .ZN(new_n257));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT65), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(G169gat), .A3(G176gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT26), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n257), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OR2_X1    g066(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n268));
  INV_X1    g067(.A(G183gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT27), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT27), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G183gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n268), .A2(new_n270), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT67), .B(G190gat), .Z(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT27), .B(G183gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n276), .B1(KEYINPUT69), .B2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n282));
  NAND2_X1  g081(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n267), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT64), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n255), .A2(KEYINPUT23), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n292), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(new_n288), .A3(new_n290), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n293), .A2(new_n297), .A3(new_n299), .A4(new_n262), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  AND4_X1   g100(.A1(KEYINPUT25), .A2(new_n262), .A3(new_n296), .A4(new_n294), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n303));
  OAI211_X1 g102(.A(G183gat), .B(G190gat), .C1(new_n303), .C2(KEYINPUT24), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n266), .A2(KEYINPUT66), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n268), .A2(new_n273), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n304), .B(new_n306), .C1(new_n307), .C2(G183gat), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n300), .A2(new_n301), .B1(new_n302), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n254), .B1(new_n286), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n210), .ZN(new_n311));
  INV_X1    g110(.A(new_n267), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n274), .A2(KEYINPUT69), .A3(new_n282), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n275), .B2(new_n274), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n280), .A2(KEYINPUT69), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n308), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT29), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n310), .B(new_n311), .C1(new_n320), .C2(new_n254), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n285), .B(new_n313), .C1(new_n275), .C2(new_n274), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n323), .A2(new_n312), .B1(new_n317), .B2(new_n318), .ZN(new_n324));
  OAI22_X1  g123(.A1(new_n324), .A2(KEYINPUT29), .B1(new_n252), .B2(new_n253), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n311), .B1(new_n325), .B2(new_n310), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n251), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n310), .B1(new_n320), .B2(new_n254), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n210), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(new_n250), .A3(new_n321), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(KEYINPUT30), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n329), .A2(new_n332), .A3(new_n250), .A4(new_n321), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT4), .ZN(new_n335));
  NOR2_X1   g134(.A1(G127gat), .A2(G134gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT71), .B(G127gat), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(G134gat), .ZN(new_n338));
  INV_X1    g137(.A(G113gat), .ZN(new_n339));
  INV_X1    g138(.A(G120gat), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT1), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n339), .B2(new_n340), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G127gat), .A2(G134gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n341), .B1(new_n345), .B2(new_n336), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G120gat), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n339), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n346), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(G113gat), .B2(G120gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n336), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n344), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n348), .A2(G120gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n358));
  OAI21_X1  g157(.A(G113gat), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT73), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n343), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n335), .B1(new_n361), .B2(new_n235), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n363), .A3(new_n237), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n351), .B1(new_n346), .B2(new_n350), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n356), .A2(new_n359), .A3(KEYINPUT73), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n365), .A2(new_n366), .B1(new_n342), .B2(new_n338), .ZN(new_n367));
  INV_X1    g166(.A(new_n235), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n362), .A2(new_n364), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT39), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n372), .A2(new_n375), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n361), .A2(new_n235), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n368), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT39), .B1(new_n387), .B2(new_n375), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n383), .B(KEYINPUT40), .C1(new_n384), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n369), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT4), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n390), .A2(new_n364), .A3(new_n374), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n375), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(KEYINPUT5), .A3(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n375), .A2(KEYINPUT5), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n362), .A2(new_n364), .A3(new_n371), .A4(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n396), .A2(new_n397), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n394), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n381), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT40), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n384), .A2(new_n388), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(new_n382), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n389), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n247), .B1(new_n334), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n330), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT37), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n329), .A2(new_n409), .A3(new_n321), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT38), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n329), .A2(new_n321), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n250), .B1(new_n413), .B2(KEYINPUT37), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n408), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT6), .B1(new_n400), .B2(new_n401), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n362), .A2(new_n364), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n417), .A2(KEYINPUT84), .A3(new_n371), .A4(new_n395), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n397), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n381), .A3(new_n394), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n381), .B1(new_n420), .B2(new_n394), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT85), .B1(new_n423), .B2(KEYINPUT6), .ZN(new_n424));
  AND4_X1   g223(.A1(KEYINPUT85), .A2(new_n400), .A3(KEYINPUT6), .A4(new_n401), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n415), .B(new_n422), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n410), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT37), .B1(new_n322), .B2(new_n326), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n251), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n429), .B2(KEYINPUT86), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n411), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n407), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n361), .A2(KEYINPUT74), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT74), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n367), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n435), .B(new_n437), .C1(new_n286), .C2(new_n309), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n316), .A2(new_n319), .A3(KEYINPUT74), .A4(new_n361), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT32), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n440), .B2(new_n441), .ZN(new_n444));
  XOR2_X1   g243(.A(G71gat), .B(G99gat), .Z(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT76), .ZN(new_n446));
  XNOR2_X1  g245(.A(G15gat), .B(G43gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT75), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n446), .B(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n442), .A2(new_n444), .A3(new_n450), .ZN(new_n451));
  OAI221_X1 g250(.A(KEYINPUT32), .B1(new_n443), .B2(new_n449), .C1(new_n440), .C2(new_n441), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT34), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n440), .A2(new_n454), .A3(new_n441), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT77), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT77), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n440), .A2(new_n457), .A3(new_n454), .A4(new_n441), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n441), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT34), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n454), .B1(new_n440), .B2(new_n441), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n440), .A2(new_n454), .A3(new_n441), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(new_n457), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n465), .A2(new_n456), .A3(new_n452), .A4(new_n451), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT36), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n462), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT78), .ZN(new_n469));
  INV_X1    g268(.A(new_n461), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n453), .A2(KEYINPUT78), .A3(new_n461), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n468), .B1(new_n473), .B2(KEYINPUT36), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n400), .A2(KEYINPUT6), .A3(new_n401), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n422), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n247), .B1(new_n477), .B2(new_n334), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n434), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT35), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n453), .A2(KEYINPUT78), .A3(new_n461), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n461), .B1(new_n453), .B2(KEYINPUT78), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n481), .A2(new_n482), .A3(new_n247), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n422), .A2(new_n475), .B1(new_n333), .B2(new_n331), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n475), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n400), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n401), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n487), .A2(new_n488), .B1(new_n421), .B2(new_n416), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT87), .B1(new_n489), .B2(new_n334), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n331), .A2(new_n333), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n462), .A2(new_n466), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n495), .A2(KEYINPUT35), .A3(new_n247), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT88), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n485), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n490), .A2(new_n494), .A3(new_n496), .A4(KEYINPUT88), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n479), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT92), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G1gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n505), .A2(KEYINPUT16), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n507), .B2(new_n504), .ZN(new_n508));
  INV_X1    g307(.A(G8gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT15), .ZN(new_n511));
  XNOR2_X1  g310(.A(G43gat), .B(G50gat), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(KEYINPUT90), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(KEYINPUT90), .B2(new_n512), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  AOI21_X1  g314(.A(G36gat), .B1(new_n515), .B2(G29gat), .ZN(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT14), .ZN(new_n518));
  MUX2_X1   g317(.A(G36gat), .B(new_n516), .S(new_n518), .Z(new_n519));
  OR2_X1    g318(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n521), .A2(KEYINPUT91), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(KEYINPUT91), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n522), .A2(new_n514), .A3(new_n519), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT17), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n508), .B(G8gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n525), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(KEYINPUT18), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n510), .A2(new_n526), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n534), .B(KEYINPUT13), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n530), .A2(new_n534), .A3(new_n532), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n535), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G169gat), .B(G197gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT12), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n549), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n535), .A2(new_n539), .A3(new_n542), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n202), .B1(new_n501), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n497), .A2(new_n498), .ZN(new_n556));
  INV_X1    g355(.A(new_n485), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n500), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n479), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(KEYINPUT93), .A3(new_n553), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT7), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  INV_X1    g366(.A(G92gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(KEYINPUT8), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G99gat), .B(G106gat), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n563), .B1(new_n526), .B2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n573), .B(KEYINPUT95), .Z(new_n574));
  NAND3_X1  g373(.A1(new_n527), .A2(new_n529), .A3(new_n572), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G134gat), .B(G162gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n576), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(new_n576), .B2(new_n579), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(KEYINPUT94), .A2(G57gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(G64gat), .Z(new_n590));
  NOR2_X1   g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT9), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(G57gat), .B2(G64gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n591), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n593), .ZN(new_n598));
  OAI22_X1  g397(.A1(new_n590), .A2(new_n594), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n603), .B(G127gat), .Z(new_n604));
  OAI21_X1  g403(.A(new_n510), .B1(new_n600), .B2(new_n599), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G155gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n588), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G120gat), .B(G148gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT97), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n572), .A2(new_n599), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n572), .A2(new_n599), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  OR3_X1    g422(.A1(new_n572), .A2(new_n621), .A3(new_n599), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT98), .ZN(new_n628));
  INV_X1    g427(.A(new_n626), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(new_n623), .B2(new_n624), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n620), .A2(new_n622), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n629), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n619), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n627), .A2(new_n635), .A3(new_n618), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n614), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n562), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n477), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g442(.A(KEYINPUT16), .B(G8gat), .Z(new_n644));
  AND3_X1   g443(.A1(new_n641), .A2(new_n334), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n509), .B1(new_n641), .B2(new_n334), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT42), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(KEYINPUT42), .B2(new_n645), .ZN(G1325gat));
  INV_X1    g447(.A(G15gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n495), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n641), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n474), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n641), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n651), .B1(new_n653), .B2(new_n649), .ZN(G1326gat));
  NAND2_X1  g453(.A1(new_n641), .A2(new_n247), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT43), .B(G22gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  AOI21_X1  g456(.A(new_n588), .B1(new_n558), .B2(new_n559), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT44), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661));
  NOR4_X1   g460(.A1(new_n501), .A2(KEYINPUT100), .A3(new_n661), .A4(new_n588), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n639), .B(KEYINPUT99), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n666), .A2(new_n554), .A3(new_n613), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n663), .A2(new_n664), .A3(new_n477), .A4(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n560), .A2(new_n659), .A3(new_n587), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n661), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT44), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n670), .A2(new_n477), .A3(new_n671), .A4(new_n667), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT101), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n668), .A2(new_n673), .A3(G29gat), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n588), .A2(new_n613), .A3(new_n639), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n562), .A2(new_n517), .A3(new_n477), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT45), .ZN(new_n677));
  INV_X1    g476(.A(new_n675), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n555), .B2(new_n561), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n517), .A4(new_n477), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n674), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n674), .A2(KEYINPUT102), .A3(new_n682), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(G1328gat));
  INV_X1    g486(.A(G36gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n679), .A2(new_n688), .A3(new_n334), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT46), .Z(new_n690));
  NAND3_X1  g489(.A1(new_n663), .A2(new_n334), .A3(new_n667), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G36gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n690), .B1(new_n693), .B2(new_n695), .ZN(G1329gat));
  NAND4_X1  g495(.A1(new_n670), .A2(new_n652), .A3(new_n671), .A4(new_n667), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G43gat), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n495), .A2(G43gat), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n562), .A2(new_n675), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT104), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n679), .A2(new_n702), .A3(new_n699), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n698), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT105), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n705), .A2(KEYINPUT105), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n706), .B1(new_n704), .B2(new_n707), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(G1330gat));
  NAND4_X1  g509(.A1(new_n670), .A2(new_n247), .A3(new_n671), .A4(new_n667), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G50gat), .ZN(new_n712));
  INV_X1    g511(.A(new_n247), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(G50gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n679), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n712), .A2(KEYINPUT48), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n712), .A2(KEYINPUT107), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n711), .B2(G50gat), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n679), .A2(new_n714), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n722));
  OAI21_X1  g521(.A(new_n716), .B1(new_n721), .B2(new_n722), .ZN(G1331gat));
  NOR4_X1   g522(.A1(new_n501), .A2(new_n553), .A3(new_n614), .A4(new_n665), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n477), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g525(.A1(new_n724), .A2(new_n334), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  AND2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(G1333gat));
  NAND2_X1  g530(.A1(new_n724), .A2(new_n652), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n495), .A2(G71gat), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n732), .A2(G71gat), .B1(new_n724), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g534(.A1(new_n724), .A2(new_n247), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g536(.A1(new_n613), .A2(new_n553), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n739));
  AND2_X1   g538(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n658), .B(new_n738), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n738), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n501), .A2(new_n588), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n743), .B2(new_n740), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(new_n639), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(new_n567), .A3(new_n477), .ZN(new_n746));
  INV_X1    g545(.A(new_n639), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n663), .A2(new_n477), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n746), .B1(new_n567), .B2(new_n749), .ZN(G1336gat));
  NAND3_X1  g549(.A1(new_n663), .A2(new_n334), .A3(new_n748), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G92gat), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n665), .A2(G92gat), .A3(new_n493), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n744), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT110), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n744), .A2(new_n757), .A3(new_n754), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n752), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT52), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT111), .A2(KEYINPUT52), .ZN(new_n761));
  AND2_X1   g560(.A1(KEYINPUT111), .A2(KEYINPUT52), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n752), .B(new_n755), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(G1337gat));
  INV_X1    g563(.A(G99gat), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n745), .A2(new_n765), .A3(new_n650), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n663), .A2(new_n652), .A3(new_n748), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(G1338gat));
  NAND3_X1  g567(.A1(new_n663), .A2(new_n247), .A3(new_n748), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n665), .A2(G106gat), .A3(new_n713), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n744), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n770), .B2(new_n772), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(G1339gat));
  INV_X1    g575(.A(new_n613), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n628), .A2(new_n778), .A3(new_n632), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n619), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n630), .A2(new_n778), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n623), .A2(new_n629), .A3(new_n624), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n781), .A2(KEYINPUT113), .A3(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n780), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n780), .A2(new_n787), .A3(KEYINPUT55), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n790), .A2(new_n553), .A3(new_n638), .A4(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n533), .A2(new_n534), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n537), .A2(new_n538), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n793), .B(new_n548), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n548), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT114), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n639), .A2(new_n552), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n587), .B1(new_n792), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n790), .A2(new_n638), .A3(new_n791), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n587), .A2(new_n798), .A3(new_n552), .A4(new_n796), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n777), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n640), .A2(new_n554), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n476), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n495), .A2(new_n334), .A3(new_n247), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(G113gat), .B1(new_n809), .B2(new_n554), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n806), .A2(new_n483), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(KEYINPUT116), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(KEYINPUT116), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n493), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n553), .A2(new_n339), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n812), .A2(new_n813), .B1(new_n817), .B2(new_n818), .ZN(G1340gat));
  OAI21_X1  g618(.A(G120gat), .B1(new_n809), .B2(new_n665), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(KEYINPUT117), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(KEYINPUT117), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n639), .A2(new_n347), .A3(new_n349), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n821), .A2(new_n822), .B1(new_n817), .B2(new_n823), .ZN(G1341gat));
  OAI21_X1  g623(.A(new_n337), .B1(new_n809), .B2(new_n777), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n777), .A2(new_n337), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n817), .B2(new_n826), .ZN(G1342gat));
  NOR2_X1   g626(.A1(new_n588), .A2(G134gat), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n493), .B(new_n828), .C1(new_n815), .C2(new_n816), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n829), .A2(KEYINPUT56), .ZN(new_n830));
  OAI21_X1  g629(.A(G134gat), .B1(new_n809), .B2(new_n588), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n829), .A2(new_n832), .A3(KEYINPUT56), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n829), .B2(KEYINPUT56), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n830), .B(new_n831), .C1(new_n833), .C2(new_n834), .ZN(G1343gat));
  NOR3_X1   g634(.A1(new_n652), .A2(new_n713), .A3(new_n334), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n806), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(G141gat), .A3(new_n554), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n652), .A2(new_n476), .A3(new_n334), .ZN(new_n839));
  XOR2_X1   g638(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n840));
  NAND2_X1  g639(.A1(new_n788), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n841), .A2(new_n553), .A3(new_n638), .A4(new_n791), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n587), .B1(new_n842), .B2(new_n799), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n777), .B1(new_n843), .B2(new_n803), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n713), .B1(new_n844), .B2(new_n805), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(KEYINPUT57), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n713), .B1(new_n804), .B2(new_n805), .ZN(new_n847));
  XNOR2_X1  g646(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n553), .B(new_n839), .C1(new_n846), .C2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n838), .B1(new_n851), .B2(G141gat), .ZN(new_n852));
  XOR2_X1   g651(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n853));
  XNOR2_X1  g652(.A(new_n852), .B(new_n853), .ZN(G1344gat));
  NOR3_X1   g653(.A1(new_n837), .A2(G148gat), .A3(new_n747), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT122), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n219), .A2(KEYINPUT59), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n839), .B1(new_n846), .B2(new_n850), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n747), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n804), .A2(new_n805), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n247), .A3(new_n849), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(KEYINPUT57), .B2(new_n845), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n864), .A2(new_n639), .A3(new_n839), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT59), .B1(new_n865), .B2(new_n219), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n859), .A2(new_n860), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n856), .B1(new_n867), .B2(new_n868), .ZN(G1345gat));
  OAI21_X1  g668(.A(G155gat), .B1(new_n858), .B2(new_n777), .ZN(new_n870));
  OR3_X1    g669(.A1(new_n837), .A2(G155gat), .A3(new_n777), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1346gat));
  OAI21_X1  g671(.A(new_n233), .B1(new_n858), .B2(new_n588), .ZN(new_n873));
  OR3_X1    g672(.A1(new_n837), .A2(new_n233), .A3(new_n588), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1347gat));
  NOR2_X1   g674(.A1(new_n477), .A2(new_n493), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n877), .B1(new_n804), .B2(new_n805), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n495), .A2(new_n247), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n881), .A2(G169gat), .A3(new_n553), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n878), .A2(new_n483), .ZN(new_n883));
  AOI21_X1  g682(.A(G169gat), .B1(new_n883), .B2(new_n553), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n884), .ZN(G1348gat));
  NAND3_X1  g684(.A1(new_n881), .A2(G176gat), .A3(new_n666), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT124), .ZN(new_n887));
  AOI21_X1  g686(.A(G176gat), .B1(new_n883), .B2(new_n639), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(G1349gat));
  NAND3_X1  g688(.A1(new_n883), .A2(new_n279), .A3(new_n613), .ZN(new_n890));
  OAI21_X1  g689(.A(G183gat), .B1(new_n880), .B2(new_n777), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g692(.A1(new_n883), .A2(new_n278), .A3(new_n587), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT125), .Z(new_n895));
  OAI21_X1  g694(.A(G190gat), .B1(new_n880), .B2(new_n588), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT61), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1351gat));
  NOR2_X1   g697(.A1(new_n652), .A2(new_n877), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n847), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(G197gat), .B1(new_n900), .B2(new_n553), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n863), .B(new_n902), .C1(KEYINPUT57), .C2(new_n845), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n903), .A2(new_n899), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n845), .A2(KEYINPUT57), .ZN(new_n905));
  AOI211_X1 g704(.A(new_n713), .B(new_n848), .C1(new_n804), .C2(new_n805), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT126), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n553), .A2(G197gat), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n901), .B1(new_n908), .B2(new_n909), .ZN(G1352gat));
  NAND3_X1  g709(.A1(new_n904), .A2(new_n666), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G204gat), .ZN(new_n912));
  INV_X1    g711(.A(G204gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n900), .A2(new_n913), .A3(new_n639), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT62), .Z(new_n915));
  NAND2_X1  g714(.A1(new_n912), .A2(new_n915), .ZN(G1353gat));
  NAND3_X1  g715(.A1(new_n864), .A2(new_n613), .A3(new_n899), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G211gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n900), .A2(new_n205), .A3(new_n613), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1354gat));
  NAND4_X1  g721(.A1(new_n907), .A2(new_n587), .A3(new_n903), .A4(new_n899), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G218gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n900), .A2(new_n206), .A3(new_n587), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT127), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n928), .A3(new_n925), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1355gat));
endmodule


