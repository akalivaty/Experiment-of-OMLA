//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT69), .B1(new_n461), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n461), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n462), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n468), .A2(G137), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(new_n466), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n464), .A2(G2105), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  NOR3_X1   g056(.A1(new_n475), .A2(new_n479), .A3(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n474), .A2(new_n467), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT70), .Z(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n464), .B1(new_n473), .B2(new_n486), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n483), .A2(G124), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n467), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n462), .A2(new_n465), .A3(new_n466), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n470), .A2(new_n472), .A3(G138), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n461), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n503), .A2(new_n506), .A3(new_n507), .A4(new_n462), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n470), .A2(new_n472), .A3(G138), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT72), .B1(new_n467), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(KEYINPUT4), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n476), .A2(new_n466), .ZN(new_n512));
  NOR3_X1   g087(.A1(new_n509), .A2(new_n512), .A3(KEYINPUT4), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n502), .B1(new_n511), .B2(new_n514), .ZN(G164));
  NAND2_X1  g090(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n517), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G50), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  AND3_X1   g103(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(G543), .B1(KEYINPUT73), .B2(KEYINPUT5), .ZN(new_n530));
  AND2_X1   g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n529), .A2(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n527), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n523), .A2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  NAND2_X1  g111(.A1(new_n526), .A2(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n518), .A2(new_n519), .B1(new_n524), .B2(new_n525), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n542), .A2(G89), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n522), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n526), .A2(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n548), .B2(new_n533), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  AOI22_X1  g125(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n522), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n542), .A2(G81), .B1(new_n526), .B2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  OAI21_X1  g135(.A(G65), .B1(new_n529), .B2(new_n530), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT77), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n561), .A2(new_n563), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n569), .A2(new_n570), .A3(G651), .A4(new_n564), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g147(.A(G53), .B(G543), .C1(new_n531), .C2(new_n532), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n573), .A2(KEYINPUT74), .A3(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n524), .A2(new_n525), .ZN(new_n575));
  NAND2_X1  g150(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n575), .A2(G53), .A3(G543), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n542), .B2(G91), .ZN(new_n580));
  INV_X1    g155(.A(G91), .ZN(new_n581));
  NOR3_X1   g156(.A1(new_n533), .A2(KEYINPUT75), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n578), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n572), .A2(new_n584), .ZN(G299));
  INV_X1    g160(.A(G171), .ZN(G301));
  INV_X1    g161(.A(G168), .ZN(G286));
  AOI22_X1  g162(.A1(new_n542), .A2(G87), .B1(new_n526), .B2(G49), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(new_n520), .A2(G61), .ZN(new_n591));
  INV_X1    g166(.A(G73), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(new_n517), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(new_n526), .B2(G48), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n542), .A2(G86), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n522), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n526), .A2(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n533), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n598), .A2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n533), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n526), .A2(KEYINPUT78), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(G54), .B1(new_n526), .B2(KEYINPUT78), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(new_n522), .ZN(new_n612));
  AND3_X1   g187(.A1(new_n606), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n603), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n603), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n583), .B1(new_n567), .B2(new_n571), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  INV_X1    g196(.A(new_n613), .ZN(new_n622));
  OAI21_X1  g197(.A(KEYINPUT79), .B1(new_n622), .B2(G559), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n613), .A2(new_n624), .A3(new_n620), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n623), .A2(G868), .A3(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n555), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(G282));
  INV_X1    g206(.A(new_n629), .ZN(G323));
  NAND3_X1  g207(.A1(new_n469), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT81), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n483), .A2(G123), .ZN(new_n639));
  OAI221_X1 g214(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n474), .C2(G111), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n489), .A2(G135), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n635), .A2(new_n636), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n638), .A2(new_n643), .A3(new_n645), .ZN(G156));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT83), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  XOR2_X1   g228(.A(G2443), .B(G2446), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n658), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT84), .ZN(new_n664));
  INV_X1    g239(.A(G14), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n665), .B1(new_n666), .B2(new_n661), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n671), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(KEYINPUT85), .ZN(new_n677));
  INV_X1    g252(.A(new_n670), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n674), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n678), .B1(new_n677), .B2(new_n671), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n677), .ZN(new_n684));
  OAI22_X1  g259(.A1(new_n681), .A2(new_n682), .B1(new_n684), .B2(new_n676), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n680), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G2096), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT88), .B(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n691), .A2(new_n696), .A3(new_n694), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n691), .A2(new_n696), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n699));
  AOI211_X1 g274(.A(new_n695), .B(new_n697), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n698), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G24), .ZN(new_n710));
  INV_X1    g285(.A(G290), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  INV_X1    g287(.A(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  OAI221_X1 g289(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n474), .C2(G107), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT91), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(KEYINPUT91), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n716), .A2(new_n717), .B1(G119), .B2(new_n483), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n489), .A2(G131), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(KEYINPUT90), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(KEYINPUT90), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G25), .B2(new_n726), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  OAI21_X1  g304(.A(new_n714), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n729), .B2(new_n728), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n709), .A2(G6), .ZN(new_n732));
  INV_X1    g307(.A(G305), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n709), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT32), .B(G1981), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n709), .A2(G22), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G166), .B2(new_n709), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1971), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n709), .A2(G23), .ZN(new_n740));
  INV_X1    g315(.A(G288), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(new_n709), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT33), .B(G1976), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n742), .B(new_n743), .Z(new_n744));
  NOR3_X1   g319(.A1(new_n736), .A2(new_n739), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT34), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n731), .A2(KEYINPUT93), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n731), .A2(new_n747), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT92), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT24), .B(G34), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n726), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT98), .Z(new_n756));
  INV_X1    g331(.A(G160), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n722), .ZN(new_n758));
  INV_X1    g333(.A(G2084), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT95), .B(G1341), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n709), .A2(G19), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(KEYINPUT94), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(KEYINPUT94), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n763), .B(new_n764), .C1(new_n555), .C2(new_n709), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n760), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n758), .A2(new_n759), .ZN(new_n767));
  NOR2_X1   g342(.A1(G168), .A2(new_n709), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n709), .B2(G21), .ZN(new_n769));
  INV_X1    g344(.A(G1966), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT31), .B(G11), .Z(new_n772));
  NOR2_X1   g347(.A1(new_n642), .A2(new_n726), .ZN(new_n773));
  INV_X1    g348(.A(G28), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(KEYINPUT30), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT100), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n774), .B2(KEYINPUT30), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n772), .B(new_n773), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n769), .A2(new_n770), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n767), .A2(new_n771), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n766), .B(new_n780), .C1(new_n761), .C2(new_n765), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n709), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n709), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1961), .ZN(new_n784));
  NOR2_X1   g359(.A1(G4), .A2(G16), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n613), .B2(G16), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT29), .B(G2090), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n726), .A2(G35), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT102), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n491), .B2(new_n725), .ZN(new_n790));
  OAI22_X1  g365(.A1(new_n786), .A2(G1348), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  AOI211_X1 g366(.A(new_n784), .B(new_n791), .C1(new_n787), .C2(new_n790), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n786), .A2(G1348), .ZN(new_n793));
  INV_X1    g368(.A(G2072), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n722), .A2(G33), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT25), .Z(new_n797));
  NAND2_X1  g372(.A1(G115), .A2(G2104), .ZN(new_n798));
  INV_X1    g373(.A(G127), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n512), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(new_n473), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT97), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n489), .A2(G139), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n797), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n795), .B1(new_n804), .B2(G29), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n793), .B1(new_n794), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n794), .B2(new_n805), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n781), .A2(new_n792), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n709), .A2(G20), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT23), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n617), .B2(new_n709), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1956), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n722), .A2(G32), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n489), .A2(G141), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT99), .ZN(new_n815));
  NAND3_X1  g390(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT26), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n480), .A2(G105), .ZN(new_n818));
  AOI211_X1 g393(.A(new_n817), .B(new_n818), .C1(new_n483), .C2(G129), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n813), .B1(new_n821), .B2(new_n722), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT27), .B(G1996), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n725), .A2(G27), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G164), .B2(new_n725), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT101), .B(G2078), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n726), .A2(G26), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n483), .A2(G128), .ZN(new_n832));
  OAI221_X1 g407(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n474), .C2(G116), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G140), .B2(new_n489), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n831), .B1(new_n835), .B2(new_n722), .ZN(new_n836));
  INV_X1    g411(.A(G2067), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n824), .A2(new_n828), .A3(new_n838), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n808), .A2(new_n812), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n751), .A2(new_n753), .A3(new_n840), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n749), .A2(KEYINPUT92), .A3(new_n750), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(G311));
  INV_X1    g418(.A(G311), .ZN(G150));
  AOI22_X1  g419(.A1(new_n542), .A2(G93), .B1(new_n526), .B2(G55), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n522), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(KEYINPUT103), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(KEYINPUT103), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n555), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n554), .A2(new_n847), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n613), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n856), .A2(new_n857), .A3(G860), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n848), .A2(new_n849), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT37), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n858), .A2(new_n861), .ZN(G145));
  NAND2_X1  g437(.A1(new_n511), .A2(new_n514), .ZN(new_n863));
  INV_X1    g438(.A(new_n501), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n498), .A2(new_n499), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n495), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n835), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n820), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n804), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n720), .A2(new_n634), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n720), .A2(new_n634), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n483), .A2(G130), .ZN(new_n874));
  OAI221_X1 g449(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n474), .C2(G118), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n489), .A2(G142), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n871), .B2(new_n872), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(KEYINPUT104), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n870), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(G160), .B(new_n491), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n642), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n885), .B(new_n887), .C1(new_n870), .C2(new_n882), .ZN(new_n888));
  XOR2_X1   g463(.A(KEYINPUT105), .B(G37), .Z(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n881), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n870), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n888), .B(new_n889), .C1(new_n891), .C2(new_n887), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g468(.A1(G299), .A2(new_n613), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT106), .B1(G299), .B2(new_n613), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n613), .B(new_n617), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n898), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n623), .A2(new_n625), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n850), .A2(new_n851), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  MUX2_X1   g482(.A(new_n903), .B(new_n904), .S(new_n907), .Z(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n711), .B(G305), .ZN(new_n910));
  XNOR2_X1  g485(.A(G303), .B(new_n741), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n909), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n909), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(G868), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n859), .A2(new_n627), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(G295));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n918), .ZN(G331));
  INV_X1    g495(.A(new_n904), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n922));
  XNOR2_X1  g497(.A(G171), .B(G168), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n852), .B2(new_n924), .ZN(new_n925));
  NOR4_X1   g500(.A1(new_n850), .A2(new_n923), .A3(KEYINPUT109), .A4(new_n851), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n923), .B1(new_n850), .B2(new_n851), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n906), .A2(KEYINPUT108), .A3(new_n923), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n921), .A2(new_n927), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n852), .A2(new_n924), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n928), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n899), .A2(new_n902), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n936), .B2(new_n913), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n912), .B1(new_n932), .B2(new_n935), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT110), .B1(new_n941), .B2(G37), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n932), .A2(new_n935), .A3(new_n912), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n939), .A2(new_n940), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT111), .ZN(new_n945));
  INV_X1    g520(.A(new_n943), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n937), .B2(new_n938), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n940), .A4(new_n942), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n931), .B(new_n930), .C1(new_n925), .C2(new_n926), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n901), .B2(new_n900), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n904), .B1(new_n952), .B2(new_n934), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n901), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n913), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n889), .A3(new_n943), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n950), .B1(new_n956), .B2(KEYINPUT43), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n945), .A2(new_n949), .A3(new_n957), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n959));
  AOI21_X1  g534(.A(new_n940), .B1(new_n947), .B2(new_n942), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(G397));
  XOR2_X1   g538(.A(new_n720), .B(new_n729), .Z(new_n964));
  INV_X1    g539(.A(G1996), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n820), .B(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n835), .B(G2067), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(G164), .B2(G1384), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT112), .B(G40), .ZN(new_n972));
  NOR4_X1   g547(.A1(new_n475), .A2(new_n479), .A3(new_n481), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n969), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n711), .A2(new_n713), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT113), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n713), .B2(new_n711), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n977), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT114), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n867), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n971), .A2(new_n973), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n770), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT4), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n467), .A2(new_n509), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n989), .B2(new_n507), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n513), .B1(new_n990), .B2(new_n510), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n984), .B1(new_n991), .B2(new_n502), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n974), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n863), .B2(new_n866), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n759), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n987), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT116), .B(G8), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G168), .A2(new_n999), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(KEYINPUT51), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G8), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n987), .B2(new_n997), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT51), .B1(new_n1006), .B2(new_n1002), .ZN(new_n1007));
  AOI211_X1 g582(.A(G168), .B(new_n999), .C1(new_n987), .C2(new_n997), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G2078), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n867), .B2(new_n984), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n970), .B(G1384), .C1(new_n863), .C2(new_n866), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT115), .B1(new_n1013), .B2(new_n973), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n971), .A2(KEYINPUT115), .A3(new_n985), .A4(new_n973), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1010), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n973), .B1(new_n994), .B2(new_n995), .ZN(new_n1020));
  NOR3_X1   g595(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1022), .A2(G1961), .ZN(new_n1023));
  AND2_X1   g598(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1024));
  NOR2_X1   g599(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT53), .B(G40), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n757), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1013), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1019), .A2(G301), .A3(new_n1023), .A4(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1013), .A2(KEYINPUT53), .A3(new_n1010), .A4(new_n973), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n986), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(G2078), .B1(new_n1032), .B2(new_n1015), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1023), .B(new_n1030), .C1(new_n1033), .C2(KEYINPUT53), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G171), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1029), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1009), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1971), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1032), .A2(new_n1039), .A3(new_n1015), .ZN(new_n1040));
  INV_X1    g615(.A(G2090), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1022), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n1000), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G303), .A2(G8), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT55), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n999), .B1(new_n994), .B2(new_n973), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n741), .A2(G1976), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT52), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G305), .A2(G1981), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1981), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT117), .B(G86), .Z(new_n1055));
  NAND2_X1  g630(.A1(new_n542), .A2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n594), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1053), .B(KEYINPUT49), .C1(new_n1054), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT49), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1057), .A2(new_n1054), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n1052), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1048), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n741), .B2(G1976), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1051), .B(new_n1062), .C1(new_n1050), .C2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1005), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1046), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1047), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT125), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1047), .A2(new_n1068), .A3(KEYINPUT125), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1023), .B(new_n1028), .C1(new_n1033), .C2(KEYINPUT53), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1074), .B(KEYINPUT54), .C1(G171), .C2(new_n1034), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1038), .A2(new_n1071), .A3(new_n1072), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1956), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n617), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  NOR2_X1   g657(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n617), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT56), .B(G2072), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n971), .A2(new_n973), .A3(new_n985), .A4(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1078), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1078), .A2(new_n1087), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1085), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT122), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1085), .B1(new_n1078), .B2(new_n1087), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n992), .B2(new_n974), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n994), .A2(KEYINPUT121), .A3(new_n973), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n837), .ZN(new_n1102));
  INV_X1    g677(.A(G1348), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n613), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1089), .B1(new_n1097), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n613), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1102), .A2(new_n1104), .A3(KEYINPUT60), .A4(new_n622), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1109), .A2(new_n1110), .B1(new_n1108), .B2(new_n1105), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1088), .A2(KEYINPUT61), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1093), .A2(new_n1112), .A3(new_n1096), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT58), .B(G1341), .Z(new_n1114));
  NAND3_X1  g689(.A1(new_n1099), .A2(new_n1100), .A3(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n971), .A2(new_n965), .A3(new_n985), .A4(new_n973), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n554), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1117), .B(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1113), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1111), .B1(new_n1122), .B2(KEYINPUT123), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1113), .A2(new_n1119), .A3(new_n1124), .A4(new_n1121), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1107), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1076), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1004), .B(KEYINPUT62), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1128), .A2(G171), .A3(new_n1034), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1009), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1129), .A2(new_n1071), .A3(new_n1072), .A4(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n1133));
  NAND3_X1  g708(.A1(new_n998), .A2(G168), .A3(new_n1000), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(new_n1069), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1065), .B(KEYINPUT118), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT63), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1137), .ZN(new_n1143));
  INV_X1    g718(.A(G1976), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1062), .A2(new_n1144), .A3(new_n741), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1053), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1136), .A2(new_n1143), .B1(new_n1048), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1132), .A2(new_n1142), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n983), .B1(new_n1127), .B2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n977), .B(KEYINPUT126), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n979), .A2(new_n975), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT48), .Z(new_n1152));
  AND4_X1   g727(.A1(new_n729), .A2(new_n966), .A3(new_n721), .A4(new_n967), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n837), .B2(new_n835), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1150), .A2(new_n1152), .B1(new_n976), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n976), .B1(new_n821), .B2(new_n967), .ZN(new_n1156));
  OR3_X1    g731(.A1(new_n976), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT46), .B1(new_n976), .B2(G1996), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT47), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1149), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g737(.A(G319), .ZN(new_n1164));
  NOR2_X1   g738(.A1(G227), .A2(new_n1164), .ZN(new_n1165));
  XOR2_X1   g739(.A(new_n1165), .B(KEYINPUT127), .Z(new_n1166));
  AND3_X1   g740(.A1(new_n668), .A2(new_n1166), .A3(new_n707), .ZN(new_n1167));
  OAI211_X1 g741(.A(new_n892), .B(new_n1167), .C1(new_n960), .C2(new_n961), .ZN(G225));
  INV_X1    g742(.A(G225), .ZN(G308));
endmodule


