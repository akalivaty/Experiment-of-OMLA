//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(KEYINPUT22), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n203), .B1(new_n210), .B2(KEYINPUT29), .ZN(new_n211));
  XOR2_X1   g010(.A(KEYINPUT75), .B(G155gat), .Z(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT2), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G155gat), .B(G162gat), .Z(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n216), .A2(KEYINPUT2), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n215), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n211), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n202), .B1(new_n222), .B2(KEYINPUT78), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n214), .A2(new_n217), .B1(new_n219), .B2(new_n215), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT29), .B1(new_n224), .B2(new_n203), .ZN(new_n225));
  INV_X1    g024(.A(new_n210), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  OAI221_X1 g027(.A(new_n222), .B1(KEYINPUT78), .B2(new_n202), .C1(new_n225), .C2(new_n226), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT79), .B(G22gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G78gat), .B(G106gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT31), .B(G50gat), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n233), .B(new_n234), .Z(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT77), .Z(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(G22gat), .A3(new_n229), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n230), .B2(new_n231), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n232), .A2(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G1gat), .B(G29gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT0), .ZN(new_n241));
  XNOR2_X1  g040(.A(G57gat), .B(G85gat), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n241), .B(new_n242), .Z(new_n243));
  INV_X1    g042(.A(KEYINPUT76), .ZN(new_n244));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245));
  XOR2_X1   g044(.A(G113gat), .B(G120gat), .Z(new_n246));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n246), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n246), .A2(KEYINPUT68), .A3(new_n245), .A4(new_n249), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(KEYINPUT4), .A3(new_n224), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT4), .B1(new_n254), .B2(new_n224), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n244), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(KEYINPUT76), .A3(new_n255), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n254), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n224), .A2(new_n203), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G225gat), .A2(G233gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n266), .A2(KEYINPUT5), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n259), .A2(new_n265), .A3(new_n267), .A4(new_n255), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n262), .A2(new_n221), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n224), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n271), .B(KEYINPUT5), .C1(new_n274), .C2(new_n267), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n243), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n270), .A2(new_n243), .A3(new_n275), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(KEYINPUT6), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT73), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(new_n289), .B2(new_n288), .ZN(new_n291));
  NOR2_X1   g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT23), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT25), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n287), .B1(new_n301), .B2(KEYINPUT24), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n301), .A2(KEYINPUT24), .ZN(new_n303));
  OAI221_X1 g102(.A(new_n288), .B1(G183gat), .B2(G190gat), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  AND4_X1   g103(.A1(KEYINPUT25), .A2(new_n293), .A3(new_n294), .A4(new_n296), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT66), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n308), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n292), .A2(KEYINPUT26), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT26), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n294), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n314), .B(new_n287), .C1(new_n316), .C2(new_n292), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n312), .B1(new_n309), .B2(new_n310), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(KEYINPUT28), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n307), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n285), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n300), .A2(new_n306), .B1(new_n313), .B2(new_n319), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(new_n284), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n210), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(KEYINPUT74), .A3(new_n285), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n328));
  INV_X1    g127(.A(new_n285), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n328), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n284), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n327), .A2(new_n330), .A3(new_n331), .A4(new_n226), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G8gat), .B(G36gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G64gat), .B(G92gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n334), .B(new_n335), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n326), .A2(new_n332), .A3(new_n336), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n338), .A2(KEYINPUT30), .A3(new_n339), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n333), .A2(KEYINPUT30), .A3(new_n337), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n239), .B1(new_n283), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n243), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n266), .B1(new_n258), .B2(new_n260), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(new_n267), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT39), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n272), .A2(new_n267), .A3(new_n273), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI221_X1 g150(.A(new_n351), .B1(new_n350), .B2(new_n349), .C1(new_n345), .C2(new_n267), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT40), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(KEYINPUT81), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n342), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n357), .B1(new_n348), .B2(new_n352), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n277), .B1(new_n358), .B2(new_n354), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n239), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n276), .A2(new_n362), .A3(KEYINPUT6), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n276), .B2(KEYINPUT6), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n280), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n339), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT37), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n336), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n338), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n329), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n324), .B2(new_n284), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n367), .B1(new_n374), .B2(new_n226), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n327), .A2(new_n330), .A3(new_n331), .A4(new_n210), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n366), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n368), .B1(new_n333), .B2(new_n337), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n367), .B1(new_n326), .B2(new_n332), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n372), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n361), .B1(new_n365), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n343), .B1(new_n360), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT69), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n324), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n313), .A2(new_n319), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n298), .A2(new_n299), .B1(new_n304), .B2(new_n305), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT69), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n386), .A2(new_n262), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n321), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT32), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(new_n392), .B2(new_n393), .ZN(new_n396));
  XOR2_X1   g195(.A(KEYINPUT70), .B(G71gat), .Z(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G99gat), .ZN(new_n398));
  XOR2_X1   g197(.A(G15gat), .B(G43gat), .Z(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n394), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  OAI221_X1 g201(.A(KEYINPUT32), .B1(new_n395), .B2(new_n400), .C1(new_n392), .C2(new_n393), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n390), .A2(new_n391), .B1(G227gat), .B2(G233gat), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT34), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n405), .A2(KEYINPUT72), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT72), .B1(new_n405), .B2(new_n406), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n405), .A2(new_n406), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT71), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n404), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n405), .A2(new_n406), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT72), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n405), .A2(KEYINPUT72), .A3(new_n406), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n405), .A2(new_n406), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n418), .A2(KEYINPUT71), .A3(new_n402), .A4(new_n403), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n412), .A2(KEYINPUT36), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n410), .A2(new_n402), .A3(new_n403), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT36), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n418), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n384), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n410), .A2(new_n404), .A3(new_n411), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n418), .A2(KEYINPUT71), .B1(new_n402), .B2(new_n403), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n361), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT84), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n283), .A2(new_n342), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n419), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(KEYINPUT84), .A3(new_n361), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT35), .ZN(new_n436));
  INV_X1    g235(.A(new_n342), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n437), .A2(new_n361), .A3(new_n421), .A4(new_n423), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT35), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n365), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n426), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G229gat), .A2(G233gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n444), .B(KEYINPUT88), .Z(new_n445));
  XOR2_X1   g244(.A(new_n445), .B(KEYINPUT13), .Z(new_n446));
  XNOR2_X1  g245(.A(G15gat), .B(G22gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT87), .ZN(new_n448));
  INV_X1    g247(.A(G1gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n447), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n449), .A2(KEYINPUT16), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(G8gat), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n450), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G43gat), .B(G50gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT15), .ZN(new_n458));
  NAND2_X1  g257(.A1(G29gat), .A2(G36gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT86), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n459), .A2(KEYINPUT86), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  OR3_X1    g261(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(KEYINPUT15), .B2(new_n457), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(KEYINPUT85), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT85), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n469), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n458), .B1(new_n471), .B2(new_n459), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n455), .B1(new_n450), .B2(new_n454), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n456), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n467), .A2(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n450), .A2(new_n454), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(G8gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n450), .A2(new_n454), .A3(new_n455), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n446), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n471), .A2(new_n459), .ZN(new_n482));
  OAI221_X1 g281(.A(KEYINPUT17), .B1(new_n462), .B2(new_n466), .C1(new_n482), .C2(new_n458), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT17), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n467), .B2(new_n472), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n478), .A2(new_n483), .A3(new_n479), .A4(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n473), .B1(new_n456), .B2(new_n474), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT18), .A4(new_n445), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n487), .A3(new_n445), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT18), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n493));
  XNOR2_X1  g292(.A(G113gat), .B(G141gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(G197gat), .ZN(new_n495));
  XOR2_X1   g294(.A(KEYINPUT11), .B(G169gat), .Z(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n497), .B(KEYINPUT12), .Z(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n489), .B(new_n492), .C1(new_n493), .C2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n488), .A3(new_n493), .ZN(new_n501));
  INV_X1    g300(.A(new_n492), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n481), .A2(new_n488), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n501), .B(new_n498), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n443), .A2(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G57gat), .B(G64gat), .Z(new_n508));
  INV_X1    g307(.A(G71gat), .ZN(new_n509));
  INV_X1    g308(.A(G78gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n508), .B1(KEYINPUT9), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(new_n509), .A3(new_n510), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT90), .B1(G71gat), .B2(G78gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n511), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n516), .A2(KEYINPUT91), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT91), .B1(new_n516), .B2(new_n517), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n512), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n509), .A2(new_n510), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n508), .A2(KEYINPUT9), .A3(new_n517), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G231gat), .A2(G233gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(G127gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n456), .A2(new_n474), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n525), .B2(new_n524), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n531), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(G155gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(new_n537), .Z(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n532), .A2(new_n533), .A3(new_n538), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT8), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n545));
  INV_X1    g344(.A(G85gat), .ZN(new_n546));
  INV_X1    g345(.A(G92gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n545), .B1(new_n544), .B2(new_n548), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n554), .A2(G85gat), .A3(G92gat), .A4(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n552), .B(new_n553), .C1(new_n546), .C2(new_n547), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT95), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(G99gat), .B(G106gat), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n548), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT94), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n556), .A2(new_n557), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n559), .A2(new_n560), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n560), .B1(new_n559), .B2(new_n567), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n483), .B(new_n485), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n560), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n551), .A2(KEYINPUT95), .A3(new_n558), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n566), .B1(new_n564), .B2(new_n565), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n560), .A3(new_n567), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n473), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n570), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(KEYINPUT96), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT96), .B1(new_n578), .B2(new_n579), .ZN(new_n582));
  INV_X1    g381(.A(new_n579), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n570), .A2(new_n583), .A3(new_n576), .A4(new_n577), .ZN(new_n584));
  XNOR2_X1  g383(.A(G134gat), .B(G162gat), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g387(.A1(new_n581), .A2(new_n582), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n587), .B(KEYINPUT92), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n578), .A2(new_n579), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n591), .B1(new_n592), .B2(new_n584), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT97), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n595));
  INV_X1    g394(.A(new_n593), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n582), .A2(new_n588), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(new_n581), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n542), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n524), .B1(new_n568), .B2(new_n569), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n574), .A2(new_n575), .A3(new_n523), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n574), .A2(KEYINPUT10), .A3(new_n575), .A4(new_n523), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G230gat), .ZN(new_n607));
  INV_X1    g406(.A(G233gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n610), .B1(new_n601), .B2(new_n603), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G120gat), .B(G148gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT98), .ZN(new_n615));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n611), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n609), .B1(new_n604), .B2(new_n605), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n617), .B1(new_n620), .B2(new_n612), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(KEYINPUT99), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT99), .B1(new_n619), .B2(new_n621), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n600), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n507), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n282), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n449), .ZN(G1324gat));
  NAND3_X1  g429(.A1(new_n507), .A2(new_n342), .A3(new_n627), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT16), .B(G8gat), .Z(new_n632));
  AND2_X1   g431(.A1(new_n632), .A2(KEYINPUT42), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OR3_X1    g433(.A1(new_n631), .A2(KEYINPUT102), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT102), .B1(new_n631), .B2(new_n634), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(G8gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT101), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n631), .A2(new_n640), .A3(G8gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT42), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n632), .B(KEYINPUT100), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n631), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n637), .A2(new_n642), .A3(new_n645), .ZN(G1325gat));
  INV_X1    g445(.A(new_n425), .ZN(new_n647));
  OAI21_X1  g446(.A(G15gat), .B1(new_n628), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n421), .A2(new_n423), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n650), .A2(G15gat), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n648), .B1(new_n628), .B2(new_n651), .ZN(G1326gat));
  OAI21_X1  g451(.A(KEYINPUT103), .B1(new_n628), .B2(new_n361), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n507), .A2(new_n654), .A3(new_n239), .A4(new_n627), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT43), .B(G22gat), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n653), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n653), .B2(new_n655), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(G1327gat));
  INV_X1    g458(.A(new_n542), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n625), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n599), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n441), .B1(new_n435), .B2(KEYINPUT35), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n505), .B(new_n662), .C1(new_n663), .C2(new_n426), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(G29gat), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n666), .A3(new_n283), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT45), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n661), .A2(new_n506), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT44), .B1(new_n443), .B2(new_n599), .ZN(new_n671));
  INV_X1    g470(.A(new_n599), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n384), .B2(new_n425), .ZN(new_n675));
  OAI221_X1 g474(.A(new_n361), .B1(new_n365), .B2(new_n382), .C1(new_n356), .C2(new_n359), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n676), .A2(new_n647), .A3(KEYINPUT104), .A4(new_n343), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n672), .B(new_n673), .C1(new_n678), .C2(new_n663), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n670), .B1(new_n671), .B2(new_n679), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n680), .A2(new_n283), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n668), .B1(new_n666), .B2(new_n681), .ZN(G1328gat));
  NOR2_X1   g481(.A1(new_n437), .A2(G36gat), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n665), .A2(KEYINPUT106), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n686));
  INV_X1    g485(.A(new_n683), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n664), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT107), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n684), .A2(new_n691), .A3(new_n685), .A4(new_n688), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n685), .B1(new_n684), .B2(new_n688), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n680), .A2(new_n342), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(G36gat), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(G1329gat));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698));
  INV_X1    g497(.A(G43gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n649), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n664), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n698), .B1(new_n701), .B2(KEYINPUT108), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n699), .B1(new_n680), .B2(new_n425), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n701), .ZN(new_n705));
  INV_X1    g504(.A(new_n701), .ZN(new_n706));
  AOI211_X1 g505(.A(new_n647), .B(new_n670), .C1(new_n671), .C2(new_n679), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n706), .B(new_n702), .C1(new_n707), .C2(new_n699), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(G1330gat));
  INV_X1    g508(.A(G50gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n239), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n664), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n680), .A2(new_n239), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(G50gat), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n715));
  AOI21_X1  g514(.A(new_n710), .B1(new_n680), .B2(new_n239), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n712), .A2(KEYINPUT110), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n664), .B2(new_n711), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(KEYINPUT48), .A3(new_n719), .ZN(new_n720));
  OAI22_X1  g519(.A1(new_n714), .A2(new_n715), .B1(new_n716), .B2(new_n720), .ZN(G1331gat));
  NOR2_X1   g520(.A1(new_n678), .A2(new_n663), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n600), .A2(new_n505), .A3(new_n625), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n283), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n342), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT49), .B(G64gat), .Z(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(G1333gat));
  NAND3_X1  g530(.A1(new_n725), .A2(new_n509), .A3(new_n649), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT84), .B1(new_n433), .B2(new_n361), .ZN(new_n733));
  AOI211_X1 g532(.A(new_n430), .B(new_n239), .C1(new_n412), .C2(new_n419), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n439), .B1(new_n735), .B2(new_n432), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n675), .B(new_n677), .C1(new_n736), .C2(new_n441), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(new_n425), .A3(new_n723), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n732), .B1(new_n509), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n239), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT111), .B(G78gat), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n743), .B(new_n744), .Z(G1335gat));
  NOR2_X1   g544(.A1(new_n542), .A2(new_n505), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n626), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n671), .B2(new_n679), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749), .B2(new_n282), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n672), .B(new_n746), .C1(new_n678), .C2(new_n663), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n737), .A2(KEYINPUT51), .A3(new_n672), .A4(new_n746), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT112), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n753), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n626), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n283), .A2(new_n546), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n750), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  AOI21_X1  g560(.A(new_n547), .B1(new_n748), .B2(new_n342), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n625), .A2(new_n437), .A3(G92gat), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n753), .B2(new_n754), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n755), .A2(new_n763), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  AOI211_X1 g567(.A(new_n437), .B(new_n747), .C1(new_n671), .C2(new_n679), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n767), .B(new_n768), .C1(new_n547), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(G1337gat));
  OAI21_X1  g570(.A(G99gat), .B1(new_n749), .B2(new_n647), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n650), .A2(G99gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n759), .B2(new_n773), .ZN(G1338gat));
  XNOR2_X1  g573(.A(KEYINPUT113), .B(G106gat), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n748), .B2(new_n239), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n625), .A2(new_n361), .A3(G106gat), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT114), .Z(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n753), .B2(new_n754), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT53), .B1(new_n776), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n755), .A2(new_n778), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n361), .B(new_n747), .C1(new_n671), .C2(new_n679), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n775), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n785), .ZN(G1339gat));
  NAND3_X1  g585(.A1(new_n489), .A2(new_n492), .A3(new_n499), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n475), .A2(new_n480), .A3(new_n446), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n445), .B1(new_n486), .B2(new_n487), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n497), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n623), .B2(new_n624), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n611), .A2(KEYINPUT54), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n618), .B1(new_n620), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT55), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(KEYINPUT55), .A3(new_n797), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n505), .A2(new_n799), .A3(new_n619), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n793), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n599), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n804), .A2(new_n620), .A3(new_n796), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n606), .A2(new_n796), .A3(new_n610), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n617), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n803), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n594), .A2(new_n598), .A3(new_n792), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n799), .A2(new_n619), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n802), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n660), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n542), .A2(new_n506), .A3(new_n599), .A4(new_n625), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n282), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n438), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n506), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n733), .A2(new_n734), .A3(new_n342), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n506), .A2(G113gat), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n819), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT115), .ZN(G1340gat));
  OAI21_X1  g624(.A(G120gat), .B1(new_n818), .B2(new_n625), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n625), .A2(G120gat), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(KEYINPUT116), .Z(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n821), .B2(new_n828), .ZN(G1341gat));
  OAI21_X1  g628(.A(G127gat), .B1(new_n818), .B2(new_n660), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n660), .A2(G127gat), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n821), .B2(new_n831), .ZN(G1342gat));
  OR3_X1    g631(.A1(new_n821), .A2(G134gat), .A3(new_n599), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n835));
  OAI21_X1  g634(.A(G134gat), .B1(new_n818), .B2(new_n599), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(G1343gat));
  NAND2_X1  g636(.A1(new_n647), .A2(new_n239), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n437), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n816), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n842), .A2(G141gat), .A3(new_n506), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n283), .A2(new_n437), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n425), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n814), .A2(new_n815), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n846), .B2(new_n239), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n808), .A2(KEYINPUT117), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n798), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n793), .B1(new_n851), .B2(new_n800), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n811), .B1(new_n852), .B2(new_n599), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n815), .B1(new_n853), .B2(new_n542), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n361), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n845), .B1(new_n847), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(G141gat), .B1(new_n859), .B2(new_n506), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g660(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n862), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n843), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(G1344gat));
  INV_X1    g665(.A(new_n842), .ZN(new_n867));
  INV_X1    g666(.A(G148gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n626), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n542), .B1(new_n802), .B2(new_n812), .ZN(new_n871));
  INV_X1    g670(.A(new_n815), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n856), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n799), .A2(new_n619), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n874), .A2(new_n848), .A3(new_n505), .A4(new_n850), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n672), .B1(new_n875), .B2(new_n793), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n660), .B1(new_n876), .B2(new_n811), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n361), .B1(new_n877), .B2(new_n815), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n873), .B1(new_n878), .B2(KEYINPUT57), .ZN(new_n879));
  INV_X1    g678(.A(new_n845), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n625), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n868), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n879), .ZN(new_n885));
  INV_X1    g684(.A(new_n881), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT120), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n870), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n846), .A2(new_n239), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n855), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n880), .B1(new_n890), .B2(new_n857), .ZN(new_n891));
  AOI211_X1 g690(.A(KEYINPUT59), .B(new_n868), .C1(new_n891), .C2(new_n626), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n869), .B1(new_n888), .B2(new_n892), .ZN(G1345gat));
  NOR2_X1   g692(.A1(new_n660), .A2(new_n212), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n212), .B1(new_n842), .B2(new_n660), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(G1346gat));
  AOI21_X1  g699(.A(G162gat), .B1(new_n867), .B2(new_n672), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n599), .A2(new_n213), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n891), .B2(new_n902), .ZN(G1347gat));
  AOI21_X1  g702(.A(new_n283), .B1(new_n814), .B2(new_n815), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n733), .A2(new_n734), .A3(new_n437), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT122), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(G169gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n505), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(KEYINPUT123), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(KEYINPUT123), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n650), .A2(new_n437), .A3(new_n239), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n904), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n505), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n916), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT124), .B1(new_n916), .B2(G169gat), .ZN(new_n918));
  OAI22_X1  g717(.A1(new_n911), .A2(new_n912), .B1(new_n917), .B2(new_n918), .ZN(G1348gat));
  INV_X1    g718(.A(G176gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n908), .A2(new_n920), .A3(new_n626), .ZN(new_n921));
  OAI21_X1  g720(.A(G176gat), .B1(new_n914), .B2(new_n625), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1349gat));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n309), .A3(new_n542), .ZN(new_n924));
  OAI21_X1  g723(.A(G183gat), .B1(new_n914), .B2(new_n660), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g726(.A1(new_n908), .A2(new_n310), .A3(new_n672), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n915), .A2(new_n672), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(G190gat), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT61), .B(new_n310), .C1(new_n915), .C2(new_n672), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(G1351gat));
  INV_X1    g732(.A(G197gat), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n425), .A2(new_n283), .A3(new_n437), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n879), .A2(new_n505), .A3(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n938), .B1(new_n937), .B2(new_n936), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n838), .A2(new_n437), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n904), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n934), .A3(new_n505), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n939), .A2(new_n943), .ZN(G1352gat));
  NOR3_X1   g743(.A1(new_n941), .A2(G204gat), .A3(new_n625), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT62), .ZN(new_n946));
  INV_X1    g745(.A(G204gat), .ZN(new_n947));
  INV_X1    g746(.A(new_n935), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n885), .A2(new_n625), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n947), .B2(new_n949), .ZN(G1353gat));
  NAND3_X1  g749(.A1(new_n942), .A2(new_n205), .A3(new_n542), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT57), .B1(new_n854), .B2(new_n239), .ZN(new_n954));
  INV_X1    g753(.A(new_n856), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n814), .B2(new_n815), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n542), .B(new_n935), .C1(new_n954), .C2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n879), .A2(KEYINPUT126), .A3(new_n542), .A4(new_n935), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n205), .B1(KEYINPUT127), .B2(new_n952), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n953), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n953), .ZN(new_n964));
  INV_X1    g763(.A(new_n962), .ZN(new_n965));
  AOI211_X1 g764(.A(new_n964), .B(new_n965), .C1(new_n959), .C2(new_n960), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n951), .B1(new_n963), .B2(new_n966), .ZN(G1354gat));
  NAND3_X1  g766(.A1(new_n942), .A2(new_n206), .A3(new_n672), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n885), .A2(new_n599), .A3(new_n948), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(new_n206), .ZN(G1355gat));
endmodule


