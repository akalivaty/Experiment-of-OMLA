//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  AND2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n206), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  AOI211_X1 g0015(.A(new_n213), .B(new_n215), .C1(G50), .C2(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n201), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n202), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n209), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NAND2_X1  g0027(.A1(new_n203), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n224), .A2(new_n227), .A3(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G226), .B(G232), .Z(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n219), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT67), .B(G264), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n237), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT84), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  OAI211_X1 g0057(.A(G1), .B(G13), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n252), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G226), .ZN(new_n261));
  INV_X1    g0061(.A(new_n258), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT68), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n263), .B2(new_n265), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  MUX2_X1   g0069(.A(G222), .B(G223), .S(G1698), .Z(new_n270));
  OAI21_X1  g0070(.A(new_n262), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n264), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT68), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G77), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n255), .B(new_n261), .C1(new_n271), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G190), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT76), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(KEYINPUT9), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n229), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT69), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n229), .A2(new_n256), .A3(KEYINPUT70), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(G20), .B2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G150), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n285), .A2(new_n286), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI221_X1 g0095(.A(KEYINPUT71), .B1(new_n291), .B2(new_n292), .C1(new_n285), .C2(new_n286), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n295), .B(new_n296), .C1(new_n229), .C2(new_n205), .ZN(new_n297));
  NAND3_X1  g0097(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n230), .ZN(new_n299));
  INV_X1    g0099(.A(G50), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n297), .A2(new_n299), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n281), .A2(KEYINPUT9), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n301), .A2(new_n230), .A3(new_n298), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT72), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n229), .B2(G1), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n251), .A2(KEYINPUT72), .A3(G20), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G50), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n303), .A2(new_n304), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n304), .B1(new_n303), .B2(new_n311), .ZN(new_n313));
  OAI211_X1 g0113(.A(KEYINPUT77), .B(new_n282), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n278), .A2(G200), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(new_n282), .C1(new_n312), .C2(new_n313), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n314), .A3(new_n315), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n303), .A2(new_n311), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n278), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n322), .B(new_n324), .C1(G179), .C2(new_n278), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n320), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G1698), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n276), .A2(G232), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n276), .A2(G238), .A3(G1698), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n269), .A2(G107), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT73), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT73), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n328), .A2(new_n329), .A3(new_n330), .A4(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n262), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n254), .B1(new_n260), .B2(G244), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n323), .ZN(new_n338));
  INV_X1    g0138(.A(new_n299), .ZN(new_n339));
  XOR2_X1   g0139(.A(KEYINPUT8), .B(G58), .Z(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT74), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT74), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n286), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n290), .A3(new_n343), .ZN(new_n344));
  XOR2_X1   g0144(.A(KEYINPUT15), .B(G87), .Z(new_n345));
  INV_X1    g0145(.A(new_n283), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n345), .A2(new_n346), .B1(G20), .B2(G77), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n339), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n301), .A2(G77), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n310), .A2(G77), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G179), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n335), .A2(new_n353), .A3(new_n336), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n338), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n352), .A2(KEYINPUT75), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT75), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n350), .A2(new_n358), .A3(new_n351), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n357), .B(new_n359), .C1(new_n337), .C2(new_n279), .ZN(new_n360));
  INV_X1    g0160(.A(G200), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n335), .B2(new_n336), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n326), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n290), .A2(G50), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n367), .B1(new_n229), .B2(G68), .C1(new_n285), .C2(new_n206), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n299), .ZN(new_n369));
  XOR2_X1   g0169(.A(new_n369), .B(KEYINPUT11), .Z(new_n370));
  NAND2_X1  g0170(.A1(new_n302), .A2(new_n202), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(KEYINPUT12), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(KEYINPUT12), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n372), .A2(new_n373), .B1(G68), .B2(new_n310), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT13), .ZN(new_n377));
  NOR2_X1   g0177(.A1(G226), .A2(G1698), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n217), .B2(G1698), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n267), .B2(new_n268), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G97), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n258), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n255), .B1(new_n259), .B2(new_n221), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n377), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n383), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n276), .A2(new_n379), .B1(G33), .B2(G97), .ZN(new_n386));
  OAI211_X1 g0186(.A(KEYINPUT13), .B(new_n385), .C1(new_n386), .C2(new_n258), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT14), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n384), .A2(new_n387), .A3(new_n388), .A4(G169), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n377), .A2(KEYINPUT78), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n382), .B2(new_n383), .ZN(new_n391));
  INV_X1    g0191(.A(new_n390), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n385), .B(new_n392), .C1(new_n386), .C2(new_n258), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n393), .A3(G179), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n384), .A2(new_n387), .A3(G169), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(KEYINPUT79), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT79), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(new_n395), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n376), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n384), .A2(new_n387), .A3(G200), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n391), .A2(new_n393), .A3(G190), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n376), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g0208(.A(G58), .B(G68), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n290), .A2(G159), .B1(new_n409), .B2(G20), .ZN(new_n410));
  AOI21_X1  g0210(.A(G20), .B1(new_n263), .B2(new_n265), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT7), .ZN(new_n412));
  OAI21_X1  g0212(.A(G68), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT3), .B(G33), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n414), .A2(KEYINPUT7), .A3(G20), .ZN(new_n415));
  OAI211_X1 g0215(.A(KEYINPUT16), .B(new_n410), .C1(new_n413), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n299), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n410), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT81), .B1(new_n264), .B2(G33), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT81), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(new_n256), .A3(KEYINPUT3), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n422), .A3(new_n265), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n267), .A2(new_n268), .A3(G20), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(KEYINPUT7), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n419), .B1(new_n426), .B2(G68), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n418), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n327), .A2(G226), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n414), .B(new_n430), .C1(G223), .C2(G1698), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G87), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n258), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n259), .A2(new_n217), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n433), .A2(new_n254), .A3(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n279), .A2(KEYINPUT83), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n279), .A2(KEYINPUT83), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT82), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n340), .B1(new_n305), .B2(new_n309), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n286), .A2(new_n301), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n441), .A3(new_n443), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n435), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G200), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n429), .A2(new_n440), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n446), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n444), .ZN(new_n454));
  INV_X1    g0254(.A(new_n428), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n274), .A2(new_n229), .A3(new_n275), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n412), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n202), .B1(new_n457), .B2(new_n424), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n455), .B1(new_n458), .B2(new_n419), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n454), .B1(new_n459), .B2(new_n418), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n460), .A2(KEYINPUT17), .A3(new_n440), .A4(new_n449), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n452), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n429), .A2(new_n447), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n435), .A2(G179), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(new_n435), .B2(new_n323), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT18), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT18), .ZN(new_n467));
  NOR4_X1   g0267(.A1(new_n433), .A2(new_n353), .A3(new_n434), .A4(new_n254), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n448), .B2(G169), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n460), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n408), .A2(new_n462), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n250), .B1(new_n366), .B2(new_n473), .ZN(new_n474));
  NOR4_X1   g0274(.A1(new_n326), .A2(new_n472), .A3(KEYINPUT84), .A4(new_n365), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT24), .ZN(new_n478));
  AOI21_X1  g0278(.A(G20), .B1(new_n274), .B2(new_n275), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT22), .B1(new_n479), .B2(G87), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n229), .A2(G107), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n481), .B(KEYINPUT23), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  INV_X1    g0283(.A(G87), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n414), .A2(new_n485), .B1(G33), .B2(G116), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n482), .B1(new_n486), .B2(G20), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n478), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n229), .B(G87), .C1(new_n267), .C2(new_n268), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n483), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n486), .A2(G20), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT24), .A4(new_n482), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n299), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n305), .B1(new_n251), .B2(G33), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G107), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n301), .A2(G107), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT89), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(KEYINPUT25), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(KEYINPUT25), .ZN(new_n499));
  MUX2_X1   g0299(.A(new_n496), .B(new_n498), .S(new_n499), .Z(new_n500));
  NAND3_X1  g0300(.A1(new_n493), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G45), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(G1), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n257), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G41), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n253), .ZN(new_n508));
  OR2_X1    g0308(.A1(G250), .A2(G1698), .ZN(new_n509));
  INV_X1    g0309(.A(G257), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n263), .A2(new_n509), .A3(new_n265), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n258), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n507), .A2(G264), .A3(new_n258), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT90), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n507), .A2(KEYINPUT90), .A3(G264), .A4(new_n258), .ZN(new_n518));
  AOI211_X1 g0318(.A(new_n508), .B(new_n514), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT91), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n520), .A3(G179), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(new_n518), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n507), .A2(new_n253), .ZN(new_n523));
  INV_X1    g0323(.A(new_n514), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT91), .B1(new_n525), .B2(new_n353), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n523), .A3(new_n515), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G169), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n521), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n501), .A2(new_n529), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n519), .A2(G200), .B1(G190), .B2(new_n527), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n531), .A2(new_n493), .A3(new_n495), .A4(new_n500), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n507), .A2(new_n258), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n219), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n274), .A2(G303), .A3(new_n275), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n212), .A2(G1698), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n414), .B(new_n537), .C1(G257), .C2(G1698), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n535), .B1(new_n539), .B2(new_n262), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n323), .B1(new_n540), .B2(new_n523), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n251), .A2(G33), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n339), .A2(G116), .A3(new_n301), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n302), .A2(new_n218), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n298), .A2(new_n230), .B1(G20), .B2(new_n218), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G283), .ZN(new_n546));
  INV_X1    g0346(.A(G97), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n546), .B(new_n229), .C1(G33), .C2(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n545), .A2(KEYINPUT20), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT20), .B1(new_n545), .B2(new_n548), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n543), .B(new_n544), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n541), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT21), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n540), .A2(new_n523), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n353), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n551), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n541), .A2(KEYINPUT21), .A3(new_n551), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT88), .ZN(new_n560));
  INV_X1    g0360(.A(new_n551), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n555), .B2(new_n438), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n258), .B1(new_n536), .B2(new_n538), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n563), .A2(new_n508), .A3(new_n535), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(new_n361), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n560), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  OR3_X1    g0366(.A1(new_n562), .A2(new_n560), .A3(new_n565), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n559), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G250), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n210), .A2(G1698), .ZN(new_n570));
  OAI211_X1 g0370(.A(KEYINPUT4), .B(new_n570), .C1(new_n267), .C2(new_n268), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n414), .A2(new_n570), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n572), .A2(new_n573), .B1(G33), .B2(G283), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n569), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n262), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n523), .B1(new_n510), .B2(new_n534), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n323), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  AOI211_X1 g0379(.A(new_n353), .B(new_n577), .C1(new_n575), .C2(new_n262), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n211), .B1(new_n457), .B2(new_n424), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT6), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n547), .A2(new_n211), .ZN(new_n584));
  NOR2_X1   g0384(.A1(G97), .A2(G107), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n211), .A2(KEYINPUT6), .A3(G97), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n588), .A2(new_n229), .B1(new_n206), .B2(new_n291), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n299), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n301), .A2(G97), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n494), .B2(G97), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT85), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT85), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n590), .A2(new_n595), .A3(new_n592), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n581), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n221), .A2(new_n327), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n210), .A2(G1698), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n414), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G33), .A2(G116), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n262), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n251), .A2(G45), .ZN(new_n604));
  AND2_X1   g0404(.A1(G33), .A2(G41), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n604), .B(G250), .C1(new_n605), .C2(new_n230), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT86), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n604), .B2(new_n253), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n503), .A2(KEYINPUT86), .A3(G274), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n603), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G200), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n258), .B1(new_n600), .B2(new_n601), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(new_n610), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G190), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT19), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n229), .B1(new_n381), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n585), .A2(new_n484), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT87), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n618), .B1(new_n283), .B2(new_n547), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n414), .A2(new_n229), .A3(G68), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n619), .A2(new_n620), .A3(KEYINPUT87), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n623), .A2(new_n624), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n345), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n627), .A2(new_n299), .B1(new_n302), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n494), .A2(G87), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n614), .A2(G179), .A3(new_n610), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n494), .A2(new_n345), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(new_n629), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n612), .A2(new_n323), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n617), .A2(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n577), .B1(new_n575), .B2(new_n262), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n639), .A2(G190), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n361), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n593), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n597), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n477), .A2(new_n533), .A3(new_n568), .A4(new_n643), .ZN(G372));
  OAI21_X1  g0444(.A(new_n593), .B1(new_n579), .B2(new_n580), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n627), .A2(new_n299), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n628), .A2(new_n302), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n634), .ZN(new_n648));
  INV_X1    g0448(.A(new_n633), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT92), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n610), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n606), .A2(new_n608), .A3(new_n609), .A4(KEYINPUT92), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n614), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G169), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n616), .B1(new_n654), .B2(new_n361), .ZN(new_n656));
  OAI22_X1  g0456(.A1(new_n650), .A2(new_n655), .B1(new_n656), .B2(new_n631), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n645), .A2(new_n657), .A3(KEYINPUT26), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n579), .A2(new_n580), .ZN(new_n659));
  INV_X1    g0459(.A(new_n596), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n595), .B1(new_n590), .B2(new_n592), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n637), .B(new_n659), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n658), .B1(KEYINPUT26), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT21), .B1(new_n541), .B2(new_n551), .ZN(new_n664));
  NOR4_X1   g0464(.A1(new_n564), .A2(new_n561), .A3(new_n553), .A4(new_n323), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n530), .A2(new_n666), .A3(new_n557), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n652), .A2(new_n653), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n603), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n670), .A2(G200), .B1(G190), .B2(new_n615), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n323), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n632), .A2(new_n671), .B1(new_n635), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(new_n532), .ZN(new_n674));
  INV_X1    g0474(.A(new_n642), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n667), .A2(new_n668), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n635), .A2(new_n672), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n663), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n477), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n407), .A2(new_n355), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n462), .B1(new_n680), .B2(new_n403), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n681), .A2(new_n471), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n320), .A2(new_n321), .ZN(new_n683));
  OAI211_X1 g0483(.A(KEYINPUT93), .B(new_n325), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT93), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n683), .B1(new_n471), .B2(new_n681), .ZN(new_n686));
  INV_X1    g0486(.A(new_n325), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n679), .A2(new_n689), .ZN(G369));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n229), .A2(G13), .ZN(new_n692));
  OR3_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .A3(G1), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT27), .B1(new_n692), .B2(G1), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n568), .B1(new_n561), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n559), .A2(new_n551), .A3(new_n697), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n691), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n530), .A2(new_n698), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n501), .A2(new_n697), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n533), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n697), .B1(new_n666), .B2(new_n557), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n533), .A2(new_n705), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n501), .A2(new_n529), .A3(new_n698), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(G399));
  NOR2_X1   g0512(.A1(new_n620), .A2(G116), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n225), .A2(new_n257), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n714), .A3(G1), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n228), .B2(new_n714), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT94), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n643), .A2(new_n568), .A3(new_n533), .A4(new_n698), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n615), .A2(new_n524), .A3(new_n522), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n556), .A2(new_n639), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(KEYINPUT96), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(KEYINPUT96), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n556), .A2(new_n639), .A3(new_n724), .A4(new_n720), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n555), .A2(new_n525), .A3(new_n670), .ZN(new_n726));
  OR3_X1    g0526(.A1(new_n726), .A2(G179), .A3(new_n639), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n723), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n697), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n719), .B(new_n731), .C1(new_n729), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT26), .B1(new_n645), .B2(new_n657), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n677), .B(new_n737), .C1(new_n662), .C2(KEYINPUT26), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT97), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT26), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n597), .A2(new_n740), .A3(new_n637), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT97), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(new_n677), .A4(new_n737), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n743), .A3(new_n676), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n736), .B1(new_n744), .B2(new_n698), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n678), .A2(new_n698), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(KEYINPUT29), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n735), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n718), .B1(new_n748), .B2(G1), .ZN(G364));
  NOR3_X1   g0549(.A1(new_n229), .A2(new_n353), .A3(new_n361), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n439), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n276), .B1(new_n751), .B2(new_n300), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n229), .A2(new_n353), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n361), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n438), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n361), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G20), .A3(G190), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n756), .A2(new_n201), .B1(new_n484), .B2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n279), .A2(G179), .A3(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n229), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n752), .B(new_n759), .C1(G97), .C2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n753), .A2(new_n279), .A3(new_n361), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT101), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(KEYINPUT101), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G77), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n229), .A2(G190), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n353), .A3(new_n361), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT32), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n770), .A2(new_n757), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT102), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n750), .A2(new_n279), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n777), .A2(G107), .B1(G68), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n763), .A2(new_n769), .A3(new_n774), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n764), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n751), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n276), .B1(new_n784), .B2(G326), .ZN(new_n785));
  INV_X1    g0585(.A(G329), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n786), .B2(new_n771), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n783), .B(new_n787), .C1(G322), .C2(new_n755), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT33), .B(G317), .ZN(new_n789));
  INV_X1    g0589(.A(new_n758), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n779), .A2(new_n789), .B1(G303), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n788), .B(new_n791), .C1(new_n792), .C2(new_n776), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n761), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n781), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n230), .B1(G20), .B2(new_n323), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n797), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT100), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n276), .A2(G355), .A3(new_n225), .ZN(new_n804));
  INV_X1    g0604(.A(new_n414), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n225), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT99), .Z(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n502), .B2(new_n248), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n228), .A2(G45), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n804), .B1(G116), .B2(new_n225), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n796), .A2(new_n797), .B1(new_n803), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n699), .A2(new_n700), .A3(new_n800), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n692), .B(KEYINPUT98), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G45), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G1), .ZN(new_n815));
  INV_X1    g0615(.A(new_n714), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n811), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AND3_X1   g0619(.A1(new_n699), .A2(new_n691), .A3(new_n700), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n701), .ZN(new_n821));
  INV_X1    g0621(.A(new_n817), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  NAND2_X1  g0624(.A1(new_n352), .A2(new_n697), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n360), .B2(new_n362), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n355), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n356), .A2(new_n698), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n746), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n678), .A2(new_n364), .A3(new_n698), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(new_n735), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n822), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n829), .A2(new_n798), .ZN(new_n835));
  INV_X1    g0635(.A(new_n771), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n755), .A2(G294), .B1(G311), .B2(new_n836), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n767), .A2(new_n218), .B1(new_n792), .B2(new_n778), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n837), .B1(new_n547), .B2(new_n761), .C1(new_n838), .C2(KEYINPUT103), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(KEYINPUT103), .B2(new_n838), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n777), .A2(G87), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n784), .A2(G303), .B1(G107), .B2(new_n790), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n840), .A2(new_n269), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G143), .A2(new_n755), .B1(new_n779), .B2(G150), .ZN(new_n844));
  INV_X1    g0644(.A(G137), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n844), .B1(new_n845), .B2(new_n751), .C1(new_n767), .C2(new_n772), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT34), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n790), .A2(G50), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n777), .A2(G68), .B1(G132), .B2(new_n836), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n847), .A2(new_n414), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n761), .A2(new_n201), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n843), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n797), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n797), .A2(new_n798), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n206), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n835), .A2(new_n817), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n834), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  OAI22_X1  g0658(.A1(new_n474), .A2(new_n475), .B1(new_n745), .B2(new_n747), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n689), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT108), .Z(new_n861));
  OAI211_X1 g0661(.A(new_n452), .B(new_n461), .C1(new_n466), .C2(new_n470), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n411), .A2(new_n412), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT7), .B1(new_n414), .B2(G20), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(G68), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n428), .B1(new_n865), .B2(new_n410), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n417), .A2(new_n866), .B1(new_n444), .B2(new_n453), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT105), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n695), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n447), .B(KEYINPUT105), .C1(new_n417), .C2(new_n866), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n862), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n869), .A2(new_n465), .A3(new_n871), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n450), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT106), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(new_n450), .A3(KEYINPUT106), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n874), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT107), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n460), .B2(new_n695), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n423), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n412), .B2(new_n456), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n410), .B1(new_n884), .B2(new_n202), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n417), .B1(new_n885), .B2(new_n455), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT107), .B(new_n870), .C1(new_n886), .C2(new_n454), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n463), .A2(new_n465), .ZN(new_n889));
  AND4_X1   g0689(.A1(new_n874), .A2(new_n888), .A3(new_n450), .A4(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(KEYINPUT38), .B(new_n873), .C1(new_n880), .C2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n888), .A2(new_n450), .A3(new_n889), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n888), .A2(new_n874), .A3(new_n450), .A4(new_n889), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n888), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n862), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n891), .B1(new_n898), .B2(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n729), .A2(new_n732), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n719), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n376), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT79), .B1(new_n396), .B2(new_n398), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n401), .A2(new_n395), .A3(new_n400), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(new_n697), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n406), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n403), .A2(new_n697), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n829), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n902), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n873), .B1(new_n880), .B2(new_n890), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n891), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n912), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT109), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT109), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n921), .B(KEYINPUT40), .C1(new_n917), .C2(new_n912), .ZN(new_n922));
  OAI211_X1 g0722(.A(G330), .B(new_n913), .C1(new_n920), .C2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(G330), .B(new_n902), .C1(new_n474), .C2(new_n475), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n477), .A2(new_n902), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n912), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n902), .A2(new_n910), .A3(new_n911), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n891), .B2(new_n916), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n921), .B1(new_n928), .B2(KEYINPUT40), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n918), .A2(KEYINPUT109), .A3(new_n919), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n923), .A2(new_n924), .B1(new_n925), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n861), .B(new_n932), .Z(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  INV_X1    g0734(.A(new_n891), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n895), .B2(new_n897), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n916), .A2(KEYINPUT39), .A3(new_n891), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n906), .A2(new_n697), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n471), .A2(new_n870), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n408), .A2(new_n907), .B1(new_n403), .B2(new_n697), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n831), .B2(new_n828), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n943), .B1(new_n917), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n933), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n933), .A2(new_n948), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n949), .B(new_n950), .C1(new_n251), .C2(new_n813), .ZN(new_n951));
  OAI21_X1  g0751(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n228), .A2(new_n952), .B1(G50), .B2(new_n202), .ZN(new_n953));
  INV_X1    g0753(.A(G13), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(G1), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT35), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n229), .B(new_n230), .C1(new_n588), .C2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n957), .B(G116), .C1(new_n956), .C2(new_n588), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT104), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT36), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n951), .A2(new_n955), .A3(new_n960), .ZN(G367));
  NOR2_X1   g0761(.A1(new_n645), .A2(new_n698), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n597), .A2(new_n642), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n593), .A2(new_n697), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n708), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n668), .B1(new_n965), .B2(new_n530), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT110), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n698), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n963), .A2(new_n533), .A3(new_n705), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT42), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n631), .A2(new_n697), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n673), .A2(new_n973), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n677), .A2(new_n973), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n970), .A2(new_n972), .B1(KEYINPUT43), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n977), .A2(new_n979), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n967), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT111), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n815), .ZN(new_n985));
  INV_X1    g0785(.A(new_n748), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n701), .A2(new_n707), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n710), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n709), .A2(new_n711), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n965), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT44), .Z(new_n992));
  NOR2_X1   g0792(.A1(new_n990), .A2(new_n965), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n986), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n714), .B(KEYINPUT41), .Z(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n985), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  OR3_X1    g0799(.A1(new_n980), .A2(new_n981), .A3(new_n967), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n982), .A2(new_n983), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n984), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n807), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n803), .B1(new_n225), .B2(new_n628), .C1(new_n1003), .C2(new_n241), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n976), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n822), .B1(new_n1005), .B2(new_n800), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n758), .A2(new_n218), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n414), .B1(new_n1007), .B2(KEYINPUT46), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n211), .B2(new_n761), .C1(new_n767), .C2(new_n792), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1007), .A2(KEYINPUT46), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G294), .B2(new_n779), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n775), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G317), .A2(new_n836), .B1(new_n1012), .B2(G97), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(new_n782), .C2(new_n751), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1009), .B(new_n1014), .C1(G303), .C2(new_n755), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n779), .A2(G159), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n276), .B1(new_n756), .B2(new_n292), .C1(new_n767), .C2(new_n300), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n771), .A2(new_n845), .B1(new_n775), .B2(new_n206), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n762), .A2(G68), .ZN(new_n1019));
  INV_X1    g0819(.A(G143), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1019), .B1(new_n201), .B2(new_n758), .C1(new_n751), .C2(new_n1020), .ZN(new_n1021));
  NOR3_X1   g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1015), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT47), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n797), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1004), .B(new_n1006), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1002), .A2(new_n1026), .ZN(G387));
  OAI21_X1  g0827(.A(new_n805), .B1(new_n775), .B2(new_n218), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G317), .A2(new_n755), .B1(new_n779), .B2(G311), .ZN(new_n1029));
  INV_X1    g0829(.A(G322), .ZN(new_n1030));
  INV_X1    g0830(.A(G303), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1029), .B1(new_n1030), .B2(new_n751), .C1(new_n767), .C2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT48), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n792), .B2(new_n761), .C1(new_n794), .C2(new_n758), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1028), .B(new_n1036), .C1(G326), .C2(new_n836), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n414), .B1(new_n286), .B2(new_n778), .C1(new_n776), .C2(new_n547), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n784), .A2(G159), .B1(new_n345), .B2(new_n762), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n202), .B2(new_n764), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G77), .B2(new_n790), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n300), .B2(new_n756), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1038), .B(new_n1042), .C1(G150), .C2(new_n836), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n797), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n704), .A2(new_n800), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n276), .A2(new_n225), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1046), .A2(new_n713), .B1(G107), .B2(new_n225), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT112), .Z(new_n1048));
  NAND3_X1  g0848(.A1(new_n341), .A2(new_n300), .A3(new_n343), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT50), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1049), .A2(KEYINPUT50), .B1(G68), .B2(G77), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1050), .A2(new_n1051), .A3(new_n502), .A4(new_n713), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1003), .B1(new_n237), .B2(G45), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1048), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n817), .B1(new_n1054), .B2(new_n802), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT113), .Z(new_n1056));
  NAND3_X1  g0856(.A1(new_n1044), .A2(new_n1045), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n986), .A2(new_n988), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n816), .B1(new_n989), .B2(new_n748), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1057), .B1(new_n985), .B2(new_n988), .C1(new_n1058), .C2(new_n1059), .ZN(G393));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n995), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n708), .A2(KEYINPUT115), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n995), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n708), .A2(KEYINPUT115), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n816), .B(new_n1061), .C1(new_n1065), .C2(new_n1058), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n965), .A2(new_n800), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n803), .B1(new_n547), .B2(new_n225), .C1(new_n1003), .C2(new_n245), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n784), .A2(G150), .B1(G159), .B2(new_n755), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT51), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G50), .B2(new_n779), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n836), .A2(G143), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n777), .A2(G87), .B1(G77), .B2(new_n762), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n341), .A2(new_n343), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n414), .B1(new_n767), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G68), .B2(new_n790), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n784), .A2(G317), .B1(G311), .B2(new_n755), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n764), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1080), .B1(G294), .B2(new_n1081), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n218), .B2(new_n761), .C1(new_n1031), .C2(new_n778), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n276), .B1(new_n777), .B2(G107), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n792), .B2(new_n758), .C1(new_n1030), .C2(new_n771), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT116), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1078), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n822), .B(new_n1069), .C1(new_n797), .C2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n1065), .B2(new_n815), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1066), .A2(new_n1089), .ZN(G390));
  INV_X1    g0890(.A(KEYINPUT119), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n831), .A2(new_n828), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n910), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n941), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(KEYINPUT117), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT117), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n945), .B2(new_n941), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n939), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n744), .A2(new_n364), .A3(new_n698), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1099), .A2(new_n828), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1094), .B(new_n899), .C1(new_n1100), .C2(new_n944), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n902), .A2(G330), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n829), .B1(new_n908), .B2(new_n909), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT118), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT118), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1103), .A2(new_n1107), .A3(new_n1104), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1091), .B1(new_n1102), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1111));
  AND4_X1   g0911(.A1(new_n1107), .A2(new_n1104), .A3(G330), .A4(new_n902), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(KEYINPUT119), .B(new_n1113), .C1(new_n1098), .C2(new_n1101), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n734), .A2(new_n829), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n910), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1098), .A2(new_n1101), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1110), .A2(new_n1114), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n815), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n940), .A2(new_n799), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n784), .A2(G128), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT54), .B(G143), .Z(new_n1123));
  AOI22_X1  g0923(.A1(new_n768), .A2(new_n1123), .B1(G137), .B2(new_n779), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1124), .A2(KEYINPUT120), .B1(new_n772), .B2(new_n761), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1122), .B(new_n1125), .C1(G132), .C2(new_n755), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(KEYINPUT120), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n758), .A2(new_n292), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n771), .A2(new_n1130), .B1(new_n775), .B2(new_n300), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1131), .A2(new_n269), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .A4(new_n1132), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n269), .B1(new_n756), .B2(new_n218), .C1(new_n767), .C2(new_n547), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G294), .B2(new_n836), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n779), .A2(G107), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n777), .A2(G68), .B1(G77), .B2(new_n762), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n784), .A2(G283), .B1(G87), .B2(new_n790), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1025), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n854), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1141), .A2(new_n340), .ZN(new_n1142));
  OR4_X1    g0942(.A1(new_n822), .A2(new_n1121), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n924), .A2(new_n859), .A3(new_n689), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1115), .A2(new_n910), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1092), .B1(new_n1109), .B2(new_n1145), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1103), .A2(new_n911), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1116), .B(new_n1100), .C1(new_n910), .C2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1144), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1119), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1102), .A2(new_n1109), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(KEYINPUT119), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1102), .A2(new_n1091), .A3(new_n1109), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1152), .A2(new_n1117), .A3(new_n1149), .A4(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n816), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1120), .B(new_n1143), .C1(new_n1150), .C2(new_n1155), .ZN(G378));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1144), .B1(new_n1119), .B2(new_n1149), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n322), .A2(new_n870), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n326), .B(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n923), .A2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1161), .B(new_n1162), .Z(new_n1165));
  NAND3_X1  g0965(.A1(new_n931), .A2(new_n1165), .A3(G330), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1164), .A2(new_n1166), .A3(new_n948), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n948), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1157), .B1(new_n1158), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1144), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1154), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n923), .A2(new_n1163), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1165), .B1(new_n931), .B2(G330), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n947), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1164), .A2(new_n1166), .A3(new_n948), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1172), .A2(new_n1177), .A3(KEYINPUT57), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1170), .A2(new_n816), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n985), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1163), .A2(new_n798), .ZN(new_n1181));
  INV_X1    g0981(.A(G124), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n257), .B1(new_n771), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n790), .A2(new_n1123), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n751), .B2(new_n1130), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n779), .A2(G132), .B1(new_n1081), .B2(G137), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n292), .B2(new_n761), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G128), .C2(new_n755), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT59), .ZN(new_n1189));
  AOI211_X1 g0989(.A(G33), .B(new_n1183), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n1189), .B2(new_n1188), .C1(new_n772), .C2(new_n775), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1191), .B1(G50), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n414), .B1(new_n1012), .B2(G58), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1019), .B(new_n1194), .C1(new_n751), .C2(new_n218), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n345), .A2(new_n1081), .B1(new_n836), .B2(G283), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G41), .B1(new_n790), .B2(G77), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n211), .C2(new_n756), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1195), .B(new_n1198), .C1(G97), .C2(new_n779), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT121), .Z(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT58), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n797), .B1(new_n1193), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n854), .A2(new_n300), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1181), .A2(new_n817), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(KEYINPUT122), .B1(new_n1180), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n815), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT122), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n1208), .A3(new_n1204), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1179), .A2(KEYINPUT123), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT123), .B1(new_n1179), .B2(new_n1210), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(G375));
  OAI22_X1  g1014(.A1(new_n910), .A2(new_n799), .B1(G68), .B2(new_n1141), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n768), .A2(G107), .B1(new_n345), .B2(new_n762), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n778), .A2(new_n218), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n771), .A2(new_n1031), .B1(new_n758), .B2(new_n547), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(new_n784), .C2(G294), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n755), .A2(G283), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n276), .B1(new_n777), .B2(G77), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1216), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n779), .A2(new_n1123), .B1(new_n762), .B2(G50), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n201), .B2(new_n775), .C1(new_n772), .C2(new_n758), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G137), .B2(new_n755), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n784), .A2(G132), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n805), .B1(new_n836), .B2(G128), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n764), .A2(new_n292), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1222), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n822), .B(new_n1215), .C1(new_n797), .C2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n1232), .B2(new_n815), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1146), .A2(new_n1144), .A3(new_n1148), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n997), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1235), .B2(new_n1149), .ZN(G381));
  INV_X1    g1036(.A(KEYINPUT123), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1172), .A2(new_n1177), .A3(KEYINPUT57), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT57), .B1(new_n1172), .B2(new_n1177), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1238), .A2(new_n1239), .A3(new_n714), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1180), .A2(KEYINPUT122), .A3(new_n1205), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1208), .B1(new_n1207), .B2(new_n1204), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1237), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(G378), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1179), .A2(KEYINPUT123), .A3(new_n1210), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(G381), .A2(G384), .ZN(new_n1248));
  INV_X1    g1048(.A(G390), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1002), .A2(new_n1026), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  OR3_X1    g1053(.A1(new_n1247), .A2(new_n1248), .A3(new_n1253), .ZN(G407));
  OAI21_X1  g1054(.A(G213), .B1(new_n1247), .B2(G343), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(G407), .A3(KEYINPUT124), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT124), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1247), .A2(new_n1248), .A3(new_n1253), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1258), .B1(new_n1259), .B2(new_n1255), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(G409));
  AOI21_X1  g1061(.A(new_n1245), .B1(new_n1179), .B2(new_n1210), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1172), .A2(new_n1177), .A3(new_n997), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n1207), .A3(new_n1204), .ZN(new_n1264));
  INV_X1    g1064(.A(G213), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n1264), .A2(G378), .B1(new_n1265), .B2(G343), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n857), .A2(KEYINPUT125), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT60), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1234), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1232), .A2(new_n1171), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1146), .A2(new_n1144), .A3(KEYINPUT60), .A4(new_n1148), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n816), .A4(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1267), .B1(new_n1272), .B2(new_n1233), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n857), .A2(KEYINPUT125), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1272), .A2(KEYINPUT125), .A3(new_n857), .A4(new_n1233), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1262), .A2(new_n1266), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT62), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n696), .A2(G213), .A3(G2897), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT126), .Z(new_n1285));
  XNOR2_X1  g1085(.A(new_n1277), .B(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1282), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  NOR4_X1   g1087(.A1(new_n1262), .A2(new_n1266), .A3(new_n1278), .A4(KEYINPUT62), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1281), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1249), .B1(new_n1002), .B2(new_n1026), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(G393), .B(new_n823), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1291), .A2(new_n1294), .A3(new_n1250), .A4(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1251), .B2(new_n1290), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT63), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1279), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1279), .A2(KEYINPUT63), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(new_n1282), .A3(new_n1299), .ZN(new_n1304));
  OAI22_X1  g1104(.A1(new_n1289), .A2(new_n1299), .B1(new_n1302), .B2(new_n1304), .ZN(G405));
  INV_X1    g1105(.A(new_n1262), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1247), .A2(new_n1306), .A3(new_n1277), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1277), .B1(new_n1247), .B2(new_n1306), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1307), .A2(new_n1308), .A3(new_n1299), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1299), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1211), .A2(new_n1212), .A3(G378), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1278), .B1(new_n1311), .B2(new_n1262), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1247), .A2(new_n1306), .A3(new_n1277), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1310), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1309), .A2(new_n1314), .ZN(G402));
endmodule


