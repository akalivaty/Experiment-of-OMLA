//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT0), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G57gat), .ZN(new_n205));
  INV_X1    g004(.A(G85gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G113gat), .ZN(new_n210));
  INV_X1    g009(.A(G113gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G120gat), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT1), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G127gat), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n214), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(G134gat), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G134gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n213), .A2(new_n214), .ZN(new_n219));
  AOI211_X1 g018(.A(KEYINPUT1), .B(G127gat), .C1(new_n210), .C2(new_n212), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G155gat), .ZN(new_n223));
  INV_X1    g022(.A(G162gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G141gat), .B(G148gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(KEYINPUT2), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G148gat), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n230), .A2(G141gat), .ZN(new_n231));
  XOR2_X1   g030(.A(KEYINPUT78), .B(G141gat), .Z(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(G148gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n225), .B1(new_n234), .B2(new_n226), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n229), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT3), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n222), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n236), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G225gat), .A2(G233gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n222), .A2(new_n236), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n236), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n242), .B(new_n243), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT5), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n217), .A2(new_n221), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n239), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n222), .A2(new_n236), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n243), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(KEYINPUT4), .ZN(new_n255));
  INV_X1    g054(.A(new_n247), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n255), .A2(new_n256), .B1(new_n241), .B2(new_n238), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n254), .B1(new_n257), .B2(new_n243), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n208), .B(new_n250), .C1(new_n258), .C2(new_n249), .ZN(new_n259));
  INV_X1    g058(.A(new_n254), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n249), .B1(new_n248), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT5), .B1(new_n257), .B2(new_n243), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n207), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT6), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n261), .A2(new_n262), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT6), .A3(new_n208), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT25), .ZN(new_n269));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT24), .ZN(new_n271));
  INV_X1    g070(.A(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n277));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n269), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n272), .A2(KEYINPUT65), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G183gat), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n271), .B1(new_n285), .B2(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n276), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n269), .B1(new_n290), .B2(KEYINPUT23), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n286), .A2(new_n291), .A3(new_n278), .A4(new_n277), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n281), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT26), .ZN(new_n294));
  INV_X1    g093(.A(new_n289), .ZN(new_n295));
  NOR3_X1   g094(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n278), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n284), .A3(KEYINPUT27), .ZN(new_n300));
  NOR2_X1   g099(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n273), .B1(new_n306), .B2(new_n301), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n307), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n299), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n299), .A2(new_n305), .A3(KEYINPUT66), .A4(new_n308), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n293), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n312), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n323));
  XNOR2_X1  g122(.A(G211gat), .B(G218gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G211gat), .A2(G218gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT22), .ZN(new_n327));
  INV_X1    g126(.A(G197gat), .ZN(new_n328));
  INV_X1    g127(.A(G204gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G197gat), .A2(G204gat), .ZN(new_n331));
  AOI221_X4 g130(.A(KEYINPUT74), .B1(new_n326), .B2(new_n327), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n333), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n323), .B(new_n325), .C1(new_n332), .C2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n335), .B1(new_n330), .B2(new_n331), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT75), .B1(new_n340), .B2(new_n324), .ZN(new_n341));
  AND2_X1   g140(.A1(G197gat), .A2(G204gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(G197gat), .A2(G204gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT74), .B1(new_n344), .B2(new_n335), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n334), .A2(new_n333), .A3(new_n336), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n324), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n338), .B(new_n339), .C1(new_n341), .C2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n325), .B1(new_n332), .B2(new_n337), .ZN(new_n350));
  INV_X1    g149(.A(new_n341), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n339), .B1(new_n352), .B2(new_n338), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n322), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n345), .A2(new_n346), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n341), .B1(new_n355), .B2(new_n325), .ZN(new_n356));
  AOI211_X1 g155(.A(KEYINPUT75), .B(new_n324), .C1(new_n345), .C2(new_n346), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT76), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(KEYINPUT77), .A3(new_n348), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n348), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n310), .A2(new_n315), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n320), .B2(new_n311), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n321), .A2(new_n360), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365));
  INV_X1    g164(.A(G64gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G92gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT30), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n363), .A2(new_n361), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n320), .A2(new_n315), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n311), .B2(new_n310), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n358), .A2(KEYINPUT77), .A3(new_n348), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT77), .B1(new_n358), .B2(new_n348), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n372), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(new_n369), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n369), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n370), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(KEYINPUT30), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n268), .A2(new_n384), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n319), .A2(new_n251), .A3(new_n293), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n251), .B1(new_n319), .B2(new_n293), .ZN(new_n387));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT34), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(KEYINPUT70), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n320), .A2(new_n222), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n319), .A2(new_n251), .A3(new_n293), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n393), .A2(new_n391), .A3(new_n388), .A4(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT70), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n388), .A3(new_n394), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT34), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n392), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT67), .B1(new_n401), .B2(KEYINPUT33), .ZN(new_n402));
  XNOR2_X1  g201(.A(G15gat), .B(G43gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(G71gat), .ZN(new_n404));
  INV_X1    g203(.A(G99gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n389), .B1(new_n386), .B2(new_n387), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(KEYINPUT32), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT67), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n402), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n406), .B2(KEYINPUT68), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n414), .B1(KEYINPUT68), .B2(new_n406), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n408), .A2(KEYINPUT32), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT69), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n408), .A2(KEYINPUT69), .A3(KEYINPUT32), .A4(new_n415), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n400), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT71), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n392), .A2(new_n397), .A3(new_n399), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n402), .A2(new_n409), .A3(new_n412), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n418), .A4(new_n419), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT71), .B(new_n400), .C1(new_n413), .C2(new_n420), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n241), .A2(new_n313), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n358), .A3(new_n348), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n325), .B1(new_n335), .B2(new_n344), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n340), .A2(new_n324), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT29), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n236), .B1(new_n432), .B2(KEYINPUT3), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n435), .B(KEYINPUT79), .Z(new_n436));
  AND2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n428), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n354), .B2(new_n359), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n352), .A2(new_n338), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT3), .B1(new_n440), .B2(new_n313), .ZN(new_n441));
  OAI211_X1 g240(.A(G228gat), .B(G233gat), .C1(new_n441), .C2(new_n239), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT80), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n428), .B1(new_n375), .B2(new_n376), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT80), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n440), .A2(new_n313), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n240), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n435), .B1(new_n447), .B2(new_n236), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n437), .B1(new_n443), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G22gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(G78gat), .B(G106gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT31), .ZN(new_n453));
  INV_X1    g252(.A(G50gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n437), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n439), .A2(new_n442), .A3(KEYINPUT80), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n445), .B1(new_n444), .B2(new_n448), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n455), .A2(KEYINPUT81), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(G22gat), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n450), .B2(new_n451), .ZN(new_n464));
  AOI211_X1 g263(.A(G22gat), .B(new_n437), .C1(new_n443), .C2(new_n449), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n456), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT82), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n460), .A2(G22gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n451), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n461), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT82), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n456), .A4(new_n463), .ZN(new_n472));
  AOI221_X4 g271(.A(new_n385), .B1(new_n426), .B2(new_n427), .C1(new_n467), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT35), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n202), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT35), .B1(new_n467), .B2(new_n472), .ZN(new_n476));
  INV_X1    g275(.A(new_n385), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT72), .ZN(new_n478));
  OR4_X1    g277(.A1(new_n478), .A2(new_n413), .A3(new_n420), .A4(new_n400), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n421), .A2(new_n478), .A3(new_n425), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n479), .A2(KEYINPUT87), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT87), .B1(new_n479), .B2(new_n480), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n476), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n472), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n426), .A2(new_n427), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n477), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(KEYINPUT88), .A3(KEYINPUT35), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n475), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n378), .A2(KEYINPUT37), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n369), .B1(new_n378), .B2(KEYINPUT37), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT38), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(new_n491), .B(KEYINPUT86), .Z(new_n492));
  NAND2_X1  g291(.A1(new_n374), .A2(new_n377), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n493), .A2(KEYINPUT84), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(KEYINPUT84), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n363), .A2(new_n361), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n496), .A2(KEYINPUT85), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(KEYINPUT85), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n494), .A2(new_n495), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT38), .B1(new_n499), .B2(KEYINPUT37), .ZN(new_n500));
  INV_X1    g299(.A(new_n490), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n268), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n492), .A2(new_n502), .A3(new_n382), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n257), .A2(new_n243), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n252), .A2(new_n243), .A3(new_n253), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(KEYINPUT39), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n506), .B(new_n207), .C1(KEYINPUT39), .C2(new_n504), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n507), .A2(new_n508), .B1(new_n208), .B2(new_n266), .ZN(new_n509));
  INV_X1    g308(.A(new_n384), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n509), .B(new_n510), .C1(new_n508), .C2(new_n507), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n503), .A2(new_n484), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n479), .A2(new_n480), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT73), .B1(new_n513), .B2(KEYINPUT36), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n485), .A2(KEYINPUT36), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT73), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n479), .A2(new_n516), .A3(new_n517), .A4(new_n480), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT83), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n484), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n467), .A2(KEYINPUT83), .A3(new_n472), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n512), .B(new_n519), .C1(new_n477), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n488), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G43gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(G50gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n454), .A2(G43gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT92), .ZN(new_n529));
  AOI22_X1  g328(.A1(KEYINPUT91), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT92), .B1(new_n454), .B2(G43gat), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n530), .B(new_n531), .C1(KEYINPUT91), .C2(new_n527), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(KEYINPUT90), .B(G29gat), .Z(new_n535));
  INV_X1    g334(.A(G36gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OR3_X1    g337(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT93), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  OR3_X1    g342(.A1(new_n528), .A2(new_n527), .A3(new_n533), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n538), .A2(new_n541), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n539), .B1(new_n537), .B2(new_n542), .ZN(new_n546));
  OAI22_X1  g345(.A1(new_n534), .A2(new_n545), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT17), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(KEYINPUT8), .A2(new_n549), .B1(new_n206), .B2(new_n368), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT101), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n206), .A2(new_n368), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G99gat), .B(G106gat), .Z(new_n556));
  OR2_X1    g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n548), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n559), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n547), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT41), .ZN(new_n563));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT99), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n560), .B(new_n562), .C1(new_n563), .C2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G190gat), .B(G218gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT102), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n563), .ZN(new_n572));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT103), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n570), .B2(KEYINPUT104), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n577), .B(new_n569), .C1(KEYINPUT104), .C2(new_n570), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G15gat), .B(G22gat), .Z(new_n580));
  INV_X1    g379(.A(KEYINPUT16), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(G1gat), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G8gat), .ZN(new_n584));
  INV_X1    g383(.A(G1gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT95), .Z(new_n588));
  XOR2_X1   g387(.A(new_n586), .B(KEYINPUT94), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n583), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(G8gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  XOR2_X1   g394(.A(G57gat), .B(G64gat), .Z(new_n596));
  AOI211_X1 g395(.A(new_n594), .B(new_n595), .C1(new_n596), .C2(KEYINPUT9), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(KEYINPUT97), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(KEYINPUT9), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n593), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n597), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT98), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n592), .B1(new_n602), .B2(KEYINPUT21), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(new_n214), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n603), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n607));
  XNOR2_X1  g406(.A(G155gat), .B(G183gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  INV_X1    g410(.A(G211gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n579), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT105), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n548), .A2(new_n591), .A3(new_n588), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n592), .A2(new_n547), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT18), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n592), .B2(new_n547), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n620), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n622), .B(KEYINPUT13), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT89), .B(G197gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT11), .B(G169gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT12), .Z(new_n636));
  OR2_X1    g435(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n630), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n559), .B(new_n601), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n561), .A2(new_n602), .A3(KEYINPUT10), .ZN(new_n643));
  INV_X1    g442(.A(new_n640), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(KEYINPUT10), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n642), .B1(new_n645), .B2(new_n641), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  INV_X1    g446(.A(G176gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(new_n329), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n646), .B(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n525), .A2(new_n618), .A3(new_n639), .A4(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n268), .B(KEYINPUT107), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g456(.A1(new_n654), .A2(new_n510), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n581), .B2(new_n584), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n581), .B2(new_n584), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n658), .A2(new_n584), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT42), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(KEYINPUT42), .B2(new_n660), .ZN(G1325gat));
  NOR2_X1   g462(.A1(new_n481), .A2(new_n482), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(G15gat), .B1(new_n654), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n519), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n654), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n666), .B1(G15gat), .B2(new_n668), .ZN(G1326gat));
  INV_X1    g468(.A(new_n523), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT108), .Z(new_n672));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n671), .B(KEYINPUT108), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT43), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n674), .A2(G22gat), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(G22gat), .B1(new_n674), .B2(new_n676), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(G1327gat));
  INV_X1    g478(.A(new_n579), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n488), .B2(new_n524), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n637), .A2(new_n638), .ZN(new_n682));
  INV_X1    g481(.A(new_n616), .ZN(new_n683));
  INV_X1    g482(.A(new_n651), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n535), .A3(new_n655), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT45), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(new_n525), .B2(new_n579), .ZN(new_n690));
  AOI211_X1 g489(.A(KEYINPUT44), .B(new_n680), .C1(new_n488), .C2(new_n524), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n685), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT109), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n694), .B(new_n685), .C1(new_n690), .C2(new_n691), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n655), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n688), .B1(new_n699), .B2(new_n535), .ZN(G1328gat));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n697), .B2(new_n384), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n696), .A2(KEYINPUT110), .A3(new_n510), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(G36gat), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n686), .A2(new_n536), .A3(new_n510), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT46), .Z(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(G1329gat));
  OAI21_X1  g506(.A(G43gat), .B1(new_n692), .B2(new_n519), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n686), .A2(new_n526), .A3(new_n665), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(KEYINPUT47), .A3(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT112), .Z(new_n711));
  OAI21_X1  g510(.A(G43gat), .B1(new_n697), .B2(new_n519), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT47), .B1(new_n712), .B2(new_n709), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n711), .B1(new_n715), .B2(new_n716), .ZN(G1330gat));
  OAI21_X1  g516(.A(G50gat), .B1(new_n692), .B2(new_n484), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n686), .A2(new_n454), .A3(new_n670), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(KEYINPUT48), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n523), .B1(new_n693), .B2(new_n695), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n721), .B2(new_n454), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n722), .A2(KEYINPUT113), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT113), .B1(new_n722), .B2(new_n723), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n720), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT114), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n720), .B(new_n728), .C1(new_n724), .C2(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1331gat));
  NAND4_X1  g529(.A1(new_n525), .A2(new_n618), .A3(new_n682), .A4(new_n684), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n698), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g532(.A(new_n731), .B(KEYINPUT115), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT49), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n510), .B1(new_n735), .B2(new_n366), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT116), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n366), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1333gat));
  NOR3_X1   g539(.A1(new_n731), .A2(G71gat), .A3(new_n664), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n734), .A2(new_n667), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(G71gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n670), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n639), .A2(new_n683), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n684), .B(new_n747), .C1(new_n690), .C2(new_n691), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n748), .A2(new_n206), .A3(new_n698), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT117), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n750), .A2(KEYINPUT51), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n681), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(new_n750), .A3(KEYINPUT51), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(KEYINPUT51), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n681), .A2(new_n754), .A3(new_n747), .A4(new_n751), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n753), .A2(new_n684), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n655), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n749), .B1(new_n757), .B2(new_n206), .ZN(G1336gat));
  NOR3_X1   g557(.A1(new_n748), .A2(new_n368), .A3(new_n384), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n510), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(new_n368), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT52), .ZN(G1337gat));
  NOR3_X1   g561(.A1(new_n748), .A2(new_n405), .A3(new_n519), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n756), .A2(new_n665), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n405), .ZN(G1338gat));
  INV_X1    g564(.A(new_n484), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n753), .A2(new_n684), .A3(new_n766), .A4(new_n755), .ZN(new_n767));
  OR3_X1    g566(.A1(new_n767), .A2(KEYINPUT118), .A3(G106gat), .ZN(new_n768));
  OAI21_X1  g567(.A(G106gat), .B1(new_n748), .B2(new_n523), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT118), .B1(new_n767), .B2(G106gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT53), .ZN(new_n772));
  INV_X1    g571(.A(G106gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n773), .A3(new_n766), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775));
  OAI21_X1  g574(.A(G106gat), .B1(new_n748), .B2(new_n484), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT119), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n774), .A2(KEYINPUT119), .A3(new_n775), .A4(new_n776), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n772), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT120), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n772), .A2(new_n779), .A3(new_n783), .A4(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1339gat));
  NAND2_X1  g584(.A1(new_n645), .A2(new_n641), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n650), .B1(new_n786), .B2(KEYINPUT54), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n645), .A2(new_n641), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(KEYINPUT54), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n787), .B1(new_n789), .B2(new_n786), .ZN(new_n790));
  INV_X1    g589(.A(new_n650), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n790), .A2(KEYINPUT55), .B1(new_n646), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(KEYINPUT55), .B2(new_n790), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n682), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n627), .A2(new_n628), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n621), .A2(new_n622), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n635), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n637), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n684), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n579), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n798), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n801), .A2(new_n680), .A3(new_n793), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n616), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n618), .A2(new_n682), .A3(new_n651), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n670), .B(new_n664), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n698), .A2(new_n510), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(G113gat), .B1(new_n808), .B2(new_n682), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n484), .A2(new_n485), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n803), .B2(new_n804), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n806), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n211), .A3(new_n639), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n813), .ZN(G1340gat));
  AOI21_X1  g613(.A(new_n209), .B1(new_n807), .B2(new_n684), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT121), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n812), .A2(new_n209), .A3(new_n684), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1341gat));
  AOI21_X1  g617(.A(G127gat), .B1(new_n812), .B2(new_n683), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n616), .A2(new_n214), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n807), .B2(new_n820), .ZN(G1342gat));
  NAND3_X1  g620(.A1(new_n812), .A2(new_n218), .A3(new_n579), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT56), .Z(new_n823));
  OAI21_X1  g622(.A(G134gat), .B1(new_n808), .B2(new_n680), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(G1343gat));
  XNOR2_X1  g624(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n639), .B(new_n792), .C1(new_n790), .C2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n579), .B1(new_n827), .B2(new_n799), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n616), .B1(new_n828), .B2(new_n802), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n804), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT57), .B1(new_n830), .B2(new_n523), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n519), .A2(new_n806), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n484), .B1(new_n803), .B2(new_n804), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n639), .ZN(new_n837));
  INV_X1    g636(.A(new_n232), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT58), .B1(new_n839), .B2(KEYINPUT123), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n833), .A2(new_n832), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n682), .A2(G141gat), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n837), .A2(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n840), .B(new_n843), .ZN(G1344gat));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n230), .A3(new_n684), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT124), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n833), .A2(new_n834), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n680), .A2(new_n793), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT125), .Z(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n801), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n616), .B1(new_n851), .B2(new_n828), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT57), .B1(new_n852), .B2(new_n804), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n848), .B1(new_n853), .B2(new_n670), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n684), .A3(new_n832), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n847), .B1(new_n855), .B2(G148gat), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT59), .B(new_n230), .C1(new_n836), .C2(new_n684), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n846), .B1(new_n856), .B2(new_n857), .ZN(G1345gat));
  AOI21_X1  g657(.A(G155gat), .B1(new_n841), .B2(new_n683), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n616), .A2(new_n223), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n836), .B2(new_n860), .ZN(G1346gat));
  AOI21_X1  g660(.A(G162gat), .B1(new_n841), .B2(new_n579), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n680), .A2(new_n224), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n836), .B2(new_n863), .ZN(G1347gat));
  NOR2_X1   g663(.A1(new_n655), .A2(new_n384), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n805), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(G169gat), .B1(new_n866), .B2(new_n682), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n811), .A2(new_n865), .ZN(new_n868));
  INV_X1    g667(.A(G169gat), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n639), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n867), .A2(new_n870), .ZN(G1348gat));
  NOR3_X1   g670(.A1(new_n866), .A2(new_n648), .A3(new_n651), .ZN(new_n872));
  AOI21_X1  g671(.A(G176gat), .B1(new_n868), .B2(new_n684), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(G1349gat));
  OAI21_X1  g673(.A(new_n285), .B1(new_n866), .B2(new_n616), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n868), .B(new_n683), .C1(new_n301), .C2(new_n306), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g677(.A1(new_n868), .A2(new_n273), .A3(new_n579), .ZN(new_n879));
  OAI21_X1  g678(.A(G190gat), .B1(new_n866), .B2(new_n680), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n880), .A2(KEYINPUT61), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(KEYINPUT61), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(G1351gat));
  AND2_X1   g682(.A1(new_n519), .A2(new_n865), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n833), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n328), .A3(new_n639), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n854), .A2(new_n884), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(new_n639), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n886), .B1(new_n888), .B2(new_n328), .ZN(G1352gat));
  NAND3_X1  g688(.A1(new_n885), .A2(new_n329), .A3(new_n684), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT62), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT126), .Z(new_n892));
  AND3_X1   g691(.A1(new_n854), .A2(new_n684), .A3(new_n884), .ZN(new_n893));
  OAI221_X1 g692(.A(new_n892), .B1(KEYINPUT62), .B2(new_n890), .C1(new_n329), .C2(new_n893), .ZN(G1353gat));
  NAND3_X1  g693(.A1(new_n885), .A2(new_n612), .A3(new_n683), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n854), .A2(new_n683), .A3(new_n884), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n896), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT63), .B1(new_n896), .B2(G211gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(G1354gat));
  AOI21_X1  g698(.A(G218gat), .B1(new_n885), .B2(new_n579), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n579), .A2(G218gat), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT127), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n887), .B2(new_n902), .ZN(G1355gat));
endmodule


