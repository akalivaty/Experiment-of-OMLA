

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792;

  NAND2_X1 U376 ( .A1(n397), .A2(n396), .ZN(n404) );
  XNOR2_X1 U377 ( .A(n588), .B(KEYINPUT38), .ZN(n722) );
  XNOR2_X1 U378 ( .A(n418), .B(n417), .ZN(n488) );
  XNOR2_X1 U379 ( .A(n461), .B(n460), .ZN(n779) );
  XNOR2_X1 U380 ( .A(n428), .B(KEYINPUT73), .ZN(n418) );
  NOR2_X1 U381 ( .A1(G953), .A2(KEYINPUT83), .ZN(n410) );
  OR2_X2 U382 ( .A1(n727), .A2(n360), .ZN(n419) );
  XNOR2_X2 U383 ( .A(n773), .B(n440), .ZN(n690) );
  NAND2_X1 U384 ( .A1(n611), .A2(n537), .ZN(n538) );
  XNOR2_X2 U385 ( .A(n593), .B(KEYINPUT33), .ZN(n753) );
  XNOR2_X2 U386 ( .A(n447), .B(n446), .ZN(n559) );
  XNOR2_X2 U387 ( .A(n525), .B(n524), .ZN(n780) );
  XNOR2_X2 U388 ( .A(n534), .B(KEYINPUT42), .ZN(n671) );
  INV_X1 U389 ( .A(n578), .ZN(n539) );
  XNOR2_X1 U390 ( .A(KEYINPUT4), .B(G101), .ZN(n482) );
  NAND2_X1 U391 ( .A1(n409), .A2(n403), .ZN(n395) );
  XNOR2_X1 U392 ( .A(n390), .B(n389), .ZN(n366) );
  NAND2_X1 U393 ( .A1(n420), .A2(n419), .ZN(n754) );
  XNOR2_X1 U394 ( .A(n638), .B(n637), .ZN(n713) );
  OR2_X1 U395 ( .A1(n645), .A2(KEYINPUT47), .ZN(n415) );
  INV_X1 U396 ( .A(n722), .ZN(n354) );
  OR2_X1 U397 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U398 ( .A1(n402), .A2(n400), .ZN(n399) );
  BUF_X2 U399 ( .A(n472), .Z(n774) );
  XNOR2_X1 U400 ( .A(G104), .B(G122), .ZN(n455) );
  XNOR2_X1 U401 ( .A(G140), .B(KEYINPUT106), .ZN(n452) );
  XNOR2_X1 U402 ( .A(KEYINPUT109), .B(KEYINPUT11), .ZN(n450) );
  XNOR2_X1 U403 ( .A(G140), .B(G137), .ZN(n524) );
  AND2_X2 U404 ( .A1(n398), .A2(n399), .ZN(n355) );
  AND2_X1 U405 ( .A1(n624), .A2(n584), .ZN(n542) );
  BUF_X1 U406 ( .A(n364), .Z(n699) );
  AND2_X2 U407 ( .A1(n539), .A2(n533), .ZN(n561) );
  XNOR2_X2 U408 ( .A(n575), .B(n560), .ZN(n601) );
  XNOR2_X2 U409 ( .A(n356), .B(n572), .ZN(n632) );
  XNOR2_X2 U410 ( .A(n432), .B(n431), .ZN(n773) );
  BUF_X2 U411 ( .A(n624), .Z(n356) );
  BUF_X2 U412 ( .A(n624), .Z(n357) );
  NAND2_X1 U413 ( .A1(n354), .A2(n371), .ZN(n370) );
  NOR2_X1 U414 ( .A1(n721), .A2(KEYINPUT114), .ZN(n371) );
  AND2_X1 U415 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U416 ( .A1(n721), .A2(KEYINPUT114), .ZN(n373) );
  XNOR2_X1 U417 ( .A(G113), .B(KEYINPUT3), .ZN(n417) );
  XNOR2_X2 U418 ( .A(G146), .B(G125), .ZN(n461) );
  XOR2_X1 U419 ( .A(KEYINPUT69), .B(G131), .Z(n480) );
  XNOR2_X1 U420 ( .A(n429), .B(G110), .ZN(n526) );
  XNOR2_X1 U421 ( .A(G104), .B(KEYINPUT81), .ZN(n429) );
  XNOR2_X1 U422 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U423 ( .A(n502), .B(KEYINPUT20), .ZN(n422) );
  INV_X1 U424 ( .A(KEYINPUT1), .ZN(n375) );
  XOR2_X1 U425 ( .A(G116), .B(KEYINPUT5), .Z(n487) );
  XNOR2_X1 U426 ( .A(n482), .B(G146), .ZN(n527) );
  INV_X1 U427 ( .A(KEYINPUT41), .ZN(n368) );
  NAND2_X1 U428 ( .A1(n359), .A2(n372), .ZN(n369) );
  NAND2_X1 U429 ( .A1(n423), .A2(n737), .ZN(n541) );
  AND2_X1 U430 ( .A1(n539), .A2(n540), .ZN(n423) );
  XNOR2_X1 U431 ( .A(n488), .B(n526), .ZN(n432) );
  XNOR2_X1 U432 ( .A(n463), .B(n462), .ZN(n682) );
  INV_X1 U433 ( .A(KEYINPUT92), .ZN(n405) );
  NAND2_X1 U434 ( .A1(n662), .A2(n501), .ZN(n391) );
  INV_X1 U435 ( .A(n640), .ZN(n385) );
  NAND2_X1 U436 ( .A1(n554), .A2(n553), .ZN(n712) );
  XNOR2_X1 U437 ( .A(n726), .B(n416), .ZN(n645) );
  INV_X1 U438 ( .A(KEYINPUT91), .ZN(n416) );
  NAND2_X1 U439 ( .A1(G953), .A2(G902), .ZN(n595) );
  NAND2_X1 U440 ( .A1(G953), .A2(KEYINPUT83), .ZN(n412) );
  INV_X1 U441 ( .A(KEYINPUT78), .ZN(n381) );
  INV_X1 U442 ( .A(n715), .ZN(n379) );
  AND2_X1 U443 ( .A1(n696), .A2(KEYINPUT44), .ZN(n630) );
  NAND2_X1 U444 ( .A1(n414), .A2(n411), .ZN(n485) );
  AND2_X1 U445 ( .A1(n413), .A2(n412), .ZN(n411) );
  NAND2_X1 U446 ( .A1(n410), .A2(n443), .ZN(n414) );
  NAND2_X1 U447 ( .A1(G237), .A2(KEYINPUT83), .ZN(n413) );
  XNOR2_X1 U448 ( .A(n441), .B(KEYINPUT15), .ZN(n657) );
  XNOR2_X1 U449 ( .A(G902), .B(KEYINPUT96), .ZN(n441) );
  NAND2_X1 U450 ( .A1(n422), .A2(G221), .ZN(n519) );
  NAND2_X1 U451 ( .A1(n442), .A2(n401), .ZN(n400) );
  NAND2_X1 U452 ( .A1(KEYINPUT64), .A2(KEYINPUT2), .ZN(n401) );
  NAND2_X1 U453 ( .A1(n657), .A2(KEYINPUT64), .ZN(n402) );
  INV_X1 U454 ( .A(G902), .ZN(n501) );
  INV_X1 U455 ( .A(n736), .ZN(n622) );
  XNOR2_X1 U456 ( .A(n392), .B(n491), .ZN(n662) );
  XNOR2_X1 U457 ( .A(KEYINPUT24), .B(KEYINPUT99), .ZN(n497) );
  XNOR2_X1 U458 ( .A(G119), .B(KEYINPUT23), .ZN(n492) );
  XOR2_X1 U459 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n468) );
  XNOR2_X1 U460 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n467) );
  XNOR2_X1 U461 ( .A(G122), .B(G116), .ZN(n430) );
  XNOR2_X1 U462 ( .A(n377), .B(n526), .ZN(n376) );
  NAND2_X1 U463 ( .A1(n632), .A2(n636), .ZN(n593) );
  NAND2_X1 U464 ( .A1(G234), .A2(G237), .ZN(n510) );
  INV_X1 U465 ( .A(G953), .ZN(n472) );
  NAND2_X1 U466 ( .A1(n369), .A2(n367), .ZN(n420) );
  NAND2_X1 U467 ( .A1(n421), .A2(n368), .ZN(n367) );
  INV_X1 U468 ( .A(KEYINPUT84), .ZN(n545) );
  XOR2_X1 U469 ( .A(KEYINPUT62), .B(n662), .Z(n663) );
  XNOR2_X1 U470 ( .A(n682), .B(n681), .ZN(n683) );
  INV_X1 U471 ( .A(n404), .ZN(n719) );
  INV_X1 U472 ( .A(KEYINPUT40), .ZN(n389) );
  NAND2_X1 U473 ( .A1(n644), .A2(n643), .ZN(n706) );
  XNOR2_X1 U474 ( .A(n388), .B(n387), .ZN(n698) );
  INV_X1 U475 ( .A(n712), .ZN(n394) );
  XNOR2_X1 U476 ( .A(n578), .B(n375), .ZN(n736) );
  AND2_X1 U477 ( .A1(n736), .A2(n737), .ZN(n636) );
  NAND2_X1 U478 ( .A1(n672), .A2(n647), .ZN(n358) );
  AND2_X1 U479 ( .A1(n370), .A2(n421), .ZN(n359) );
  OR2_X1 U480 ( .A1(n610), .A2(KEYINPUT41), .ZN(n360) );
  INV_X1 U481 ( .A(G237), .ZN(n443) );
  INV_X1 U482 ( .A(KEYINPUT2), .ZN(n408) );
  AND2_X1 U483 ( .A1(n442), .A2(KEYINPUT64), .ZN(n361) );
  NAND2_X1 U484 ( .A1(n355), .A2(n395), .ZN(n362) );
  NAND2_X1 U485 ( .A1(n355), .A2(n395), .ZN(n363) );
  NAND2_X1 U486 ( .A1(n355), .A2(n395), .ZN(n407) );
  AND2_X2 U487 ( .A1(n407), .A2(n404), .ZN(n364) );
  AND2_X2 U488 ( .A1(n363), .A2(n404), .ZN(n365) );
  AND2_X1 U489 ( .A1(n362), .A2(n404), .ZN(n762) );
  XNOR2_X1 U490 ( .A(n378), .B(KEYINPUT71), .ZN(n580) );
  NAND2_X1 U491 ( .A1(n660), .A2(KEYINPUT2), .ZN(n406) );
  XNOR2_X1 U492 ( .A(n406), .B(n405), .ZN(n397) );
  NAND2_X1 U493 ( .A1(n366), .A2(n671), .ZN(n550) );
  XNOR2_X1 U494 ( .A(n366), .B(G131), .ZN(G33) );
  NAND2_X1 U495 ( .A1(n372), .A2(n370), .ZN(n727) );
  NAND2_X1 U496 ( .A1(n722), .A2(KEYINPUT114), .ZN(n374) );
  XNOR2_X2 U497 ( .A(n532), .B(n531), .ZN(n578) );
  XNOR2_X1 U498 ( .A(n780), .B(n376), .ZN(n700) );
  XNOR2_X1 U499 ( .A(n530), .B(n527), .ZN(n377) );
  XNOR2_X2 U500 ( .A(n481), .B(n480), .ZN(n525) );
  XNOR2_X2 U501 ( .A(n471), .B(G134), .ZN(n481) );
  NAND2_X1 U502 ( .A1(n380), .A2(n379), .ZN(n378) );
  XNOR2_X1 U503 ( .A(n382), .B(n381), .ZN(n380) );
  NAND2_X1 U504 ( .A1(n571), .A2(n570), .ZN(n382) );
  NAND2_X1 U505 ( .A1(n383), .A2(n562), .ZN(n565) );
  NAND2_X1 U506 ( .A1(n557), .A2(n558), .ZN(n383) );
  NAND2_X1 U507 ( .A1(n384), .A2(n646), .ZN(n647) );
  NAND2_X1 U508 ( .A1(n706), .A2(n713), .ZN(n384) );
  NAND2_X1 U509 ( .A1(n385), .A2(n639), .ZN(n642) );
  NAND2_X1 U510 ( .A1(n754), .A2(n561), .ZN(n534) );
  XNOR2_X1 U511 ( .A(n386), .B(n582), .ZN(n592) );
  NAND2_X1 U512 ( .A1(n580), .A2(n581), .ZN(n386) );
  NOR2_X2 U513 ( .A1(n655), .A2(n661), .ZN(n656) );
  NAND2_X1 U514 ( .A1(n422), .A2(G217), .ZN(n507) );
  INV_X1 U515 ( .A(n767), .ZN(n396) );
  NAND2_X1 U516 ( .A1(n364), .A2(G472), .ZN(n664) );
  INV_X1 U517 ( .A(n697), .ZN(n387) );
  NAND2_X1 U518 ( .A1(n699), .A2(G217), .ZN(n388) );
  NAND2_X1 U519 ( .A1(n762), .A2(G210), .ZN(n692) );
  NAND2_X1 U520 ( .A1(n544), .A2(n543), .ZN(n546) );
  NOR2_X2 U521 ( .A1(n583), .A2(n712), .ZN(n390) );
  XNOR2_X2 U522 ( .A(n391), .B(G472), .ZN(n624) );
  XNOR2_X1 U523 ( .A(n489), .B(n490), .ZN(n392) );
  AND2_X1 U524 ( .A1(n562), .A2(n393), .ZN(n710) );
  INV_X1 U525 ( .A(n708), .ZN(n393) );
  AND2_X1 U526 ( .A1(n562), .A2(n394), .ZN(n669) );
  AND2_X2 U527 ( .A1(n601), .A2(n561), .ZN(n562) );
  INV_X1 U528 ( .A(n656), .ZN(n409) );
  NAND2_X1 U529 ( .A1(n656), .A2(n361), .ZN(n398) );
  AND2_X1 U530 ( .A1(n658), .A2(n408), .ZN(n403) );
  OR2_X2 U531 ( .A1(n700), .A2(G902), .ZN(n532) );
  NAND2_X1 U532 ( .A1(n485), .A2(G214), .ZN(n457) );
  INV_X1 U533 ( .A(n726), .ZN(n568) );
  XNOR2_X1 U534 ( .A(n415), .B(KEYINPUT79), .ZN(n569) );
  NAND2_X1 U535 ( .A1(n610), .A2(KEYINPUT41), .ZN(n421) );
  AND2_X1 U536 ( .A1(n539), .A2(n737), .ZN(n639) );
  BUF_X1 U537 ( .A(n536), .Z(n631) );
  AND2_X1 U538 ( .A1(n724), .A2(n611), .ZN(n424) );
  AND2_X1 U539 ( .A1(n588), .A2(n606), .ZN(n425) );
  XOR2_X1 U540 ( .A(n604), .B(KEYINPUT34), .Z(n426) );
  AND2_X1 U541 ( .A1(n720), .A2(n600), .ZN(n427) );
  XNOR2_X1 U542 ( .A(n609), .B(KEYINPUT66), .ZN(n626) );
  OR2_X1 U543 ( .A1(n629), .A2(n628), .ZN(n650) );
  AND2_X1 U544 ( .A1(n649), .A2(n650), .ZN(n651) );
  INV_X1 U545 ( .A(G107), .ZN(n528) );
  XNOR2_X1 U546 ( .A(n527), .B(n483), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n529), .B(n528), .ZN(n530) );
  INV_X1 U548 ( .A(KEYINPUT64), .ZN(n658) );
  BUF_X1 U549 ( .A(n661), .Z(n767) );
  INV_X1 U550 ( .A(KEYINPUT63), .ZN(n667) );
  XNOR2_X2 U551 ( .A(G119), .B(KEYINPUT72), .ZN(n428) );
  XNOR2_X1 U552 ( .A(n430), .B(G107), .ZN(n469) );
  XNOR2_X1 U553 ( .A(n469), .B(KEYINPUT16), .ZN(n431) );
  INV_X2 U554 ( .A(G143), .ZN(n433) );
  XNOR2_X2 U555 ( .A(n433), .B(G128), .ZN(n471) );
  XNOR2_X1 U556 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n434) );
  XNOR2_X1 U557 ( .A(n461), .B(n434), .ZN(n435) );
  XNOR2_X1 U558 ( .A(n471), .B(n435), .ZN(n439) );
  NAND2_X1 U559 ( .A1(n774), .A2(G224), .ZN(n436) );
  XNOR2_X1 U560 ( .A(n436), .B(KEYINPUT97), .ZN(n437) );
  XNOR2_X1 U561 ( .A(n437), .B(n482), .ZN(n438) );
  XNOR2_X1 U562 ( .A(n439), .B(n438), .ZN(n440) );
  INV_X1 U563 ( .A(n657), .ZN(n442) );
  OR2_X2 U564 ( .A1(n690), .A2(n442), .ZN(n447) );
  NAND2_X1 U565 ( .A1(n501), .A2(n443), .ZN(n448) );
  NAND2_X1 U566 ( .A1(n448), .A2(G210), .ZN(n445) );
  XNOR2_X1 U567 ( .A(KEYINPUT87), .B(KEYINPUT98), .ZN(n444) );
  BUF_X2 U568 ( .A(n559), .Z(n588) );
  NAND2_X1 U569 ( .A1(n448), .A2(G214), .ZN(n584) );
  INV_X1 U570 ( .A(n584), .ZN(n721) );
  XNOR2_X1 U571 ( .A(G143), .B(G113), .ZN(n449) );
  XNOR2_X1 U572 ( .A(n450), .B(n449), .ZN(n454) );
  XNOR2_X1 U573 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n451) );
  XNOR2_X1 U574 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U575 ( .A(n454), .B(n453), .ZN(n459) );
  XNOR2_X1 U576 ( .A(n455), .B(KEYINPUT12), .ZN(n456) );
  XNOR2_X1 U577 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U578 ( .A(n459), .B(n458), .ZN(n463) );
  XNOR2_X1 U579 ( .A(KEYINPUT68), .B(KEYINPUT10), .ZN(n460) );
  XNOR2_X1 U580 ( .A(n480), .B(n779), .ZN(n462) );
  NAND2_X1 U581 ( .A1(n682), .A2(n501), .ZN(n466) );
  INV_X1 U582 ( .A(KEYINPUT13), .ZN(n464) );
  XNOR2_X1 U583 ( .A(n464), .B(G475), .ZN(n465) );
  XNOR2_X1 U584 ( .A(n466), .B(n465), .ZN(n554) );
  INV_X1 U585 ( .A(n554), .ZN(n479) );
  XNOR2_X1 U586 ( .A(n468), .B(n467), .ZN(n470) );
  XNOR2_X1 U587 ( .A(n470), .B(n469), .ZN(n476) );
  AND2_X1 U588 ( .A1(G234), .A2(n472), .ZN(n473) );
  XNOR2_X1 U589 ( .A(n473), .B(KEYINPUT8), .ZN(n494) );
  NAND2_X1 U590 ( .A1(n494), .A2(G217), .ZN(n474) );
  XNOR2_X1 U591 ( .A(n481), .B(n474), .ZN(n475) );
  XNOR2_X1 U592 ( .A(n476), .B(n475), .ZN(n764) );
  NAND2_X1 U593 ( .A1(n764), .A2(n501), .ZN(n478) );
  INV_X1 U594 ( .A(G478), .ZN(n477) );
  XNOR2_X1 U595 ( .A(n478), .B(n477), .ZN(n553) );
  NAND2_X1 U596 ( .A1(n479), .A2(n553), .ZN(n610) );
  XOR2_X1 U597 ( .A(KEYINPUT80), .B(KEYINPUT105), .Z(n483) );
  XNOR2_X1 U598 ( .A(n525), .B(n484), .ZN(n491) );
  NAND2_X1 U599 ( .A1(n485), .A2(G210), .ZN(n486) );
  XNOR2_X1 U600 ( .A(n487), .B(n486), .ZN(n490) );
  XNOR2_X1 U601 ( .A(n488), .B(G137), .ZN(n489) );
  XNOR2_X1 U602 ( .A(G110), .B(G128), .ZN(n493) );
  XNOR2_X1 U603 ( .A(n493), .B(n492), .ZN(n496) );
  NAND2_X1 U604 ( .A1(n494), .A2(G221), .ZN(n495) );
  XNOR2_X1 U605 ( .A(n496), .B(n495), .ZN(n500) );
  XNOR2_X1 U606 ( .A(n524), .B(n497), .ZN(n498) );
  XNOR2_X1 U607 ( .A(n779), .B(n498), .ZN(n499) );
  XNOR2_X1 U608 ( .A(n500), .B(n499), .ZN(n697) );
  NAND2_X1 U609 ( .A1(n697), .A2(n501), .ZN(n509) );
  NAND2_X1 U610 ( .A1(n657), .A2(G234), .ZN(n502) );
  INV_X1 U611 ( .A(KEYINPUT100), .ZN(n503) );
  XNOR2_X1 U612 ( .A(n503), .B(KEYINPUT101), .ZN(n505) );
  XNOR2_X1 U613 ( .A(KEYINPUT25), .B(KEYINPUT86), .ZN(n504) );
  XNOR2_X1 U614 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U615 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U616 ( .A(n509), .B(n508), .ZN(n536) );
  XNOR2_X1 U617 ( .A(n510), .B(KEYINPUT14), .ZN(n720) );
  INV_X1 U618 ( .A(n720), .ZN(n511) );
  NOR2_X1 U619 ( .A1(n511), .A2(n595), .ZN(n512) );
  XNOR2_X1 U620 ( .A(n512), .B(KEYINPUT113), .ZN(n513) );
  NOR2_X1 U621 ( .A1(G900), .A2(n513), .ZN(n515) );
  AND2_X1 U622 ( .A1(n774), .A2(G952), .ZN(n594) );
  AND2_X1 U623 ( .A1(n720), .A2(n594), .ZN(n514) );
  OR2_X1 U624 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U625 ( .A(n516), .B(KEYINPUT88), .ZN(n540) );
  INV_X1 U626 ( .A(KEYINPUT102), .ZN(n517) );
  XNOR2_X1 U627 ( .A(n517), .B(KEYINPUT21), .ZN(n518) );
  XNOR2_X2 U628 ( .A(n519), .B(n518), .ZN(n732) );
  AND2_X1 U629 ( .A1(n540), .A2(n732), .ZN(n520) );
  NAND2_X1 U630 ( .A1(n631), .A2(n520), .ZN(n573) );
  INV_X1 U631 ( .A(n573), .ZN(n521) );
  NAND2_X1 U632 ( .A1(n357), .A2(n521), .ZN(n523) );
  INV_X1 U633 ( .A(KEYINPUT28), .ZN(n522) );
  XNOR2_X1 U634 ( .A(n523), .B(n522), .ZN(n533) );
  NAND2_X1 U635 ( .A1(G227), .A2(n774), .ZN(n529) );
  INV_X1 U636 ( .A(G469), .ZN(n531) );
  XNOR2_X1 U637 ( .A(n732), .B(KEYINPUT103), .ZN(n535) );
  INV_X1 U638 ( .A(n535), .ZN(n611) );
  INV_X1 U639 ( .A(n536), .ZN(n537) );
  XNOR2_X2 U640 ( .A(n538), .B(KEYINPUT67), .ZN(n737) );
  XNOR2_X1 U641 ( .A(n541), .B(KEYINPUT85), .ZN(n544) );
  XNOR2_X1 U642 ( .A(n542), .B(KEYINPUT30), .ZN(n543) );
  XNOR2_X2 U643 ( .A(n546), .B(n545), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n552), .A2(n354), .ZN(n548) );
  INV_X1 U645 ( .A(KEYINPUT39), .ZN(n547) );
  XNOR2_X1 U646 ( .A(n548), .B(n547), .ZN(n583) );
  INV_X1 U647 ( .A(KEYINPUT46), .ZN(n549) );
  XNOR2_X1 U648 ( .A(n550), .B(n549), .ZN(n581) );
  INV_X1 U649 ( .A(n553), .ZN(n551) );
  AND2_X1 U650 ( .A1(n551), .A2(n554), .ZN(n606) );
  NAND2_X1 U651 ( .A1(n552), .A2(n425), .ZN(n688) );
  XNOR2_X2 U652 ( .A(n555), .B(KEYINPUT112), .ZN(n708) );
  AND2_X2 U653 ( .A1(n708), .A2(n712), .ZN(n726) );
  INV_X1 U654 ( .A(KEYINPUT47), .ZN(n563) );
  NOR2_X1 U655 ( .A1(n563), .A2(KEYINPUT90), .ZN(n556) );
  NAND2_X1 U656 ( .A1(n726), .A2(n556), .ZN(n558) );
  NAND2_X1 U657 ( .A1(n568), .A2(KEYINPUT90), .ZN(n557) );
  AND2_X2 U658 ( .A1(n559), .A2(n584), .ZN(n575) );
  INV_X1 U659 ( .A(KEYINPUT19), .ZN(n560) );
  NAND2_X1 U660 ( .A1(n563), .A2(KEYINPUT90), .ZN(n564) );
  NAND2_X1 U661 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U662 ( .A1(n688), .A2(n566), .ZN(n567) );
  XNOR2_X1 U663 ( .A(n567), .B(KEYINPUT89), .ZN(n571) );
  NAND2_X1 U664 ( .A1(n569), .A2(n562), .ZN(n570) );
  INV_X1 U665 ( .A(KEYINPUT6), .ZN(n572) );
  NOR2_X1 U666 ( .A1(n712), .A2(n573), .ZN(n574) );
  AND2_X1 U667 ( .A1(n632), .A2(n574), .ZN(n586) );
  NAND2_X1 U668 ( .A1(n586), .A2(n575), .ZN(n577) );
  INV_X1 U669 ( .A(KEYINPUT36), .ZN(n576) );
  XNOR2_X1 U670 ( .A(n577), .B(n576), .ZN(n579) );
  XNOR2_X1 U671 ( .A(n622), .B(KEYINPUT95), .ZN(n615) );
  AND2_X1 U672 ( .A1(n579), .A2(n615), .ZN(n715) );
  XOR2_X1 U673 ( .A(KEYINPUT70), .B(KEYINPUT48), .Z(n582) );
  OR2_X1 U674 ( .A1(n583), .A2(n708), .ZN(n680) );
  AND2_X1 U675 ( .A1(n622), .A2(n584), .ZN(n585) );
  NAND2_X1 U676 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U677 ( .A(n587), .B(KEYINPUT43), .ZN(n590) );
  INV_X1 U678 ( .A(n588), .ZN(n589) );
  NAND2_X1 U679 ( .A1(n590), .A2(n589), .ZN(n670) );
  AND2_X1 U680 ( .A1(n680), .A2(n670), .ZN(n591) );
  NAND2_X1 U681 ( .A1(n592), .A2(n591), .ZN(n659) );
  XNOR2_X1 U682 ( .A(n659), .B(KEYINPUT82), .ZN(n655) );
  INV_X1 U683 ( .A(n594), .ZN(n599) );
  INV_X1 U684 ( .A(G898), .ZN(n597) );
  INV_X1 U685 ( .A(n595), .ZN(n596) );
  NAND2_X1 U686 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U687 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U688 ( .A1(n601), .A2(n427), .ZN(n603) );
  INV_X1 U689 ( .A(KEYINPUT0), .ZN(n602) );
  XNOR2_X2 U690 ( .A(n603), .B(n602), .ZN(n635) );
  NAND2_X1 U691 ( .A1(n635), .A2(n753), .ZN(n605) );
  INV_X1 U692 ( .A(KEYINPUT75), .ZN(n604) );
  XNOR2_X1 U693 ( .A(n605), .B(n426), .ZN(n607) );
  NAND2_X1 U694 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X2 U695 ( .A(n608), .B(KEYINPUT35), .ZN(n696) );
  NOR2_X2 U696 ( .A1(n696), .A2(KEYINPUT44), .ZN(n609) );
  INV_X1 U697 ( .A(n610), .ZN(n724) );
  NAND2_X1 U698 ( .A1(n635), .A2(n424), .ZN(n614) );
  XNOR2_X1 U699 ( .A(KEYINPUT77), .B(KEYINPUT22), .ZN(n612) );
  XNOR2_X1 U700 ( .A(n612), .B(KEYINPUT76), .ZN(n613) );
  XNOR2_X1 U701 ( .A(n614), .B(n613), .ZN(n623) );
  INV_X1 U702 ( .A(n631), .ZN(n733) );
  OR2_X1 U703 ( .A1(n632), .A2(n733), .ZN(n617) );
  INV_X1 U704 ( .A(n615), .ZN(n616) );
  NOR2_X1 U705 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U706 ( .A1(n623), .A2(n618), .ZN(n621) );
  INV_X1 U707 ( .A(KEYINPUT65), .ZN(n619) );
  XNOR2_X1 U708 ( .A(n619), .B(KEYINPUT32), .ZN(n620) );
  XNOR2_X1 U709 ( .A(n621), .B(n620), .ZN(n678) );
  AND2_X1 U710 ( .A1(n622), .A2(n623), .ZN(n634) );
  NOR2_X1 U711 ( .A1(n356), .A2(n733), .ZN(n625) );
  NAND2_X1 U712 ( .A1(n634), .A2(n625), .ZN(n673) );
  AND2_X1 U713 ( .A1(n678), .A2(n673), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n626), .A2(n629), .ZN(n627) );
  XNOR2_X1 U715 ( .A(n627), .B(KEYINPUT74), .ZN(n652) );
  INV_X1 U716 ( .A(KEYINPUT44), .ZN(n628) );
  XNOR2_X1 U717 ( .A(n630), .B(KEYINPUT94), .ZN(n648) );
  NOR2_X1 U718 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n672) );
  INV_X1 U720 ( .A(n635), .ZN(n640) );
  NAND2_X1 U721 ( .A1(n636), .A2(n357), .ZN(n742) );
  OR2_X1 U722 ( .A1(n640), .A2(n742), .ZN(n638) );
  INV_X1 U723 ( .A(KEYINPUT31), .ZN(n637) );
  INV_X1 U724 ( .A(KEYINPUT104), .ZN(n641) );
  XNOR2_X1 U725 ( .A(n642), .B(n641), .ZN(n644) );
  INV_X1 U726 ( .A(n357), .ZN(n643) );
  INV_X1 U727 ( .A(n645), .ZN(n646) );
  NOR2_X1 U728 ( .A1(n648), .A2(n358), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n654) );
  INV_X1 U730 ( .A(KEYINPUT45), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n654), .B(n653), .ZN(n661) );
  BUF_X2 U732 ( .A(n659), .Z(n787) );
  INV_X1 U733 ( .A(n787), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n664), .B(n663), .ZN(n666) );
  INV_X1 U735 ( .A(G952), .ZN(n665) );
  AND2_X1 U736 ( .A1(n665), .A2(G953), .ZN(n766) );
  NOR2_X2 U737 ( .A1(n666), .A2(n766), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(G57) );
  XOR2_X1 U739 ( .A(G146), .B(n669), .Z(G48) );
  XNOR2_X1 U740 ( .A(n670), .B(G140), .ZN(G42) );
  XNOR2_X1 U741 ( .A(n671), .B(G137), .ZN(G39) );
  XNOR2_X1 U742 ( .A(n672), .B(G101), .ZN(G3) );
  XNOR2_X1 U743 ( .A(n673), .B(G110), .ZN(G12) );
  NOR2_X1 U744 ( .A1(n706), .A2(n708), .ZN(n677) );
  XOR2_X1 U745 ( .A(KEYINPUT115), .B(KEYINPUT26), .Z(n675) );
  XNOR2_X1 U746 ( .A(G107), .B(KEYINPUT27), .ZN(n674) );
  XNOR2_X1 U747 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n677), .B(n676), .ZN(G9) );
  XNOR2_X1 U749 ( .A(n678), .B(G119), .ZN(G21) );
  NOR2_X1 U750 ( .A1(n713), .A2(n708), .ZN(n679) );
  XOR2_X1 U751 ( .A(G116), .B(n679), .Z(G18) );
  XNOR2_X1 U752 ( .A(n680), .B(G134), .ZN(G36) );
  NAND2_X1 U753 ( .A1(n365), .A2(G475), .ZN(n684) );
  XNOR2_X1 U754 ( .A(KEYINPUT122), .B(KEYINPUT59), .ZN(n681) );
  XNOR2_X1 U755 ( .A(n684), .B(n683), .ZN(n685) );
  NOR2_X2 U756 ( .A1(n685), .A2(n766), .ZN(n687) );
  XOR2_X1 U757 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n686) );
  XNOR2_X1 U758 ( .A(n687), .B(n686), .ZN(G60) );
  XNOR2_X1 U759 ( .A(n688), .B(G143), .ZN(G45) );
  XOR2_X1 U760 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n689) );
  XNOR2_X1 U761 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U762 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X2 U763 ( .A1(n693), .A2(n766), .ZN(n695) );
  XOR2_X1 U764 ( .A(KEYINPUT93), .B(KEYINPUT56), .Z(n694) );
  XNOR2_X1 U765 ( .A(n695), .B(n694), .ZN(G51) );
  XOR2_X1 U766 ( .A(n696), .B(G122), .Z(G24) );
  NOR2_X1 U767 ( .A1(n698), .A2(n766), .ZN(G66) );
  NAND2_X1 U768 ( .A1(n699), .A2(G469), .ZN(n704) );
  BUF_X1 U769 ( .A(n700), .Z(n702) );
  XOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n701) );
  XNOR2_X1 U771 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U772 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U773 ( .A1(n705), .A2(n766), .ZN(G54) );
  NOR2_X1 U774 ( .A1(n706), .A2(n712), .ZN(n707) );
  XOR2_X1 U775 ( .A(G104), .B(n707), .Z(G6) );
  XNOR2_X1 U776 ( .A(KEYINPUT116), .B(KEYINPUT29), .ZN(n709) );
  XNOR2_X1 U777 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U778 ( .A(G128), .B(n711), .ZN(G30) );
  NOR2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U780 ( .A(G113), .B(n714), .Z(G15) );
  XNOR2_X1 U781 ( .A(G125), .B(n715), .ZN(n716) );
  XNOR2_X1 U782 ( .A(n716), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U783 ( .A1(n767), .A2(n787), .ZN(n717) );
  NOR2_X1 U784 ( .A1(n717), .A2(KEYINPUT2), .ZN(n718) );
  NOR2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n759) );
  NAND2_X1 U786 ( .A1(G952), .A2(n720), .ZN(n752) );
  NAND2_X1 U787 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U788 ( .A(KEYINPUT119), .B(n723), .Z(n725) );
  NAND2_X1 U789 ( .A1(n725), .A2(n724), .ZN(n729) );
  OR2_X1 U790 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U791 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U792 ( .A1(n730), .A2(n753), .ZN(n731) );
  XOR2_X1 U793 ( .A(KEYINPUT120), .B(n731), .Z(n749) );
  NOR2_X1 U794 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U795 ( .A(KEYINPUT49), .B(n734), .Z(n735) );
  NOR2_X1 U796 ( .A1(n356), .A2(n735), .ZN(n741) );
  NOR2_X1 U797 ( .A1(n737), .A2(n736), .ZN(n739) );
  XNOR2_X1 U798 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n738) );
  XNOR2_X1 U799 ( .A(n739), .B(n738), .ZN(n740) );
  NAND2_X1 U800 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U801 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U802 ( .A(n744), .B(KEYINPUT118), .ZN(n745) );
  XNOR2_X1 U803 ( .A(n745), .B(KEYINPUT51), .ZN(n747) );
  INV_X1 U804 ( .A(n754), .ZN(n746) );
  NOR2_X1 U805 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U806 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U807 ( .A(n750), .B(KEYINPUT52), .ZN(n751) );
  NOR2_X1 U808 ( .A1(n752), .A2(n751), .ZN(n756) );
  AND2_X1 U809 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U811 ( .A(n757), .B(KEYINPUT121), .ZN(n758) );
  NOR2_X1 U812 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U813 ( .A1(n774), .A2(n760), .ZN(n761) );
  XOR2_X1 U814 ( .A(KEYINPUT53), .B(n761), .Z(G75) );
  NAND2_X1 U815 ( .A1(n365), .A2(G478), .ZN(n763) );
  XOR2_X1 U816 ( .A(n764), .B(n763), .Z(n765) );
  NOR2_X1 U817 ( .A1(n766), .A2(n765), .ZN(G63) );
  NAND2_X1 U818 ( .A1(n396), .A2(n774), .ZN(n771) );
  NAND2_X1 U819 ( .A1(G953), .A2(G224), .ZN(n768) );
  XNOR2_X1 U820 ( .A(KEYINPUT61), .B(n768), .ZN(n769) );
  NAND2_X1 U821 ( .A1(n769), .A2(G898), .ZN(n770) );
  NAND2_X1 U822 ( .A1(n771), .A2(n770), .ZN(n778) );
  XNOR2_X1 U823 ( .A(G101), .B(KEYINPUT124), .ZN(n772) );
  XNOR2_X1 U824 ( .A(n773), .B(n772), .ZN(n776) );
  NOR2_X1 U825 ( .A1(G898), .A2(n774), .ZN(n775) );
  NOR2_X1 U826 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U827 ( .A(n778), .B(n777), .ZN(G69) );
  XNOR2_X1 U828 ( .A(n779), .B(KEYINPUT4), .ZN(n782) );
  INV_X1 U829 ( .A(n780), .ZN(n781) );
  XNOR2_X1 U830 ( .A(n782), .B(n781), .ZN(n786) );
  XOR2_X1 U831 ( .A(G227), .B(n786), .Z(n783) );
  NAND2_X1 U832 ( .A1(n783), .A2(G900), .ZN(n784) );
  NAND2_X1 U833 ( .A1(G953), .A2(n784), .ZN(n785) );
  XOR2_X1 U834 ( .A(KEYINPUT126), .B(n785), .Z(n791) );
  XNOR2_X1 U835 ( .A(n787), .B(n786), .ZN(n788) );
  NOR2_X1 U836 ( .A1(n788), .A2(G953), .ZN(n789) );
  XOR2_X1 U837 ( .A(KEYINPUT125), .B(n789), .Z(n790) );
  NOR2_X1 U838 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U839 ( .A(KEYINPUT127), .B(n792), .ZN(G72) );
endmodule

