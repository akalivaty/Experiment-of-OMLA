//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  AND2_X1   g002(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n205));
  OAI211_X1 g004(.A(new_n202), .B(new_n203), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(KEYINPUT67), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(new_n204), .B2(new_n205), .ZN(new_n211));
  AOI21_X1  g010(.A(G190gat), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n206), .B1(new_n212), .B2(new_n202), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT68), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT26), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(KEYINPUT68), .B(new_n206), .C1(new_n212), .C2(new_n202), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n215), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(KEYINPUT24), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(KEYINPUT65), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n216), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n216), .A2(new_n226), .ZN(new_n231));
  NOR2_X1   g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g032(.A(KEYINPUT66), .B(new_n216), .C1(new_n225), .C2(new_n227), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n218), .B(KEYINPUT23), .Z(new_n236));
  XOR2_X1   g035(.A(new_n220), .B(KEYINPUT64), .Z(new_n237));
  NAND4_X1  g036(.A1(new_n235), .A2(KEYINPUT25), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n220), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n217), .A2(KEYINPUT24), .ZN(new_n241));
  NOR3_X1   g040(.A1(new_n241), .A2(new_n232), .A3(new_n231), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT29), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G211gat), .B(G218gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(KEYINPUT72), .ZN(new_n251));
  XNOR2_X1  g050(.A(G197gat), .B(G204gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT22), .ZN(new_n253));
  INV_X1    g052(.A(G211gat), .ZN(new_n254));
  INV_X1    g053(.A(G218gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n256), .B(new_n252), .C1(new_n250), .C2(KEYINPUT72), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n258), .A2(KEYINPUT73), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT73), .B1(new_n258), .B2(new_n259), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n248), .B1(new_n223), .B2(new_n244), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT75), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT75), .ZN(new_n266));
  AOI211_X1 g065(.A(new_n266), .B(new_n248), .C1(new_n223), .C2(new_n244), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n249), .B(new_n263), .C1(new_n265), .C2(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(KEYINPUT74), .B(KEYINPUT29), .Z(new_n269));
  AOI22_X1  g068(.A1(new_n245), .A2(new_n269), .B1(G226gat), .B2(G233gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n262), .B1(new_n270), .B2(new_n264), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT30), .ZN(new_n273));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  OR3_X1    g075(.A1(new_n272), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n276), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n273), .B1(new_n272), .B2(new_n276), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G1gat), .B(G29gat), .ZN(new_n282));
  INV_X1    g081(.A(G85gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT0), .B(G57gat), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G225gat), .A2(G233gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT2), .ZN(new_n290));
  INV_X1    g089(.A(G155gat), .ZN(new_n291));
  INV_X1    g090(.A(G162gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G141gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n295), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n291), .A2(new_n292), .ZN(new_n304));
  XNOR2_X1  g103(.A(G141gat), .B(G148gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n294), .B(new_n304), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT69), .ZN(new_n311));
  XNOR2_X1  g110(.A(G113gat), .B(G120gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G127gat), .B(G134gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n315));
  INV_X1    g114(.A(G120gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G113gat), .ZN(new_n317));
  INV_X1    g116(.A(G113gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G120gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n317), .A2(new_n319), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n314), .A2(new_n315), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n317), .A2(new_n319), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(new_n320), .A3(new_n315), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n313), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n289), .B1(new_n310), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n331));
  AND2_X1   g130(.A1(G127gat), .A2(G134gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(G127gat), .A2(G134gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT69), .B1(new_n324), .B2(new_n334), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n335), .A2(KEYINPUT1), .A3(new_n321), .ZN(new_n336));
  INV_X1    g135(.A(new_n326), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n331), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT71), .A3(new_n326), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n341));
  INV_X1    g140(.A(new_n299), .ZN(new_n342));
  OAI21_X1  g141(.A(G141gat), .B1(new_n342), .B2(new_n297), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n343), .A2(new_n301), .B1(new_n294), .B2(new_n293), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n304), .A2(new_n294), .ZN(new_n345));
  XOR2_X1   g144(.A(G141gat), .B(G148gat), .Z(new_n346));
  NAND2_X1  g145(.A1(new_n290), .A2(KEYINPUT76), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT2), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n345), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n341), .B1(new_n344), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n303), .A2(new_n307), .A3(KEYINPUT78), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n330), .B1(new_n340), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n344), .A2(new_n351), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n330), .B(new_n356), .C1(new_n336), .C2(new_n337), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT79), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n327), .A2(new_n359), .A3(new_n330), .A4(new_n356), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n329), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n365));
  XNOR2_X1  g164(.A(new_n327), .B(new_n356), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n366), .B2(new_n289), .ZN(new_n367));
  OAI211_X1 g166(.A(KEYINPUT80), .B(new_n329), .C1(new_n355), .C2(new_n361), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n364), .A2(KEYINPUT82), .A3(new_n367), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n323), .A2(KEYINPUT71), .A3(new_n326), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT71), .B1(new_n323), .B2(new_n326), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n330), .B(new_n354), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT83), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n340), .A2(new_n378), .A3(new_n330), .A4(new_n354), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT4), .B1(new_n328), .B2(new_n308), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(new_n365), .A3(new_n329), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n287), .B1(new_n373), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n382), .ZN(new_n384));
  AOI211_X1 g183(.A(new_n286), .B(new_n384), .C1(new_n371), .C2(new_n372), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n383), .A2(new_n385), .A3(KEYINPUT6), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n373), .A2(new_n382), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(KEYINPUT6), .A3(new_n286), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n281), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n269), .B1(new_n308), .B2(KEYINPUT3), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n262), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n258), .B2(new_n259), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n308), .B1(new_n394), .B2(KEYINPUT3), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n257), .A2(new_n250), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n269), .B1(new_n257), .B2(new_n250), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n309), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n352), .A3(new_n353), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n393), .B1(new_n392), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT87), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT87), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n352), .A2(new_n353), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n405), .A2(new_n399), .B1(new_n262), .B2(new_n391), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n403), .B(new_n404), .C1(new_n406), .C2(new_n393), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(G22gat), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n403), .B1(new_n406), .B2(new_n393), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT88), .B1(new_n409), .B2(G22gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n402), .A2(new_n407), .A3(KEYINPUT88), .A4(G22gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(G78gat), .B(G106gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G50gat), .ZN(new_n414));
  XOR2_X1   g213(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n409), .A2(G22gat), .ZN(new_n418));
  OAI21_X1  g217(.A(G22gat), .B1(new_n396), .B2(new_n401), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT86), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n409), .A2(KEYINPUT86), .A3(G22gat), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n416), .B(KEYINPUT85), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT40), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n310), .A2(new_n328), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n381), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n289), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n287), .B1(new_n431), .B2(KEYINPUT39), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n288), .B1(new_n381), .B2(new_n429), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT39), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n366), .A2(new_n289), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n428), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n431), .B(KEYINPUT39), .C1(new_n289), .C2(new_n366), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n286), .B1(new_n433), .B2(new_n434), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(KEYINPUT40), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(new_n383), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n427), .B1(new_n442), .B2(new_n280), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n387), .A2(new_n286), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n384), .B1(new_n371), .B2(new_n372), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT6), .B1(new_n445), .B2(new_n287), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT38), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT37), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n268), .A2(new_n449), .A3(new_n271), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n450), .A2(new_n276), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n272), .A2(KEYINPUT37), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n276), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n249), .B(new_n262), .C1(new_n265), .C2(new_n267), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n263), .B1(new_n270), .B2(new_n264), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(KEYINPUT37), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n448), .ZN(new_n458));
  OAI22_X1  g257(.A1(new_n454), .A2(new_n458), .B1(new_n272), .B2(new_n276), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n447), .A2(new_n388), .A3(new_n460), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n390), .A2(new_n427), .B1(new_n443), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G227gat), .A2(G233gat), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n245), .A2(new_n338), .A3(new_n339), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n340), .A2(new_n223), .A3(new_n244), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT32), .ZN(new_n467));
  OR3_X1    g266(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT34), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT34), .B1(new_n466), .B2(new_n467), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n464), .A2(new_n463), .A3(new_n465), .ZN(new_n471));
  XNOR2_X1  g270(.A(G15gat), .B(G43gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(G71gat), .B(G99gat), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n472), .B(new_n473), .Z(new_n474));
  OAI211_X1 g273(.A(new_n471), .B(new_n474), .C1(new_n466), .C2(KEYINPUT33), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n464), .A2(new_n465), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT33), .ZN(new_n477));
  INV_X1    g276(.A(new_n474), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n476), .B(new_n463), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n468), .A2(new_n475), .A3(new_n479), .A4(new_n469), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT36), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n426), .A2(new_n481), .A3(new_n483), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n487), .A2(new_n280), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT89), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n488), .B(new_n492), .C1(new_n386), .C2(new_n389), .ZN(new_n493));
  NOR2_X1   g292(.A1(KEYINPUT89), .A2(KEYINPUT35), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n491), .B1(new_n447), .B2(new_n388), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n494), .A3(new_n488), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n462), .A2(new_n486), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500));
  INV_X1    g299(.A(G1gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT16), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(G1gat), .B2(new_n500), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n504), .B(G8gat), .Z(new_n505));
  INV_X1    g304(.A(G43gat), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n506), .A2(G50gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(G50gat), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT15), .ZN(new_n509));
  NAND2_X1  g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR3_X1   g311(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(KEYINPUT94), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n510), .B1(new_n516), .B2(new_n513), .ZN(new_n517));
  AOI211_X1 g316(.A(new_n517), .B(new_n509), .C1(new_n513), .C2(new_n516), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT92), .B(G50gat), .Z(new_n519));
  OAI21_X1  g318(.A(new_n507), .B1(new_n519), .B2(G43gat), .ZN(new_n520));
  XOR2_X1   g319(.A(KEYINPUT91), .B(KEYINPUT15), .Z(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n522), .A2(KEYINPUT93), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(KEYINPUT93), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT95), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n527), .B(new_n518), .C1(new_n523), .C2(new_n524), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n515), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI211_X1 g330(.A(KEYINPUT17), .B(new_n515), .C1(new_n526), .C2(new_n528), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n505), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n529), .A2(new_n505), .ZN(new_n534));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n529), .B(new_n505), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n535), .B(KEYINPUT13), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n533), .A2(KEYINPUT18), .A3(new_n534), .A4(new_n535), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n544));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G169gat), .B(G197gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT12), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n538), .A2(new_n541), .A3(new_n542), .A4(new_n549), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G71gat), .ZN(new_n554));
  INV_X1    g353(.A(G78gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT96), .ZN(new_n557));
  XNOR2_X1  g356(.A(G57gat), .B(G64gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT9), .ZN(new_n559));
  OAI22_X1  g358(.A1(new_n558), .A2(new_n559), .B1(new_n554), .B2(new_n555), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(G64gat), .B1(KEYINPUT97), .B2(G57gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(KEYINPUT98), .A2(G57gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(KEYINPUT97), .A2(KEYINPUT98), .A3(G57gat), .A4(G64gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n556), .A2(new_n559), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n554), .A2(new_n555), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G92gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT100), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n283), .B(new_n571), .C1(new_n572), .C2(KEYINPUT7), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n572), .B2(KEYINPUT7), .ZN(new_n574));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT8), .A2(new_n575), .B1(new_n283), .B2(new_n571), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  OAI211_X1 g376(.A(KEYINPUT100), .B(new_n577), .C1(new_n283), .C2(new_n571), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G99gat), .B(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n574), .A2(new_n580), .A3(new_n576), .A4(new_n578), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n582), .A2(KEYINPUT101), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT101), .B1(new_n582), .B2(new_n583), .ZN(new_n585));
  OAI211_X1 g384(.A(KEYINPUT10), .B(new_n570), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n583), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n569), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n583), .A3(new_n582), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT10), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n588), .B2(new_n589), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT104), .ZN(new_n597));
  XNOR2_X1  g396(.A(G120gat), .B(G148gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  OR3_X1    g399(.A1(new_n595), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT105), .B1(new_n592), .B2(new_n593), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT105), .ZN(new_n603));
  INV_X1    g402(.A(new_n593), .ZN(new_n604));
  AOI211_X1 g403(.A(new_n603), .B(new_n604), .C1(new_n586), .C2(new_n591), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n597), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n600), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n553), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT21), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n505), .B1(new_n611), .B2(new_n569), .ZN(new_n612));
  INV_X1    g411(.A(G183gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G127gat), .B(G155gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT99), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n616), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n569), .A2(new_n611), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n254), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n621), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n620), .B(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n584), .A2(new_n585), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n529), .B2(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n628), .A2(KEYINPUT102), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n531), .B2(new_n532), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(KEYINPUT102), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G190gat), .B(G218gat), .Z(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT103), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n633), .A2(KEYINPUT103), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n632), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n639), .B1(new_n632), .B2(new_n634), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n625), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n499), .A2(new_n610), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n386), .A2(new_n389), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n280), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(G8gat), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n650), .A2(KEYINPUT106), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(KEYINPUT106), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT16), .B(G8gat), .Z(new_n653));
  NAND3_X1  g452(.A1(new_n645), .A2(new_n280), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n656));
  OAI22_X1  g455(.A1(new_n651), .A2(new_n652), .B1(new_n655), .B2(new_n656), .ZN(G1325gat));
  AOI21_X1  g456(.A(G15gat), .B1(new_n645), .B2(new_n485), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n486), .A2(KEYINPUT107), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n486), .A2(KEYINPUT107), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n661), .A2(G15gat), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n658), .B1(new_n645), .B2(new_n662), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n427), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT43), .B(G22gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  OAI21_X1  g465(.A(KEYINPUT44), .B1(new_n499), .B2(new_n643), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n447), .A2(new_n388), .A3(new_n460), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n444), .A2(new_n437), .A3(new_n440), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n426), .B1(new_n669), .B2(new_n281), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n280), .B1(new_n447), .B2(new_n388), .ZN(new_n671));
  OAI22_X1  g470(.A1(new_n668), .A2(new_n670), .B1(new_n671), .B2(new_n426), .ZN(new_n672));
  INV_X1    g471(.A(new_n486), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n493), .A2(new_n495), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n494), .B1(new_n497), .B2(new_n488), .ZN(new_n675));
  OAI22_X1  g474(.A1(new_n672), .A2(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n641), .B2(new_n642), .ZN(new_n679));
  INV_X1    g478(.A(new_n642), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n640), .A3(KEYINPUT109), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n676), .A2(new_n677), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n610), .A2(new_n625), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n646), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n687), .A2(KEYINPUT110), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT110), .B1(new_n687), .B2(new_n688), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(G29gat), .A3(new_n690), .ZN(new_n691));
  OAI221_X1 g490(.A(new_n486), .B1(new_n671), .B2(new_n426), .C1(new_n668), .C2(new_n670), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n496), .A2(new_n498), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n643), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n694), .A2(new_n686), .ZN(new_n695));
  INV_X1    g494(.A(G29gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(new_n646), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n691), .A2(new_n699), .ZN(G1328gat));
  INV_X1    g499(.A(G36gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n695), .A2(new_n701), .A3(new_n280), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT46), .Z(new_n703));
  OAI21_X1  g502(.A(G36gat), .B1(new_n687), .B2(new_n281), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1329gat));
  OAI21_X1  g504(.A(G43gat), .B1(new_n687), .B2(new_n486), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n695), .A2(new_n506), .A3(new_n485), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(KEYINPUT47), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n661), .ZN(new_n709));
  OAI21_X1  g508(.A(G43gat), .B1(new_n687), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(new_n707), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n708), .B1(new_n711), .B2(KEYINPUT47), .ZN(G1330gat));
  AND3_X1   g511(.A1(new_n695), .A2(new_n519), .A3(new_n427), .ZN(new_n713));
  INV_X1    g512(.A(new_n519), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n499), .A2(KEYINPUT44), .A3(new_n682), .ZN(new_n715));
  INV_X1    g514(.A(new_n643), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n677), .B1(new_n676), .B2(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n427), .B(new_n686), .C1(new_n715), .C2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n713), .B1(new_n714), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT48), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT112), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n718), .A2(new_n721), .A3(new_n714), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n718), .B2(new_n714), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n722), .A2(new_n723), .A3(new_n713), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n725));
  OAI21_X1  g524(.A(new_n720), .B1(new_n724), .B2(new_n725), .ZN(G1331gat));
  INV_X1    g525(.A(new_n553), .ZN(new_n727));
  INV_X1    g526(.A(new_n644), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n676), .A2(new_n727), .A3(new_n608), .A4(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n688), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT97), .B(G57gat), .Z(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1332gat));
  NOR2_X1   g531(.A1(new_n281), .A2(new_n609), .ZN(new_n733));
  AND4_X1   g532(.A1(new_n727), .A2(new_n676), .A3(new_n728), .A4(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  AND2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n734), .B2(new_n735), .ZN(G1333gat));
  INV_X1    g537(.A(new_n485), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n729), .A2(KEYINPUT113), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT113), .B1(new_n729), .B2(new_n739), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(new_n554), .A3(new_n741), .ZN(new_n742));
  OR3_X1    g541(.A1(new_n729), .A2(new_n554), .A3(new_n709), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1334gat));
  NOR2_X1   g545(.A1(new_n729), .A2(new_n426), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT115), .B(G78gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1335gat));
  AOI211_X1 g548(.A(new_n553), .B(new_n625), .C1(new_n667), .C2(new_n684), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n608), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n751), .A2(new_n283), .A3(new_n688), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n625), .A2(new_n553), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n694), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(KEYINPUT116), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n609), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n756), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(KEYINPUT116), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n694), .A2(new_n758), .A3(new_n753), .A4(new_n759), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(G85gat), .B1(new_n761), .B2(new_n646), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n752), .A2(new_n762), .ZN(G1336gat));
  INV_X1    g562(.A(KEYINPUT117), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n685), .A2(new_n608), .A3(new_n280), .A4(new_n753), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G92gat), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n757), .A2(new_n571), .A3(new_n280), .A4(new_n760), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n764), .B(KEYINPUT52), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n764), .A2(KEYINPUT52), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n764), .A2(KEYINPUT52), .ZN(new_n770));
  AND4_X1   g569(.A1(new_n769), .A2(new_n766), .A3(new_n770), .A4(new_n767), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n768), .A2(new_n771), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n751), .B2(new_n709), .ZN(new_n773));
  INV_X1    g572(.A(G99gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n761), .A2(new_n774), .A3(new_n485), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n757), .A2(new_n427), .A3(new_n760), .ZN(new_n777));
  INV_X1    g576(.A(G106gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n750), .A2(G106gat), .A3(new_n608), .A4(new_n427), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n780), .A3(KEYINPUT53), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1339gat));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n602), .B2(new_n605), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n586), .A2(new_n604), .A3(new_n591), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n594), .A2(KEYINPUT54), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n600), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n600), .A4(new_n789), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n601), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n551), .B2(new_n552), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n535), .B1(new_n533), .B2(new_n534), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n539), .A2(new_n540), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n548), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n552), .A2(new_n608), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n682), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n552), .A2(new_n798), .ZN(new_n801));
  INV_X1    g600(.A(new_n794), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n679), .A2(new_n801), .A3(new_n681), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n625), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n644), .A2(new_n553), .A3(new_n608), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n806), .A2(new_n688), .A3(new_n280), .ZN(new_n807));
  INV_X1    g606(.A(new_n487), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n727), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(new_n318), .ZN(G1340gat));
  NOR2_X1   g610(.A1(new_n809), .A2(new_n609), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(new_n316), .ZN(G1341gat));
  INV_X1    g612(.A(new_n625), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(KEYINPUT118), .B(G127gat), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n815), .B(new_n816), .ZN(G1342gat));
  NOR2_X1   g616(.A1(new_n809), .A2(new_n643), .ZN(new_n818));
  INV_X1    g617(.A(G134gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT56), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n821), .B(new_n823), .C1(new_n819), .C2(new_n818), .ZN(G1343gat));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825));
  INV_X1    g624(.A(new_n799), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n825), .B(new_n826), .C1(new_n727), .C2(new_n794), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT119), .B1(new_n795), .B2(new_n799), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n643), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n625), .B1(new_n829), .B2(new_n803), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n427), .B1(new_n830), .B2(new_n805), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT57), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n833), .B(new_n427), .C1(new_n804), .C2(new_n805), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n673), .A2(new_n688), .A3(new_n280), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n832), .A2(new_n553), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G141gat), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n661), .A2(new_n426), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n553), .A2(new_n296), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT120), .Z(new_n842));
  AND3_X1   g641(.A1(new_n807), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n839), .A2(KEYINPUT121), .A3(KEYINPUT58), .A4(new_n844), .ZN(new_n845));
  OR2_X1    g644(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n846));
  NAND2_X1  g645(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n836), .B1(new_n831), .B2(KEYINPUT57), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n296), .B1(new_n848), .B2(new_n553), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n846), .B(new_n847), .C1(new_n849), .C2(new_n843), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n845), .A2(new_n850), .ZN(G1344gat));
  NAND2_X1  g650(.A1(new_n807), .A2(new_n840), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n342), .A2(new_n297), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n855), .A3(new_n608), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n716), .A2(new_n802), .A3(new_n801), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n625), .B1(new_n829), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n833), .B(new_n427), .C1(new_n859), .C2(new_n805), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT57), .B1(new_n806), .B2(new_n426), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n860), .A2(new_n608), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n835), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n857), .B1(new_n863), .B2(G148gat), .ZN(new_n864));
  AOI211_X1 g663(.A(KEYINPUT59), .B(new_n855), .C1(new_n848), .C2(new_n608), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n856), .B1(new_n864), .B2(new_n865), .ZN(G1345gat));
  AOI21_X1  g665(.A(G155gat), .B1(new_n853), .B2(new_n625), .ZN(new_n867));
  INV_X1    g666(.A(new_n848), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n814), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n867), .B1(new_n869), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g669(.A(G162gat), .B1(new_n853), .B2(new_n716), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n868), .A2(new_n292), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n683), .ZN(G1347gat));
  OAI211_X1 g672(.A(new_n688), .B(new_n808), .C1(new_n804), .C2(new_n805), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n281), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n553), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(G169gat), .ZN(G1348gat));
  NOR2_X1   g676(.A1(new_n806), .A2(new_n646), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n808), .A3(new_n733), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(G176gat), .ZN(G1349gat));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n875), .A2(new_n625), .ZN(new_n882));
  NAND2_X1  g681(.A1(KEYINPUT122), .A2(G183gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n209), .A2(new_n211), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n613), .A2(KEYINPUT122), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n875), .A2(new_n625), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n881), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(KEYINPUT60), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n884), .A2(new_n888), .ZN(new_n893));
  INV_X1    g692(.A(new_n890), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(KEYINPUT124), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n875), .A2(new_n203), .A3(new_n683), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n875), .A2(new_n716), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(G190gat), .ZN(new_n900));
  AOI211_X1 g699(.A(KEYINPUT61), .B(new_n203), .C1(new_n875), .C2(new_n716), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT125), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n897), .B(new_n904), .C1(new_n900), .C2(new_n901), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1351gat));
  NOR3_X1   g705(.A1(new_n661), .A2(new_n646), .A3(new_n281), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n860), .A2(new_n861), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G197gat), .B1(new_n908), .B2(new_n727), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n806), .A2(new_n426), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n907), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n910), .A2(new_n907), .A3(KEYINPUT126), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(G197gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n909), .B1(new_n916), .B2(new_n727), .ZN(G1352gat));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT127), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n878), .B1(KEYINPUT127), .B2(new_n918), .ZN(new_n920));
  INV_X1    g719(.A(G204gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n840), .A2(new_n921), .A3(new_n733), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OR3_X1    g722(.A1(new_n920), .A2(new_n919), .A3(new_n922), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n862), .A2(new_n907), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n923), .B(new_n924), .C1(new_n925), .C2(new_n921), .ZN(G1353gat));
  NAND4_X1  g725(.A1(new_n860), .A2(new_n625), .A3(new_n861), .A4(new_n907), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n927), .B2(G211gat), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n625), .A2(new_n254), .ZN(new_n930));
  OAI22_X1  g729(.A1(new_n928), .A2(new_n929), .B1(new_n915), .B2(new_n930), .ZN(G1354gat));
  AOI21_X1  g730(.A(new_n682), .B1(new_n913), .B2(new_n914), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n716), .A2(G218gat), .ZN(new_n933));
  OAI22_X1  g732(.A1(new_n932), .A2(G218gat), .B1(new_n908), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(G1355gat));
endmodule


