//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT64), .B1(new_n191), .B2(G143), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(new_n189), .A3(G146), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G128), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n191), .A2(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n189), .A2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n195), .A2(new_n198), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n195), .A2(new_n207), .B1(new_n209), .B2(new_n203), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n206), .B1(new_n205), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G224), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G953), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n211), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G110), .B(G122), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G104), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT81), .A2(G107), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT81), .A2(G107), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT3), .B1(new_n222), .B2(G107), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(G107), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(KEYINPUT81), .A2(G107), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT81), .A2(G107), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n227), .A2(new_n217), .A3(G104), .A4(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G101), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n229), .A2(new_n230), .A3(new_n223), .A4(new_n224), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n226), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G116), .B(G119), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n235), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n233), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n240), .B(G101), .C1(new_n221), .C2(new_n225), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n232), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(G104), .B1(new_n227), .B2(new_n228), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n222), .A2(G107), .ZN(new_n244));
  OAI21_X1  g058(.A(G101), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n233), .A2(KEYINPUT5), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT5), .ZN(new_n247));
  INV_X1    g061(.A(G119), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G116), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n249), .A2(G113), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n231), .A2(new_n245), .A3(new_n251), .A4(new_n238), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n216), .B1(new_n242), .B2(new_n252), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT85), .B(KEYINPUT6), .Z(new_n254));
  AND2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT84), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n242), .A2(new_n216), .A3(new_n252), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT6), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n256), .B1(new_n258), .B2(new_n253), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n242), .A2(new_n252), .ZN(new_n260));
  INV_X1    g074(.A(new_n216), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n262), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n257), .ZN(new_n263));
  AOI211_X1 g077(.A(new_n215), .B(new_n255), .C1(new_n259), .C2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  INV_X1    g079(.A(new_n211), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT88), .B1(new_n210), .B2(new_n205), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT7), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(new_n213), .ZN(new_n269));
  OR2_X1    g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n266), .A2(new_n269), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(new_n257), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n216), .B(KEYINPUT8), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n250), .A2(KEYINPUT86), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n249), .A2(G113), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT86), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(new_n246), .A3(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n279), .A2(new_n238), .A3(new_n231), .A4(new_n245), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n245), .A2(new_n231), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n251), .A2(new_n238), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n281), .A2(KEYINPUT87), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT87), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n274), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n265), .B1(new_n272), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n188), .B1(new_n264), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n259), .A2(new_n263), .ZN(new_n290));
  INV_X1    g104(.A(new_n215), .ZN(new_n291));
  INV_X1    g105(.A(new_n255), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n270), .A2(new_n271), .A3(new_n257), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n284), .A2(new_n286), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n273), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n293), .A2(new_n297), .A3(new_n187), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G214), .B1(G237), .B2(G902), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT89), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT89), .ZN(new_n302));
  INV_X1    g116(.A(new_n300), .ZN(new_n303));
  AOI211_X1 g117(.A(new_n302), .B(new_n303), .C1(new_n289), .C2(new_n298), .ZN(new_n304));
  INV_X1    g118(.A(G128), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n305), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n195), .A2(new_n306), .ZN(new_n307));
  AOI211_X1 g121(.A(new_n197), .B(new_n190), .C1(new_n192), .C2(new_n194), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n231), .B(new_n245), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT10), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n232), .A2(new_n210), .A3(new_n241), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT11), .ZN(new_n313));
  INV_X1    g127(.A(G134), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(G137), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(G137), .ZN(new_n316));
  INV_X1    g130(.A(G137), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT11), .A3(G134), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G131), .ZN(new_n320));
  INV_X1    g134(.A(G131), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n315), .A2(new_n318), .A3(new_n321), .A4(new_n316), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n193), .B1(new_n189), .B2(G146), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n191), .A2(KEYINPUT64), .A3(G143), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n201), .B(new_n198), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n200), .A2(new_n203), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n329), .A2(KEYINPUT10), .A3(new_n231), .A4(new_n245), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n311), .A2(new_n312), .A3(new_n324), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n282), .A2(new_n204), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n309), .ZN(new_n333));
  NOR2_X1   g147(.A1(KEYINPUT82), .A2(KEYINPUT12), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n323), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n324), .B1(new_n332), .B2(new_n309), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n331), .B(new_n335), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  XOR2_X1   g153(.A(G110), .B(G140), .Z(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT80), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT69), .B(G953), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n342), .A2(G227), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n341), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT83), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n338), .B1(new_n333), .B2(new_n323), .ZN(new_n347));
  INV_X1    g161(.A(new_n334), .ZN(new_n348));
  AOI211_X1 g162(.A(new_n324), .B(new_n348), .C1(new_n332), .C2(new_n309), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n344), .A4(new_n331), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n311), .A2(new_n312), .A3(new_n330), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n323), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n331), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n345), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n346), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G469), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n265), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n339), .A2(new_n345), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n354), .A2(new_n344), .A3(new_n331), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(G469), .A3(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n358), .A2(new_n265), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n359), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT9), .B(G234), .ZN(new_n367));
  OAI21_X1  g181(.A(G221), .B1(new_n367), .B2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n301), .A2(new_n304), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n371));
  XNOR2_X1  g185(.A(G113), .B(G122), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(new_n222), .ZN(new_n373));
  INV_X1    g187(.A(G237), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT68), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT68), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G237), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n342), .A3(G214), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n189), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n378), .A2(new_n342), .A3(G143), .A4(G214), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g196(.A1(KEYINPUT18), .A2(G131), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(G125), .B(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n191), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G140), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n388), .A2(KEYINPUT73), .A3(G125), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n385), .B2(KEYINPUT73), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n387), .B1(new_n390), .B2(G146), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n382), .A2(KEYINPUT17), .A3(G131), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT91), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n321), .B1(new_n380), .B2(new_n381), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT91), .A3(KEYINPUT17), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n380), .A2(new_n321), .A3(new_n381), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(new_n396), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT17), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n395), .A2(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT16), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(new_n388), .A3(G125), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n205), .A2(G140), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n388), .A2(G125), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT73), .ZN(new_n406));
  OR3_X1    g220(.A1(new_n388), .A2(KEYINPUT73), .A3(G125), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n402), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT74), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n403), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n390), .A2(KEYINPUT74), .A3(new_n402), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n191), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT74), .B1(new_n390), .B2(new_n402), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n409), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n413), .A2(new_n414), .A3(G146), .A4(new_n403), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(KEYINPUT75), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT75), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n417), .B(new_n191), .C1(new_n410), .C2(new_n411), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n392), .B1(new_n401), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n373), .B1(new_n420), .B2(KEYINPUT92), .ZN(new_n421));
  INV_X1    g235(.A(new_n392), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n416), .A2(new_n418), .ZN(new_n423));
  INV_X1    g237(.A(new_n397), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT91), .B1(new_n396), .B2(KEYINPUT17), .ZN(new_n425));
  INV_X1    g239(.A(new_n396), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n380), .A2(new_n321), .A3(new_n381), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI22_X1  g242(.A1(new_n424), .A2(new_n425), .B1(new_n428), .B2(KEYINPUT17), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n422), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT92), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n373), .B(KEYINPUT90), .Z(new_n433));
  AOI22_X1  g247(.A1(new_n421), .A2(new_n432), .B1(new_n420), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n371), .B1(new_n434), .B2(G902), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n420), .A2(new_n433), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n422), .B(KEYINPUT92), .C1(new_n423), .C2(new_n429), .ZN(new_n437));
  INV_X1    g251(.A(new_n373), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n420), .A2(KEYINPUT92), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT93), .A3(new_n265), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n435), .A2(new_n442), .A3(G475), .ZN(new_n443));
  MUX2_X1   g257(.A(new_n385), .B(new_n390), .S(KEYINPUT19), .Z(new_n444));
  OAI211_X1 g258(.A(new_n428), .B(new_n415), .C1(G146), .C2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n438), .B1(new_n446), .B2(new_n392), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n436), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(G475), .A2(G902), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(KEYINPUT20), .A3(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G478), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n457));
  XNOR2_X1  g271(.A(G116), .B(G122), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT94), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n227), .A2(new_n228), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G128), .B(G143), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n463), .A2(new_n314), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n314), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT14), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G116), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(KEYINPUT14), .A3(G122), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G107), .ZN(new_n470));
  OAI22_X1  g284(.A1(new_n464), .A2(new_n465), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  OR3_X1    g285(.A1(new_n462), .A2(new_n471), .A3(KEYINPUT96), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT96), .B1(new_n462), .B2(new_n471), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n475), .A2(new_n305), .A3(G143), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n314), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n463), .A2(new_n475), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n464), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n460), .A2(new_n461), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n462), .ZN(new_n481));
  INV_X1    g295(.A(G217), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n367), .A2(new_n482), .A3(G953), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n474), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n474), .B2(new_n481), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n457), .B1(new_n486), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n485), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n474), .A2(new_n481), .A3(new_n483), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n457), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n265), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G953), .ZN(new_n494));
  INV_X1    g308(.A(G952), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n495), .A2(KEYINPUT97), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(KEYINPUT97), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(G234), .B2(G237), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n265), .B(new_n342), .C1(G234), .C2(G237), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT21), .B(G898), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n443), .A2(new_n455), .A3(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n370), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT23), .B1(new_n305), .B2(G119), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT72), .B1(new_n248), .B2(G128), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G110), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g324(.A(G119), .B(G128), .Z(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT24), .B(G110), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n416), .A2(new_n418), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n508), .A2(new_n509), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n511), .A2(new_n512), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n415), .B(new_n386), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(G221), .A2(G234), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n342), .A2(KEYINPUT76), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT76), .B1(new_n342), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT22), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n523), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT22), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n521), .ZN(new_n527));
  AOI21_X1  g341(.A(G137), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n527), .A3(G137), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(KEYINPUT77), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT77), .ZN(new_n532));
  INV_X1    g346(.A(new_n530), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n532), .B1(new_n533), .B2(new_n528), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n519), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n515), .A2(new_n530), .A3(new_n529), .A4(new_n518), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n265), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n539), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n536), .A2(new_n265), .A3(new_n537), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n482), .B1(G234), .B2(new_n265), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n536), .A2(new_n537), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT79), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n536), .A2(KEYINPUT79), .A3(new_n537), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n545), .A2(G902), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT32), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n323), .A2(new_n210), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n314), .A2(G137), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n317), .A2(G134), .ZN(new_n558));
  OAI21_X1  g372(.A(G131), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n322), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n329), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT30), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n322), .A2(new_n559), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT65), .B1(new_n204), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT65), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n329), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n564), .A2(new_n566), .A3(KEYINPUT30), .A4(new_n556), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT66), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n563), .B1(new_n327), .B2(new_n328), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n570), .A2(new_n565), .B1(new_n323), .B2(new_n210), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n571), .A2(KEYINPUT66), .A3(KEYINPUT30), .A4(new_n564), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n569), .A2(new_n239), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n378), .A2(new_n342), .A3(G210), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT27), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT26), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT27), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n378), .A2(new_n342), .A3(new_n577), .A4(G210), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n576), .B1(new_n575), .B2(new_n578), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n230), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n575), .A2(new_n578), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT26), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(G101), .A3(new_n584), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n239), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n564), .A2(new_n566), .A3(new_n587), .A4(new_n556), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT67), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n586), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n555), .B1(new_n573), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n581), .A2(new_n585), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n571), .A2(KEYINPUT67), .A3(new_n587), .A4(new_n564), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n588), .A2(new_n589), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n569), .A2(new_n239), .A3(new_n572), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT31), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(KEYINPUT28), .A3(new_n596), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n587), .B1(new_n556), .B2(new_n561), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT28), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n556), .A2(new_n561), .A3(new_n587), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n593), .A2(new_n599), .B1(new_n594), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(G472), .A2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n554), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n594), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT31), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT31), .B1(new_n597), .B2(new_n598), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(KEYINPUT32), .A3(new_n607), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n603), .A2(new_n602), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT70), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT29), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n594), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n571), .A2(new_n564), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n595), .A2(new_n596), .B1(new_n620), .B2(new_n239), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n617), .B(new_n619), .C1(new_n621), .C2(new_n602), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT71), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n620), .A2(new_n239), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n590), .B2(new_n591), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT28), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n627), .A2(KEYINPUT71), .A3(new_n617), .A4(new_n619), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n600), .A2(new_n586), .A3(new_n604), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n618), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n595), .A2(new_n596), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n586), .B1(new_n598), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n265), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n629), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n553), .B1(new_n615), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n505), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  INV_X1    g452(.A(new_n368), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n359), .B2(new_n365), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n546), .A2(new_n640), .A3(new_n552), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n642), .B(G472), .C1(new_n606), .C2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n613), .A2(new_n607), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n613), .A2(new_n265), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n642), .B1(new_n646), .B2(G472), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n641), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(G478), .B1(new_n490), .B2(new_n265), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n474), .A2(new_n481), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT33), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n650), .B(new_n652), .C1(new_n486), .C2(KEYINPUT99), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n650), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n490), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n456), .A2(G902), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n649), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n443), .B2(new_n455), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n502), .B(new_n303), .C1(new_n289), .C2(new_n298), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n648), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT100), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT34), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G104), .ZN(G6));
  AND4_X1   g479(.A1(new_n443), .A2(new_n661), .A3(new_n455), .A4(new_n493), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n648), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT101), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT35), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G107), .ZN(G9));
  AND2_X1   g484(.A1(new_n531), .A2(new_n534), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT36), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n671), .A2(new_n672), .A3(new_n515), .A4(new_n518), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n519), .B1(new_n535), .B2(KEYINPUT36), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n673), .A2(new_n551), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n544), .B2(new_n545), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n645), .A2(new_n676), .A3(new_n647), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n505), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  NAND2_X1  g494(.A1(new_n443), .A2(new_n455), .ZN(new_n681));
  INV_X1    g495(.A(new_n493), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n499), .B1(new_n500), .B2(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n635), .A2(new_n609), .A3(new_n614), .ZN(new_n686));
  INV_X1    g500(.A(new_n675), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n546), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n303), .B1(new_n289), .B2(new_n298), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n688), .A3(new_n689), .A4(new_n640), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n685), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(G475), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n421), .A2(new_n432), .ZN(new_n695));
  AOI21_X1  g509(.A(G902), .B1(new_n695), .B2(new_n436), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n694), .B1(new_n696), .B2(KEYINPUT93), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n454), .B1(new_n697), .B2(new_n435), .ZN(new_n698));
  INV_X1    g512(.A(new_n684), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n493), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT102), .B1(new_n700), .B2(new_n690), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  XOR2_X1   g517(.A(new_n684), .B(KEYINPUT39), .Z(new_n704));
  NAND2_X1  g518(.A1(new_n640), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n705), .B(KEYINPUT40), .Z(new_n706));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n707));
  AOI211_X1 g521(.A(new_n698), .B(new_n682), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n594), .A2(new_n626), .B1(new_n597), .B2(new_n598), .ZN(new_n709));
  OAI21_X1  g523(.A(G472), .B1(new_n709), .B2(G902), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n615), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n264), .A2(new_n188), .A3(new_n288), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n187), .B1(new_n293), .B2(new_n297), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT38), .ZN(new_n716));
  NOR4_X1   g530(.A1(new_n712), .A2(new_n716), .A3(new_n303), .A4(new_n688), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n708), .B(new_n717), .C1(new_n707), .C2(new_n706), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G143), .ZN(G45));
  AOI211_X1 g533(.A(new_n684), .B(new_n659), .C1(new_n443), .C2(new_n455), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n691), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G146), .ZN(G48));
  AND2_X1   g536(.A1(new_n549), .A2(new_n550), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n723), .A2(new_n551), .B1(new_n544), .B2(new_n545), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n357), .A2(new_n358), .A3(new_n265), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n358), .B1(new_n357), .B2(new_n265), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n725), .A2(new_n726), .A3(new_n639), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n686), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n660), .A3(new_n661), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND2_X1  g545(.A1(new_n666), .A2(new_n728), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT104), .B(G116), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G18));
  AND3_X1   g548(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n443), .A2(new_n455), .A3(new_n727), .A4(new_n503), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  AOI21_X1  g552(.A(new_n682), .B1(new_n443), .B2(new_n455), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n646), .A2(G472), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n611), .A2(new_n612), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n586), .B1(new_n627), .B2(new_n617), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n607), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n553), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n502), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n727), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n739), .A2(new_n745), .A3(new_n747), .A4(new_n689), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  INV_X1    g563(.A(new_n727), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n299), .A2(new_n300), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n744), .A2(new_n676), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n720), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  NAND3_X1  g570(.A1(new_n289), .A2(new_n300), .A3(new_n298), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n686), .A2(new_n724), .A3(new_n640), .A4(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n720), .A2(new_n759), .A3(KEYINPUT42), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT42), .B1(new_n720), .B2(new_n759), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n321), .ZN(G33));
  NAND2_X1  g577(.A1(new_n685), .A2(new_n759), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  XOR2_X1   g579(.A(new_n757), .B(KEYINPUT107), .Z(new_n766));
  NAND3_X1  g580(.A1(new_n360), .A2(KEYINPUT45), .A3(new_n361), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(G469), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT45), .B1(new_n360), .B2(new_n361), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n364), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT105), .A3(new_n359), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n771), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT105), .B1(new_n772), .B2(new_n359), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(new_n368), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n704), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n681), .A2(new_n659), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT43), .B1(new_n681), .B2(new_n659), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n688), .B1(new_n645), .B2(new_n647), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT106), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n766), .B(new_n779), .C1(new_n780), .C2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n780), .B2(new_n788), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  NAND2_X1  g605(.A1(new_n777), .A2(new_n368), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT47), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n777), .A2(new_n794), .A3(new_n368), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n686), .A2(new_n724), .A3(new_n757), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n793), .A2(new_n720), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  NOR2_X1   g612(.A1(new_n750), .A2(new_n757), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n712), .A2(new_n724), .A3(new_n799), .A4(new_n499), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n698), .A3(new_n659), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n785), .A2(KEYINPUT112), .A3(new_n499), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n783), .A2(new_n499), .A3(new_n784), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n750), .B(new_n757), .C1(new_n804), .C2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n803), .B1(new_n808), .B2(new_n753), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n793), .A2(new_n795), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n725), .A2(new_n726), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n639), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n766), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n814));
  INV_X1    g628(.A(new_n745), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n804), .B2(new_n807), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n716), .A2(new_n303), .A3(new_n727), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT114), .Z(new_n819));
  AND3_X1   g633(.A1(new_n816), .A2(KEYINPUT50), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT50), .B1(new_n816), .B2(new_n819), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n809), .B(new_n817), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n808), .A2(new_n636), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT48), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT48), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n808), .A2(new_n827), .A3(new_n636), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n816), .A2(new_n752), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n498), .B1(new_n801), .B2(new_n660), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n813), .A2(new_n816), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n814), .A2(new_n823), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n809), .B1(new_n820), .B2(new_n821), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(new_n837), .B2(KEYINPUT51), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT115), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n838), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n829), .A2(new_n832), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n824), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n729), .A2(new_n732), .A3(new_n737), .A4(new_n748), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n301), .A2(new_n304), .A3(new_n502), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n443), .A2(new_n455), .A3(new_n493), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n648), .B(new_n846), .C1(new_n847), .C2(new_n660), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n370), .B(new_n504), .C1(new_n636), .C2(new_n677), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n760), .A2(new_n761), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n744), .A2(new_n369), .A3(new_n757), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n660), .A3(new_n699), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n369), .A2(new_n757), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n487), .A2(new_n492), .A3(new_n699), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n698), .A2(new_n686), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n676), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n759), .A2(new_n847), .A3(new_n699), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT108), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT108), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n635), .A2(new_n609), .A3(new_n614), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n715), .A2(new_n640), .A3(new_n300), .A4(new_n856), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n720), .A2(new_n853), .B1(new_n864), .B2(new_n698), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n861), .B(new_n764), .C1(new_n865), .C2(new_n676), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n851), .A2(new_n852), .A3(new_n860), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT109), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n682), .B(new_n751), .C1(new_n443), .C2(new_n455), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n727), .A2(new_n746), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n553), .A3(new_n744), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n869), .A2(new_n871), .B1(new_n735), .B2(new_n736), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n728), .B(new_n661), .C1(new_n847), .C2(new_n660), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n873), .A3(new_n848), .A4(new_n849), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n762), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT109), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n860), .A4(new_n866), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n720), .B1(new_n754), .B2(new_n691), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n676), .A2(new_n640), .A3(new_n699), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT110), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n711), .A3(new_n869), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n702), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n702), .A2(new_n878), .A3(new_n881), .A4(KEYINPUT52), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n868), .A2(new_n877), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(KEYINPUT53), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n890), .A2(new_n867), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n867), .A2(KEYINPUT109), .B1(new_n884), .B2(new_n885), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(KEYINPUT53), .A3(new_n877), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n892), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT111), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI211_X1 g712(.A(KEYINPUT111), .B(new_n892), .C1(new_n889), .C2(new_n895), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI22_X1  g714(.A1(new_n844), .A2(new_n900), .B1(G952), .B2(G953), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n811), .B(KEYINPUT49), .Z(new_n902));
  NOR4_X1   g716(.A1(new_n902), .A2(new_n553), .A3(new_n303), .A4(new_n639), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(new_n712), .A3(new_n716), .A4(new_n781), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n904), .ZN(G75));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(KEYINPUT56), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n889), .A2(new_n891), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(G902), .ZN(new_n909));
  INV_X1    g723(.A(G210), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n290), .A2(new_n292), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n291), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT55), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n914), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n907), .B(new_n916), .C1(new_n909), .C2(new_n910), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n342), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n915), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT117), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT117), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n915), .A2(new_n922), .A3(new_n917), .A4(new_n919), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(G51));
  NAND2_X1  g738(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n893), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n363), .B(KEYINPUT57), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n357), .ZN(new_n929));
  OR3_X1    g743(.A1(new_n909), .A2(new_n769), .A3(new_n768), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n918), .B1(new_n929), .B2(new_n930), .ZN(G54));
  AOI21_X1  g745(.A(new_n265), .B1(new_n889), .B2(new_n891), .ZN(new_n932));
  NAND2_X1  g746(.A1(KEYINPUT58), .A2(G475), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT118), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n436), .A3(new_n447), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n932), .A2(new_n448), .A3(new_n934), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n919), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G60));
  NAND2_X1  g754(.A1(G478), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT59), .Z(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n898), .B2(new_n899), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT120), .ZN(new_n945));
  INV_X1    g759(.A(new_n657), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n945), .B1(new_n944), .B2(new_n946), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n926), .A2(new_n657), .A3(new_n943), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n919), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(G63));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT60), .Z(new_n953));
  NAND4_X1  g767(.A1(new_n908), .A2(new_n673), .A3(new_n674), .A4(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n908), .A2(new_n953), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n919), .B(new_n954), .C1(new_n955), .C2(new_n723), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(KEYINPUT121), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(KEYINPUT121), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G66));
  OAI21_X1  g775(.A(G953), .B1(new_n501), .B2(new_n212), .ZN(new_n962));
  INV_X1    g776(.A(new_n342), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n962), .B1(new_n851), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n912), .B1(G898), .B2(new_n342), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT122), .Z(new_n966));
  XNOR2_X1  g780(.A(new_n964), .B(new_n966), .ZN(G69));
  NAND2_X1  g781(.A1(new_n569), .A2(new_n572), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT123), .Z(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(new_n444), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n702), .A2(new_n878), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n718), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n847), .A2(new_n660), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n977), .A2(new_n704), .A3(new_n759), .A4(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n797), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n790), .A2(new_n974), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT124), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n971), .B1(new_n984), .B2(new_n963), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n963), .A2(G900), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n778), .A2(new_n636), .A3(new_n704), .A4(new_n869), .ZN(new_n987));
  AND4_X1   g801(.A1(new_n852), .A2(new_n797), .A3(new_n764), .A4(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n790), .A2(new_n972), .A3(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n970), .B(new_n986), .C1(new_n989), .C2(new_n963), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n342), .B1(G227), .B2(G900), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n990), .B2(KEYINPUT126), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n991), .B(new_n993), .Z(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n989), .B2(new_n874), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n598), .A2(new_n632), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT127), .Z(new_n999));
  NOR2_X1   g813(.A1(new_n999), .A2(new_n586), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n918), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n996), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n984), .B2(new_n851), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n999), .A2(new_n586), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n633), .B1(new_n598), .B2(new_n597), .ZN(new_n1006));
  AOI211_X1 g820(.A(new_n1006), .B(new_n1002), .C1(new_n889), .C2(new_n895), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1005), .A2(new_n1007), .ZN(G57));
endmodule


