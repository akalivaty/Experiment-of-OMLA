//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  AND2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT65), .B(G20), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n202), .A2(new_n203), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(new_n215), .A2(KEYINPUT0), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G226), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n224), .B1(new_n201), .B2(new_n225), .C1(new_n203), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n212), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n216), .A2(new_n223), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT69), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n250), .A2(new_n251), .B1(G1), .B2(G13), .ZN(new_n252));
  NAND4_X1  g0052(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n217), .A2(G33), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT15), .B(G87), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n206), .A2(new_n217), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n254), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT72), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT72), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n264), .B(new_n254), .C1(new_n257), .C2(new_n261), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G13), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G20), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n252), .A2(new_n269), .A3(new_n253), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n206), .B1(new_n209), .B2(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n269), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n271), .A2(new_n272), .B1(new_n206), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G107), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n218), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G232), .A2(G1698), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n226), .B2(G1698), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n280), .B(new_n284), .C1(new_n278), .C2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  INV_X1    g0088(.A(G45), .ZN(new_n289));
  AOI21_X1  g0089(.A(G1), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT67), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n218), .B1(new_n291), .B2(new_n282), .ZN(new_n292));
  NAND3_X1  g0092(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G244), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n290), .A2(KEYINPUT66), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n282), .A2(new_n291), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(new_n281), .A3(new_n293), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT66), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n296), .A2(new_n298), .A3(G274), .A4(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n287), .A2(new_n295), .A3(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(G179), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n275), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n270), .A2(KEYINPUT70), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT70), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n252), .A2(new_n269), .A3(new_n310), .A4(new_n253), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n258), .B1(new_n209), .B2(G20), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n312), .A2(new_n313), .B1(new_n273), .B2(new_n258), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT3), .B(G33), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT7), .B1(new_n315), .B2(G20), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT7), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n278), .A2(new_n217), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n318), .A3(G68), .ZN(new_n319));
  INV_X1    g0119(.A(G159), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT78), .B1(new_n260), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT78), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n259), .A2(new_n322), .A3(G159), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G58), .A2(G68), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT77), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(KEYINPUT77), .A2(G58), .A3(G68), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n220), .A3(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n321), .A2(new_n323), .B1(new_n328), .B2(G20), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n319), .A2(new_n329), .A3(KEYINPUT16), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n254), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n278), .A2(new_n317), .A3(new_n210), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n210), .A2(KEYINPUT65), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT65), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(new_n315), .ZN(new_n337));
  OAI211_X1 g0137(.A(G68), .B(new_n332), .C1(new_n337), .C2(new_n317), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT16), .B1(new_n338), .B2(new_n329), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n314), .B1(new_n331), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n294), .A2(G232), .ZN(new_n341));
  INV_X1    g0141(.A(G33), .ZN(new_n342));
  INV_X1    g0142(.A(G87), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(G223), .A2(G1698), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n225), .B2(G1698), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n344), .B1(new_n346), .B2(new_n315), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n341), .B(new_n302), .C1(new_n283), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G169), .ZN(new_n349));
  INV_X1    g0149(.A(G179), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n348), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n340), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT18), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT18), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n340), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n348), .A2(G200), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n347), .A2(new_n283), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n357), .A2(G190), .A3(new_n302), .A4(new_n341), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n339), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(new_n254), .A3(new_n330), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n359), .A2(new_n361), .A3(KEYINPUT17), .A4(new_n314), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT17), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n356), .A2(new_n358), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n340), .B2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n353), .A2(new_n355), .A3(new_n362), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n303), .A2(G200), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n266), .A2(new_n274), .A3(new_n367), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n368), .A2(KEYINPUT73), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n287), .A2(new_n295), .A3(G190), .A4(new_n302), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT71), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n368), .B2(KEYINPUT73), .ZN(new_n372));
  AOI211_X1 g0172(.A(new_n308), .B(new_n366), .C1(new_n369), .C2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT10), .ZN(new_n374));
  INV_X1    g0174(.A(G1698), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n315), .A2(G222), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT68), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n376), .B(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n278), .A2(new_n375), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n379), .A2(G223), .B1(G77), .B2(new_n278), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n283), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n298), .A2(new_n299), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n302), .B1(new_n225), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G190), .ZN(new_n385));
  OAI21_X1  g0185(.A(G200), .B1(new_n381), .B2(new_n383), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(KEYINPUT74), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n259), .A2(G150), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n388), .B1(new_n255), .B2(new_n258), .C1(new_n205), .C2(new_n210), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(new_n254), .B1(new_n201), .B2(new_n273), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n209), .A2(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n312), .A2(G50), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT9), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n385), .A2(new_n386), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n374), .B(new_n387), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n393), .B(KEYINPUT9), .ZN(new_n398));
  INV_X1    g0198(.A(new_n396), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(KEYINPUT74), .C2(KEYINPUT10), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  MUX2_X1   g0201(.A(G226), .B(G232), .S(G1698), .Z(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(new_n315), .B1(G33), .B2(G97), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n403), .A2(new_n283), .B1(new_n382), .B2(new_n226), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n302), .A2(KEYINPUT75), .ZN(new_n405));
  INV_X1    g0205(.A(G274), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n292), .B2(new_n293), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT75), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(new_n301), .A4(new_n296), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n404), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT13), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT76), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n405), .A2(new_n409), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n402), .A2(new_n315), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G97), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(new_n284), .B1(new_n294), .B2(G238), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n411), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT76), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n410), .A2(new_n411), .ZN(new_n421));
  AND4_X1   g0221(.A1(G190), .A2(new_n412), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n413), .A2(new_n411), .A3(new_n417), .ZN(new_n423));
  OAI21_X1  g0223(.A(G200), .B1(new_n423), .B2(new_n418), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n273), .A2(new_n203), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n425), .B(KEYINPUT12), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n255), .B2(new_n206), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n254), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT11), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n271), .A2(G68), .A3(new_n391), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n429), .B2(new_n430), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n424), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n422), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n435), .ZN(new_n438));
  OAI21_X1  g0238(.A(G169), .B1(new_n423), .B2(new_n418), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT14), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n412), .A2(new_n420), .A3(G179), .A4(new_n421), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT14), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n442), .B(G169), .C1(new_n423), .C2(new_n418), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n437), .B1(new_n438), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n384), .A2(new_n350), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(new_n393), .C1(G169), .C2(new_n384), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n373), .A2(new_n401), .A3(new_n445), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n209), .A2(G33), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n252), .A2(new_n269), .A3(new_n253), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(KEYINPUT81), .A3(G116), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT81), .ZN(new_n453));
  INV_X1    g0253(.A(G116), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n273), .A2(new_n454), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT82), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n342), .A2(G97), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n458), .B1(new_n336), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n217), .A2(KEYINPUT82), .A3(new_n459), .A4(new_n460), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n252), .A2(new_n253), .B1(G20), .B2(new_n454), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n464), .A2(KEYINPUT20), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT20), .B1(new_n464), .B2(new_n465), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n456), .B(new_n457), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n289), .A2(G1), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT5), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G41), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n288), .A2(KEYINPUT5), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n298), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n209), .B(G45), .C1(new_n288), .C2(KEYINPUT5), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT80), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n288), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n474), .A2(G270), .B1(new_n407), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n315), .A2(G257), .A3(new_n375), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n315), .A2(G264), .A3(G1698), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n278), .A2(G303), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n284), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n305), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT21), .B1(new_n468), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n468), .A2(new_n486), .A3(KEYINPUT21), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT83), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n480), .A2(new_n485), .A3(G179), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n468), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(new_n468), .B2(new_n491), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n488), .B(new_n489), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n468), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n480), .A2(new_n485), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G200), .ZN(new_n499));
  INV_X1    g0299(.A(G190), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n497), .B(new_n499), .C1(new_n500), .C2(new_n498), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n210), .A2(G107), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT86), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n268), .B(new_n503), .C1(new_n504), .C2(KEYINPUT25), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(KEYINPUT25), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n507), .A2(new_n508), .B1(new_n451), .B2(G107), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n315), .A2(G257), .A3(G1698), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n315), .A2(G250), .A3(new_n375), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G294), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n284), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n474), .A2(G264), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n407), .A2(new_n479), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n514), .A2(KEYINPUT87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n514), .A2(KEYINPUT87), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n517), .A3(new_n521), .A4(new_n515), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n519), .A2(G200), .B1(new_n522), .B2(G190), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT85), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT23), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G116), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n503), .A2(new_n525), .B1(G20), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(KEYINPUT23), .A2(G107), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n336), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n333), .B(new_n335), .C1(new_n276), .C2(new_n277), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT84), .B1(new_n530), .B2(new_n343), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT22), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT84), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n315), .A2(new_n217), .A3(new_n533), .A4(G87), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n531), .B2(new_n534), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n529), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT24), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT24), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n539), .B(new_n529), .C1(new_n535), .C2(new_n536), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n524), .B1(new_n541), .B2(new_n254), .ZN(new_n542));
  INV_X1    g0342(.A(new_n254), .ZN(new_n543));
  AOI211_X1 g0343(.A(KEYINPUT85), .B(new_n543), .C1(new_n538), .C2(new_n540), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n509), .B(new_n523), .C1(new_n542), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n474), .A2(G257), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n517), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n315), .A2(G250), .A3(G1698), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n460), .ZN(new_n549));
  INV_X1    g0349(.A(G244), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(G1698), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT4), .B1(new_n315), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n315), .A2(KEYINPUT4), .A3(new_n551), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT79), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n315), .A2(KEYINPUT79), .A3(KEYINPUT4), .A4(new_n551), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n547), .B1(new_n559), .B2(new_n284), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n350), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT6), .ZN(new_n562));
  INV_X1    g0362(.A(G97), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(new_n279), .ZN(new_n564));
  NOR2_X1   g0364(.A1(G97), .A2(G107), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n279), .A2(KEYINPUT6), .A3(G97), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(new_n336), .B1(G77), .B2(new_n259), .ZN(new_n569));
  OAI211_X1 g0369(.A(G107), .B(new_n332), .C1(new_n337), .C2(new_n317), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n543), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n273), .A2(new_n563), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n450), .B2(new_n563), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n283), .B1(new_n553), .B2(new_n558), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n305), .B1(new_n575), .B2(new_n547), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n561), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(G200), .B1(new_n575), .B2(new_n547), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n571), .A2(new_n573), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n559), .A2(new_n284), .ZN(new_n580));
  INV_X1    g0380(.A(new_n547), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n578), .B(new_n579), .C1(new_n582), .C2(new_n500), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n550), .A2(G1698), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(G238), .B2(G1698), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n526), .B1(new_n586), .B2(new_n278), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n284), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n469), .A2(new_n406), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n298), .B(new_n589), .C1(G250), .C2(new_n469), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(G179), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT19), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n255), .B2(new_n563), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n565), .A2(new_n343), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n415), .A2(new_n593), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n336), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n315), .A2(new_n217), .A3(G68), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(new_n254), .B1(new_n273), .B2(new_n256), .ZN(new_n600));
  INV_X1    g0400(.A(new_n256), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n451), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n592), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n591), .A2(new_n305), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n591), .A2(G200), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n588), .A2(G190), .A3(new_n590), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n451), .A2(G87), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n600), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n584), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n509), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n531), .A2(new_n534), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT22), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n539), .B1(new_n616), .B2(new_n529), .ZN(new_n617));
  INV_X1    g0417(.A(new_n540), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n254), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT85), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n541), .A2(new_n524), .A3(new_n254), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n612), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(G179), .A2(new_n519), .B1(new_n522), .B2(G169), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n545), .B(new_n611), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n448), .A2(new_n502), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g0425(.A(new_n625), .B(KEYINPUT88), .Z(G372));
  NAND2_X1  g0426(.A1(new_n362), .A2(new_n365), .ZN(new_n627));
  INV_X1    g0427(.A(new_n437), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n308), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n444), .A2(new_n438), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n353), .A2(new_n355), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n401), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n447), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT90), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n577), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n600), .A2(new_n607), .A3(new_n608), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n588), .A2(KEYINPUT89), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT89), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(new_n587), .B2(new_n284), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n590), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G200), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n305), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n638), .A2(new_n643), .B1(new_n603), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n561), .A2(new_n574), .A3(KEYINPUT90), .A4(new_n576), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n637), .A2(new_n645), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n603), .A2(new_n644), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT26), .B1(new_n610), .B2(new_n577), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n584), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n545), .A2(new_n652), .A3(new_n645), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n509), .B1(new_n542), .B2(new_n544), .ZN(new_n655));
  INV_X1    g0455(.A(new_n623), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n496), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n651), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n635), .B1(new_n448), .B2(new_n659), .ZN(G369));
  INV_X1    g0460(.A(KEYINPUT91), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n217), .A2(new_n268), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G213), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(KEYINPUT27), .B2(new_n662), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(G343), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n468), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n661), .B1(new_n496), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n495), .A2(KEYINPUT91), .A3(new_n669), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n668), .B(new_n670), .C1(new_n502), .C2(new_n669), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n655), .A2(new_n656), .A3(new_n666), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n657), .A2(new_n545), .ZN(new_n673));
  INV_X1    g0473(.A(new_n666), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n622), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n672), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n671), .A2(G330), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n655), .A2(new_n656), .A3(new_n674), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n657), .A2(new_n495), .A3(new_n545), .A4(new_n674), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n213), .ZN(new_n681));
  OR3_X1    g0481(.A1(new_n681), .A2(KEYINPUT92), .A3(G41), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT92), .B1(new_n681), .B2(G41), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n595), .A2(G116), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n685), .A2(new_n209), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n222), .B2(new_n685), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT28), .Z(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT93), .B1(new_n659), .B2(new_n666), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT29), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n495), .B1(new_n655), .B2(new_n656), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n653), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT93), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(new_n696), .A3(new_n674), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n691), .A2(new_n692), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n637), .A2(new_n645), .A3(new_n647), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT26), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n649), .B(KEYINPUT94), .Z(new_n701));
  NOR3_X1   g0501(.A1(new_n610), .A2(KEYINPUT26), .A3(new_n577), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n584), .A2(KEYINPUT95), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT95), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n577), .A2(new_n583), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n545), .A2(new_n645), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n700), .B(new_n703), .C1(new_n707), .C2(new_n694), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n692), .B1(new_n708), .B2(new_n674), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n698), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  INV_X1    g0512(.A(new_n489), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n487), .ZN(new_n714));
  INV_X1    g0514(.A(new_n494), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n492), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n714), .A2(new_n716), .A3(new_n501), .A4(new_n674), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n657), .A3(new_n545), .A4(new_n611), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  AND4_X1   g0520(.A1(new_n514), .A2(new_n515), .A3(new_n588), .A4(new_n590), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n491), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n722), .B2(new_n582), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n560), .A2(new_n721), .A3(new_n491), .A4(KEYINPUT30), .ZN(new_n724));
  AOI21_X1  g0524(.A(G179), .B1(new_n480), .B2(new_n485), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n582), .A2(new_n518), .A3(new_n725), .A4(new_n642), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT31), .B1(new_n727), .B2(new_n666), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n712), .B1(new_n719), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n711), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n690), .B1(new_n732), .B2(G1), .ZN(G364));
  NOR2_X1   g0533(.A1(new_n336), .A2(new_n267), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G45), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G1), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n685), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT96), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n218), .B1(G20), .B2(new_n305), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n336), .B1(new_n500), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n563), .ZN(new_n746));
  INV_X1    g0546(.A(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G179), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(G20), .A3(G190), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n278), .B1(new_n750), .B2(G87), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n350), .A2(new_n500), .A3(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n336), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n350), .A2(new_n747), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n336), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n500), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n751), .B1(new_n202), .B2(new_n753), .C1(new_n757), .C2(new_n201), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n336), .A2(new_n500), .A3(new_n754), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n746), .B(new_n758), .C1(G68), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n217), .A2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n743), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G159), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT32), .Z(new_n766));
  NAND2_X1  g0566(.A1(new_n762), .A2(new_n748), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT100), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G107), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n350), .A2(G200), .ZN(new_n770));
  AND3_X1   g0570(.A1(new_n762), .A2(KEYINPUT99), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(KEYINPUT99), .B1(new_n762), .B2(new_n770), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G77), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n761), .A2(new_n766), .A3(new_n769), .A4(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G283), .A2(new_n768), .B1(new_n773), .B2(G311), .ZN(new_n776));
  INV_X1    g0576(.A(G303), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n278), .B1(new_n749), .B2(new_n777), .C1(new_n753), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G326), .B2(new_n756), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n760), .A2(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n764), .A2(G329), .B1(G294), .B2(new_n744), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n776), .A2(new_n780), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n741), .B1(new_n775), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G13), .A2(G33), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n741), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT98), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n248), .A2(new_n289), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n681), .A2(new_n315), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(G45), .B2(new_n221), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT97), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n681), .A2(new_n278), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G355), .B1(new_n454), .B2(new_n681), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n739), .B(new_n785), .C1(new_n791), .C2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n671), .B2(new_n789), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT101), .Z(new_n803));
  NAND2_X1  g0603(.A1(new_n671), .A2(G330), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n685), .B2(new_n736), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n671), .A2(G330), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NOR2_X1   g0609(.A1(new_n307), .A2(new_n666), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n369), .A2(new_n372), .B1(new_n275), .B2(new_n666), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(new_n308), .ZN(new_n813));
  INV_X1    g0613(.A(new_n697), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n696), .B1(new_n695), .B2(new_n674), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n813), .A2(new_n666), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n695), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n730), .B1(new_n624), .B2(new_n717), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G330), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n737), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n821), .B2(new_n819), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n278), .B1(new_n750), .B2(G50), .ZN(new_n824));
  INV_X1    g0624(.A(new_n764), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n824), .B1(new_n745), .B2(new_n202), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n753), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n756), .A2(G137), .B1(new_n828), .B2(G143), .ZN(new_n829));
  INV_X1    g0629(.A(G150), .ZN(new_n830));
  INV_X1    g0630(.A(new_n773), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n830), .B2(new_n759), .C1(new_n831), .C2(new_n320), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT34), .Z(new_n833));
  AOI211_X1 g0633(.A(new_n827), .B(new_n833), .C1(G68), .C2(new_n768), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n278), .B1(new_n749), .B2(new_n279), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n835), .B(new_n746), .C1(G294), .C2(new_n828), .ZN(new_n836));
  INV_X1    g0636(.A(G283), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n757), .A2(new_n777), .B1(new_n837), .B2(new_n759), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G311), .B2(new_n764), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n768), .A2(G87), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n773), .A2(G116), .ZN(new_n841));
  AND4_X1   g0641(.A1(new_n836), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n740), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n740), .A2(new_n786), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n739), .B1(new_n206), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n813), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n843), .B(new_n845), .C1(new_n787), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n823), .A2(new_n847), .ZN(G384));
  OR2_X1    g0648(.A1(new_n568), .A2(KEYINPUT35), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n568), .A2(KEYINPUT35), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n849), .A2(G116), .A3(new_n219), .A4(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT36), .Z(new_n852));
  NAND4_X1  g0652(.A1(new_n222), .A2(G77), .A3(new_n326), .A4(new_n327), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n203), .A2(G50), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT102), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n209), .B(G13), .C1(new_n853), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n448), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n634), .B1(new_n711), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT39), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT16), .B1(new_n319), .B2(new_n329), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n314), .B1(new_n331), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT103), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT103), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n314), .B(new_n864), .C1(new_n331), .C2(new_n861), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n665), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n366), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT38), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n359), .A2(new_n361), .A3(new_n314), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n340), .A2(new_n665), .ZN(new_n872));
  AND4_X1   g0672(.A1(new_n870), .A2(new_n871), .A3(new_n352), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n863), .A2(new_n351), .A3(new_n865), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n866), .A2(new_n874), .A3(new_n871), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(KEYINPUT37), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n366), .A2(new_n340), .A3(new_n665), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n871), .A2(new_n352), .A3(new_n872), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n871), .A2(new_n870), .A3(new_n352), .A4(new_n872), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n860), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  INV_X1    g0685(.A(new_n868), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n885), .B1(new_n876), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n875), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n881), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(KEYINPUT38), .A3(new_n868), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n887), .A2(new_n890), .A3(KEYINPUT39), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n630), .A2(new_n666), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n884), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n632), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n894), .A2(new_n665), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n810), .B1(new_n695), .B2(new_n817), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n889), .B2(new_n868), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n898), .A2(new_n877), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n438), .A2(new_n666), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n628), .A2(new_n630), .A3(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n438), .B(new_n666), .C1(new_n437), .C2(new_n444), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n897), .A2(new_n899), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n896), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n859), .B(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n813), .B1(new_n901), .B2(new_n902), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n820), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n910), .B2(new_n899), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT40), .B1(new_n877), .B2(new_n883), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n858), .A2(new_n820), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(G330), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n209), .B2(new_n734), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n907), .A2(new_n917), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n857), .B1(new_n919), .B2(new_n920), .ZN(G367));
  NAND2_X1  g0721(.A1(new_n600), .A2(new_n608), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n666), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n645), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n649), .B2(new_n923), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT104), .ZN(new_n927));
  INV_X1    g0727(.A(new_n679), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n666), .A2(new_n574), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n704), .A2(new_n706), .A3(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n577), .A2(new_n674), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n577), .B1(new_n930), .B2(new_n657), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n674), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n927), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n677), .B1(new_n930), .B2(new_n931), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n684), .B(KEYINPUT41), .ZN(new_n944));
  INV_X1    g0744(.A(new_n711), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT107), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n495), .A2(new_n674), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n672), .B(new_n947), .C1(new_n673), .C2(new_n675), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n804), .A2(new_n679), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n679), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(G330), .A3(new_n671), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n945), .A2(new_n946), .A3(new_n821), .A4(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT106), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n930), .A2(new_n931), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n679), .B2(new_n678), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n954), .A2(new_n955), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n679), .A2(new_n678), .A3(new_n932), .ZN(new_n961));
  XNOR2_X1  g0761(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n960), .A2(new_n677), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n677), .B1(new_n960), .B2(new_n964), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n952), .A2(new_n821), .A3(new_n710), .A4(new_n698), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT107), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n953), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n944), .B1(new_n970), .B2(new_n732), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n943), .B1(new_n971), .B2(new_n736), .ZN(new_n972));
  INV_X1    g0772(.A(new_n793), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n791), .B1(new_n213), .B2(new_n256), .C1(new_n241), .C2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n739), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n773), .A2(G50), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n315), .B1(new_n749), .B2(new_n202), .C1(new_n753), .C2(new_n830), .ZN(new_n979));
  INV_X1    g0779(.A(new_n767), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n979), .B1(G77), .B2(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G143), .A2(new_n756), .B1(new_n760), .B2(G159), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n764), .A2(G137), .B1(G68), .B2(new_n744), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n978), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n749), .A2(new_n454), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT46), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n315), .B(new_n986), .C1(G303), .C2(new_n828), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n980), .A2(G97), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n764), .A2(G317), .B1(new_n760), .B2(G294), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n756), .A2(G311), .B1(G107), .B2(new_n744), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n831), .A2(new_n837), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n984), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT47), .Z(new_n994));
  OAI221_X1 g0794(.A(new_n977), .B1(new_n789), .B2(new_n925), .C1(new_n994), .C2(new_n741), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n972), .A2(new_n995), .ZN(G387));
  AOI22_X1  g0796(.A1(new_n798), .A2(new_n687), .B1(new_n279), .B2(new_n681), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n687), .A2(KEYINPUT109), .ZN(new_n998));
  NAND2_X1  g0798(.A1(G68), .A2(G77), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(new_n289), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(KEYINPUT109), .B2(new_n687), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n258), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n201), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT50), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n973), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1007), .A2(KEYINPUT110), .B1(new_n238), .B2(new_n289), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1007), .A2(KEYINPUT110), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n997), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1010), .A2(new_n791), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n315), .B1(new_n753), .B2(new_n201), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n757), .A2(new_n320), .B1(new_n258), .B2(new_n759), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n601), .C2(new_n744), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n764), .A2(G150), .B1(G77), .B2(new_n750), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT111), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n773), .A2(G68), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n768), .A2(G97), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n744), .A2(G283), .B1(new_n750), .B2(G294), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G311), .A2(new_n760), .B1(new_n828), .B2(G317), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n778), .B2(new_n757), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G303), .B2(new_n773), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1020), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT112), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(KEYINPUT48), .B2(new_n1023), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT113), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(KEYINPUT113), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(KEYINPUT49), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n315), .B1(new_n764), .B2(G326), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n454), .C2(new_n767), .ZN(new_n1033));
  AOI21_X1  g0833(.A(KEYINPUT49), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1019), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n739), .B(new_n1011), .C1(new_n1035), .C2(new_n740), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n676), .A2(new_n789), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1036), .A2(new_n1037), .B1(new_n736), .B2(new_n952), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n968), .A2(new_n685), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n732), .B2(new_n952), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(G393));
  INV_X1    g0841(.A(new_n967), .ZN(new_n1042));
  AND3_X1   g0842(.A1(new_n1042), .A2(KEYINPUT115), .A3(new_n968), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT115), .B1(new_n1042), .B2(new_n968), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n685), .B(new_n970), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n930), .A2(new_n788), .A3(new_n931), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n791), .B1(new_n563), .B2(new_n213), .C1(new_n245), .C2(new_n973), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT114), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n738), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n745), .A2(new_n206), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n278), .B(new_n1052), .C1(G68), .C2(new_n750), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n773), .A2(new_n1002), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n764), .A2(G143), .B1(new_n760), .B2(G50), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1053), .A2(new_n840), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n756), .A2(G150), .B1(new_n828), .B2(G159), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT51), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n773), .A2(G294), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n278), .B1(new_n749), .B2(new_n837), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n760), .B2(G303), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n764), .A2(G322), .B1(G116), .B2(new_n744), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n769), .A2(new_n1059), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n756), .A2(G317), .B1(new_n828), .B2(G311), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT52), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1056), .A2(new_n1058), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1049), .B(new_n1051), .C1(new_n740), .C2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n967), .A2(new_n736), .B1(new_n1046), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1045), .A2(new_n1068), .ZN(G390));
  NOR3_X1   g0869(.A1(new_n821), .A2(new_n813), .A3(new_n904), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(KEYINPUT116), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n818), .A2(new_n811), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n903), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n892), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1074), .A2(new_n1075), .B1(new_n884), .B2(new_n891), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n878), .A2(new_n882), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n885), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n892), .B1(new_n890), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n708), .A2(new_n674), .A3(new_n846), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n811), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1080), .B1(new_n1082), .B2(new_n903), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1072), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1083), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n884), .A2(new_n891), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n897), .A2(new_n904), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n892), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1088), .A3(new_n1071), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n903), .B1(new_n731), .B2(new_n846), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1073), .B1(new_n1091), .B2(new_n1070), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n904), .B1(new_n821), .B2(new_n813), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n731), .A2(new_n846), .A3(new_n903), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1093), .A2(new_n1094), .A3(new_n811), .A4(new_n1081), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n858), .A2(new_n731), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n859), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n684), .B1(new_n1090), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1090), .B2(new_n1098), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1090), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1086), .A2(new_n786), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n844), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n738), .B1(new_n1002), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(G294), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n825), .A2(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n757), .A2(new_n837), .B1(new_n279), .B2(new_n759), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n278), .B1(new_n749), .B2(new_n343), .C1(new_n753), .C2(new_n454), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1052), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n768), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1109), .B1(new_n203), .B2(new_n1110), .C1(new_n563), .C2(new_n831), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n315), .B1(new_n767), .B2(new_n201), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G125), .B2(new_n764), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT117), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n756), .A2(G128), .ZN(new_n1115));
  INV_X1    g0915(.A(G137), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n759), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G159), .B2(new_n744), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n749), .A2(new_n830), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT53), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n1119), .A2(new_n1120), .B1(new_n826), .B2(new_n753), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n1120), .B2(new_n1119), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1118), .B(new_n1122), .C1(new_n831), .C2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1111), .B1(new_n1114), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1104), .B1(new_n1125), .B2(new_n740), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1101), .A2(new_n736), .B1(new_n1102), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1100), .A2(new_n1127), .ZN(G378));
  NAND3_X1  g0928(.A1(new_n397), .A2(new_n400), .A3(new_n447), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n393), .A2(new_n665), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n397), .A2(new_n400), .A3(new_n447), .A4(new_n1130), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n786), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n278), .A2(new_n288), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n750), .B2(G77), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n202), .B2(new_n767), .C1(new_n825), .C2(new_n837), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT118), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n756), .A2(G116), .B1(G68), .B2(new_n744), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT119), .Z(new_n1144));
  AOI22_X1  g0944(.A1(G97), .A2(new_n760), .B1(new_n828), .B2(G107), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n256), .C2(new_n831), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT58), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(KEYINPUT58), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1139), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1123), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n828), .A2(G128), .B1(new_n750), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G150), .B2(new_n744), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G125), .A2(new_n756), .B1(new_n760), .B2(G132), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n831), .C2(new_n1116), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n980), .A2(G159), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G33), .B(G41), .C1(new_n764), .C2(G124), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n740), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n844), .A2(new_n201), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1138), .A2(new_n737), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n820), .A2(new_n909), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n887), .A2(new_n890), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT40), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(G330), .B1(new_n910), .B2(new_n912), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1134), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1169), .A2(new_n1170), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n908), .B1(new_n890), .B2(new_n1078), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n712), .B1(new_n1167), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1137), .B1(new_n1178), .B2(new_n911), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n906), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1175), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1073), .A2(new_n1168), .A3(new_n903), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n895), .A3(new_n893), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1178), .A2(new_n911), .A3(new_n1137), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1181), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1180), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1166), .B1(new_n1186), .B2(new_n736), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n711), .A2(new_n858), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n635), .A3(new_n1097), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT120), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT120), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n859), .A2(new_n1191), .A3(new_n1097), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(new_n1090), .C2(new_n1098), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT121), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT121), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n906), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n685), .B1(new_n1194), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1193), .B2(new_n1186), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1187), .B1(new_n1200), .B2(new_n1201), .ZN(G375));
  NAND2_X1  g1002(.A1(new_n904), .A2(new_n786), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n738), .B1(G68), .B2(new_n1103), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n773), .A2(G150), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n315), .B1(new_n749), .B2(new_n320), .C1(new_n753), .C2(new_n1116), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G58), .B2(new_n980), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n764), .A2(G128), .B1(new_n760), .B2(new_n1151), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n756), .A2(G132), .B1(G50), .B2(new_n744), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1205), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n773), .A2(G107), .B1(G116), .B2(new_n760), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT122), .Z(new_n1212));
  OAI221_X1 g1012(.A(new_n278), .B1(new_n563), .B2(new_n749), .C1(new_n757), .C2(new_n1105), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G303), .B2(new_n764), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n745), .A2(new_n256), .B1(new_n837), .B2(new_n753), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT123), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(new_n206), .C2(new_n1110), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1210), .B1(new_n1212), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1204), .B1(new_n1218), .B2(new_n740), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1096), .A2(new_n736), .B1(new_n1203), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n944), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1098), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1096), .B1(new_n859), .B2(new_n1097), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1220), .B1(new_n1222), .B2(new_n1223), .ZN(G381));
  NOR2_X1   g1024(.A1(G393), .A2(G396), .ZN(new_n1225));
  INV_X1    g1025(.A(G384), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1227), .A2(G390), .A3(G381), .ZN(new_n1228));
  INV_X1    g1028(.A(G387), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1100), .A2(new_n1127), .ZN(new_n1230));
  INV_X1    g1030(.A(G375), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(G407));
  INV_X1    g1032(.A(G343), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1231), .A2(new_n1233), .A3(new_n1230), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(G407), .A2(G213), .A3(new_n1234), .ZN(G409));
  NAND3_X1  g1035(.A1(G387), .A2(new_n1045), .A3(new_n1068), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT127), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(G393), .B(G396), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1229), .A2(G390), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1236), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(G387), .B(G390), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n1238), .A3(new_n1237), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1223), .A2(KEYINPUT60), .A3(new_n1098), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n685), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1223), .B1(KEYINPUT60), .B2(new_n1098), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1220), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1226), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G384), .B(new_n1220), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1233), .A2(G213), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT125), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n736), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(KEYINPUT124), .A3(new_n1165), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1193), .A2(new_n1221), .A3(new_n1186), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT124), .B1(new_n1257), .B2(new_n1165), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1256), .B(new_n1230), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G378), .B(new_n1187), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1257), .A2(new_n1165), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT124), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1259), .A3(new_n1258), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1256), .B1(new_n1268), .B2(new_n1230), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1254), .B(new_n1255), .C1(new_n1264), .C2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT126), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1230), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT125), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT62), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1255), .B1(new_n1264), .B2(new_n1269), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1233), .A2(G213), .A3(G2897), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1253), .B(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1270), .A2(KEYINPUT62), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1246), .B1(new_n1277), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1271), .A2(new_n1285), .A3(new_n1276), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1270), .A2(new_n1285), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1286), .A2(new_n1245), .A3(new_n1281), .A4(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1284), .A2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(G375), .A2(new_n1230), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1263), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1244), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1243), .B1(new_n1238), .B2(new_n1237), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1242), .A2(new_n1244), .A3(new_n1291), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1295), .A2(new_n1254), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1254), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(G402));
endmodule


