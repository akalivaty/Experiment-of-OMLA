//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g023(.A(G2106), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n449), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n459), .A2(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(new_n454), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n459), .A2(KEYINPUT67), .B1(G567), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  OR3_X1    g047(.A1(new_n472), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n467), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n472), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n468), .A2(new_n477), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n471), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(G160));
  INV_X1    g057(.A(new_n474), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(KEYINPUT70), .A3(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n470), .A2(G2105), .A3(new_n473), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n474), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n484), .A2(new_n487), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NAND2_X1  g069(.A1(new_n486), .A2(G126), .ZN(new_n495));
  OR3_X1    g070(.A1(new_n471), .A2(KEYINPUT71), .A3(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT71), .B1(new_n471), .B2(G114), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n496), .A2(G2104), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n468), .A2(new_n477), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR4_X1   g077(.A1(new_n501), .A2(KEYINPUT4), .A3(new_n502), .A4(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT4), .B1(new_n474), .B2(new_n502), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n506), .B(KEYINPUT4), .C1(new_n474), .C2(new_n502), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n500), .B1(new_n505), .B2(new_n507), .ZN(G164));
  AND2_X1   g083(.A1(KEYINPUT73), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT73), .A2(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT6), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n511), .A2(G50), .A3(G543), .A4(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n511), .A2(G88), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT73), .B(G651), .ZN(new_n518));
  AND2_X1   g093(.A1(G75), .A2(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n516), .B2(G62), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n515), .B(new_n517), .C1(new_n518), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT74), .ZN(new_n522));
  INV_X1    g097(.A(new_n518), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n525), .A2(new_n527), .A3(G62), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n523), .B1(new_n528), .B2(new_n519), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n529), .A2(new_n530), .A3(new_n515), .A4(new_n517), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n522), .A2(new_n531), .ZN(G166));
  NAND3_X1  g107(.A1(new_n511), .A2(G543), .A3(new_n514), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n511), .A2(new_n514), .A3(new_n516), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT7), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n535), .A2(new_n538), .A3(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(new_n537), .A2(G90), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n534), .A2(G52), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n518), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  AOI22_X1  g127(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n518), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n513), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n555));
  XOR2_X1   g130(.A(KEYINPUT75), .B(G43), .Z(new_n556));
  NAND3_X1  g131(.A1(new_n555), .A2(G543), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(G81), .A3(new_n516), .ZN(new_n558));
  AND3_X1   g133(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n566), .A2(new_n536), .B1(new_n567), .B2(new_n512), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n534), .A2(new_n569), .A3(G53), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT9), .B1(new_n533), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G299));
  INV_X1    g149(.A(G166), .ZN(G303));
  NAND4_X1  g150(.A1(new_n511), .A2(G49), .A3(G543), .A4(new_n514), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n511), .A2(G87), .A3(new_n514), .A4(new_n516), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  NAND3_X1  g154(.A1(new_n555), .A2(G86), .A3(new_n516), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n555), .A2(G48), .A3(G543), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n580), .B(new_n581), .C1(new_n518), .C2(new_n582), .ZN(G305));
  NAND4_X1  g158(.A1(new_n511), .A2(G85), .A3(new_n514), .A4(new_n516), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n511), .A2(G47), .A3(G543), .A4(new_n514), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n584), .B(new_n585), .C1(new_n586), .C2(new_n518), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n516), .A2(G66), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n512), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G54), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n593), .B1(new_n533), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n511), .A2(KEYINPUT76), .A3(G543), .A4(new_n514), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n555), .A2(KEYINPUT10), .A3(G92), .A4(new_n516), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n511), .A2(G92), .A3(new_n514), .A4(new_n516), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n597), .A2(KEYINPUT77), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(KEYINPUT77), .B1(new_n597), .B2(new_n602), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n589), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n533), .A2(new_n594), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n606), .A2(G54), .A3(new_n596), .ZN(new_n607));
  INV_X1    g182(.A(new_n592), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n602), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n597), .A2(KEYINPUT77), .A3(new_n602), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n611), .A2(KEYINPUT78), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n588), .B1(new_n614), .B2(G868), .ZN(G321));
  XOR2_X1   g190(.A(G321), .B(KEYINPUT79), .Z(G284));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n573), .ZN(G297));
  XNOR2_X1  g193(.A(G297), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n614), .B1(new_n620), .B2(G860), .ZN(G148));
  NOR3_X1   g196(.A1(new_n603), .A2(new_n604), .A3(new_n589), .ZN(new_n622));
  AOI21_X1  g197(.A(KEYINPUT78), .B1(new_n611), .B2(new_n612), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(G111), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n628), .A2(KEYINPUT82), .B1(new_n629), .B2(G2105), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(KEYINPUT82), .B2(new_n628), .ZN(new_n631));
  INV_X1    g206(.A(G135), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n631), .B1(new_n474), .B2(new_n632), .C1(new_n633), .C2(new_n485), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2096), .Z(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n636));
  NOR3_X1   g211(.A1(new_n472), .A2(new_n465), .A3(G2105), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT13), .B(G2100), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n635), .A2(new_n640), .ZN(G156));
  INV_X1    g216(.A(KEYINPUT86), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT84), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2430), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT85), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n642), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(G14), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n657), .B2(new_n659), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n655), .A2(new_n656), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n655), .A2(new_n656), .ZN(new_n664));
  NAND4_X1  g239(.A1(new_n663), .A2(KEYINPUT86), .A3(new_n658), .A4(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2067), .B(G2678), .Z(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  AND3_X1   g250(.A1(new_n675), .A2(KEYINPUT17), .A3(new_n672), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n672), .B1(new_n675), .B2(KEYINPUT17), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n676), .A2(new_n677), .A3(new_n671), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XOR2_X1   g258(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n689), .A2(KEYINPUT88), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(KEYINPUT88), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n692), .A2(new_n685), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n695));
  OAI221_X1 g270(.A(new_n691), .B1(new_n686), .B2(new_n690), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1991), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G1996), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(G1996), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n682), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(new_n682), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n703), .A2(new_n704), .A3(new_n699), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n702), .B2(new_n705), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(G229));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n477), .A3(G127), .ZN(new_n710));
  NAND2_X1  g285(.A1(G115), .A2(G2104), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n471), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n466), .A2(G103), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT25), .ZN(new_n714));
  AOI211_X1 g289(.A(new_n712), .B(new_n714), .C1(G139), .C2(new_n483), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G29), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G29), .B2(G33), .ZN(new_n717));
  INV_X1    g292(.A(G2072), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT31), .B(G11), .Z(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G28), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT94), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n723), .A2(KEYINPUT94), .B1(new_n722), .B2(G28), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n720), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n719), .B(new_n726), .C1(new_n721), .C2(new_n634), .ZN(new_n727));
  NOR2_X1   g302(.A1(G16), .A2(G21), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G168), .B2(G16), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1966), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n717), .A2(new_n718), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n727), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n721), .A2(G26), .ZN(new_n733));
  OR2_X1    g308(.A1(G104), .A2(G2105), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n734), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n735));
  INV_X1    g310(.A(G140), .ZN(new_n736));
  INV_X1    g311(.A(G128), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n735), .B1(new_n474), .B2(new_n736), .C1(new_n737), .C2(new_n485), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(new_n721), .ZN(new_n740));
  MUX2_X1   g315(.A(new_n733), .B(new_n740), .S(KEYINPUT28), .Z(new_n741));
  INV_X1    g316(.A(G2067), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  AND2_X1   g318(.A1(KEYINPUT89), .A2(G16), .ZN(new_n744));
  NOR2_X1   g319(.A1(KEYINPUT89), .A2(G16), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G19), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n746), .ZN(new_n750));
  INV_X1    g325(.A(G1341), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NOR2_X1   g328(.A1(G5), .A2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G171), .B2(G16), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n753), .B1(new_n755), .B2(G1961), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n752), .B(new_n756), .C1(G1961), .C2(new_n755), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n732), .A2(new_n743), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n721), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n721), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G29), .A2(G35), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G162), .B2(G29), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n762), .B1(new_n766), .B2(G2090), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n721), .A2(G32), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT26), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n771), .A2(new_n772), .B1(G105), .B2(new_n466), .ZN(new_n773));
  INV_X1    g348(.A(G129), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n485), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G141), .B2(new_n483), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT92), .Z(new_n777));
  OAI21_X1  g352(.A(new_n768), .B1(new_n777), .B2(new_n721), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT27), .B(G1996), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT93), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n782), .B2(KEYINPUT24), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n783), .A2(new_n784), .B1(KEYINPUT24), .B2(new_n782), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G160), .B2(G29), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G2084), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(G2084), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n778), .A2(new_n780), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n781), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n758), .A2(new_n767), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G4), .A2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n614), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1348), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n766), .A2(G2090), .ZN(new_n797));
  OAI21_X1  g372(.A(G20), .B1(new_n744), .B2(new_n745), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT23), .Z(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G299), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1956), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT96), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n792), .A2(new_n796), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n746), .A2(G22), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G166), .B2(new_n746), .ZN(new_n806));
  INV_X1    g381(.A(G1971), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G16), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G6), .ZN(new_n810));
  INV_X1    g385(.A(G305), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n809), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT32), .B(G1981), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n809), .A2(G23), .ZN(new_n815));
  INV_X1    g390(.A(G288), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n809), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT33), .B(G1976), .Z(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT90), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n808), .A2(new_n814), .A3(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT34), .Z(new_n822));
  MUX2_X1   g397(.A(G24), .B(G290), .S(new_n746), .Z(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(G1986), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n721), .A2(G25), .ZN(new_n825));
  OR2_X1    g400(.A1(G95), .A2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n827));
  INV_X1    g402(.A(G131), .ZN(new_n828));
  INV_X1    g403(.A(G119), .ZN(new_n829));
  OAI221_X1 g404(.A(new_n827), .B1(new_n474), .B2(new_n828), .C1(new_n829), .C2(new_n485), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(new_n721), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT35), .B(G1991), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n822), .A2(new_n824), .A3(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(KEYINPUT36), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(KEYINPUT36), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n804), .B1(new_n837), .B2(new_n838), .ZN(G311));
  XOR2_X1   g414(.A(G311), .B(KEYINPUT97), .Z(G150));
  INV_X1    g415(.A(G55), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n533), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n525), .A2(new_n527), .ZN(new_n845));
  INV_X1    g420(.A(G67), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n523), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT99), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n537), .A2(G93), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(new_n851), .A3(new_n523), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n843), .A2(new_n849), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n614), .A2(G559), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT39), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT98), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n853), .A2(new_n559), .ZN(new_n862));
  AOI22_X1  g437(.A1(G55), .A2(new_n534), .B1(new_n537), .B2(G93), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n749), .A2(new_n863), .A3(new_n849), .A4(new_n852), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n860), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n866), .B1(new_n860), .B2(new_n861), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n855), .B1(new_n869), .B2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(G160), .B(new_n634), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n638), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n715), .A2(new_n776), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n777), .B2(new_n715), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n873), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n483), .A2(G142), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n471), .A2(G118), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(G130), .B2(new_n486), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n739), .ZN(new_n882));
  XNOR2_X1  g457(.A(G164), .B(new_n831), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n493), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n876), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(KEYINPUT100), .B(G37), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n876), .A2(new_n885), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g465(.A1(new_n816), .A2(G290), .ZN(new_n891));
  NAND2_X1  g466(.A1(G72), .A2(G543), .ZN(new_n892));
  INV_X1    g467(.A(G60), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n845), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n523), .ZN(new_n895));
  NAND4_X1  g470(.A1(G288), .A2(new_n584), .A3(new_n895), .A4(new_n585), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n522), .A2(G305), .A3(new_n531), .ZN(new_n898));
  AOI21_X1  g473(.A(G305), .B1(new_n522), .B2(new_n531), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(G166), .A2(new_n811), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n522), .A2(G305), .A3(new_n531), .ZN(new_n902));
  XNOR2_X1  g477(.A(G290), .B(G288), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI211_X1 g479(.A(KEYINPUT101), .B(KEYINPUT102), .C1(new_n900), .C2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(new_n904), .A3(KEYINPUT101), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n900), .A2(new_n904), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT42), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n908), .A2(new_n909), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n898), .A2(new_n899), .A3(new_n897), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n903), .B1(new_n901), .B2(new_n902), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n916), .B(new_n911), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n915), .B1(new_n919), .B2(new_n906), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT103), .B1(new_n920), .B2(new_n912), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n573), .A2(new_n609), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n573), .A2(new_n609), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT41), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(KEYINPUT41), .A3(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n866), .B1(new_n614), .B2(new_n620), .ZN(new_n929));
  AOI211_X1 g504(.A(G559), .B(new_n865), .C1(new_n605), .C2(new_n613), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n624), .A2(new_n865), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n614), .A2(new_n620), .A3(new_n866), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n924), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n914), .A2(new_n921), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(KEYINPUT104), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n931), .A2(new_n934), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n909), .B1(new_n908), .B2(new_n913), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n920), .A2(KEYINPUT103), .A3(new_n912), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n914), .A2(new_n921), .A3(new_n935), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(G868), .B1(new_n937), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n853), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(G868), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n936), .A2(KEYINPUT104), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n941), .A3(new_n943), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n951), .B2(G868), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n947), .B1(new_n946), .B2(new_n952), .ZN(G295));
  INV_X1    g528(.A(new_n949), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n946), .B1(new_n945), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT105), .B1(new_n951), .B2(G868), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT106), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n947), .B(new_n958), .C1(new_n946), .C2(new_n952), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n957), .A2(new_n959), .ZN(G331));
  NAND2_X1  g535(.A1(new_n910), .A2(new_n916), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n961), .A2(new_n906), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n964));
  OAI21_X1  g539(.A(G286), .B1(G171), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(G301), .A2(KEYINPUT107), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(new_n866), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(KEYINPUT108), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n967), .B(new_n866), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n970), .B2(KEYINPUT108), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n971), .A2(new_n924), .ZN(new_n972));
  INV_X1    g547(.A(new_n970), .ZN(new_n973));
  INV_X1    g548(.A(new_n928), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n963), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n924), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(new_n962), .C1(new_n971), .C2(new_n974), .ZN(new_n978));
  AND4_X1   g553(.A1(KEYINPUT43), .A2(new_n976), .A3(new_n887), .A4(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G37), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n971), .B2(new_n974), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n963), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT43), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT44), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n981), .B2(new_n983), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n976), .A2(new_n887), .A3(new_n978), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n987), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n985), .B1(new_n989), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g565(.A(new_n738), .B(G2067), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1996), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n993), .B2(new_n776), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n993), .B2(new_n777), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n830), .B(new_n833), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT112), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n504), .A2(KEYINPUT72), .ZN(new_n1000));
  INV_X1    g575(.A(new_n503), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n507), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n500), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1384), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1384), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(KEYINPUT109), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n481), .A2(G40), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1008), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G290), .A2(G1986), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT110), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n999), .A2(new_n1014), .B1(new_n1017), .B2(KEYINPUT48), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1017), .A2(KEYINPUT48), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n831), .A2(new_n834), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT125), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n995), .A2(new_n1021), .B1(new_n742), .B2(new_n739), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n1018), .A2(new_n1019), .B1(new_n1014), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1013), .A2(new_n993), .ZN(new_n1024));
  NAND2_X1  g599(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1025));
  XOR2_X1   g600(.A(new_n1024), .B(new_n1025), .Z(new_n1026));
  INV_X1    g601(.A(KEYINPUT127), .ZN(new_n1027));
  NOR2_X1   g602(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n992), .A2(new_n776), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n1013), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1027), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1033));
  OR3_X1    g608(.A1(new_n1032), .A2(KEYINPUT47), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT47), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1023), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1010), .A2(KEYINPUT45), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1009), .B1(G164), .B2(G1384), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1012), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n761), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1010), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n1040), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1961), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1037), .A2(new_n1041), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n476), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n476), .A2(new_n1048), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT123), .ZN(new_n1051));
  OAI211_X1 g626(.A(KEYINPUT53), .B(G40), .C1(new_n1051), .C2(G2078), .ZN(new_n1052));
  AOI211_X1 g627(.A(new_n1052), .B(new_n480), .C1(new_n1051), .C2(G2078), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1049), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1038), .B(new_n1054), .C1(new_n1008), .C2(new_n1011), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1047), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G171), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1012), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1060), .A2(KEYINPUT53), .A3(new_n761), .A4(new_n1038), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1047), .A2(G301), .A3(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1062), .A2(KEYINPUT54), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1056), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1059), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G8), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1010), .B2(new_n1040), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n816), .A2(G1976), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT52), .ZN(new_n1070));
  INV_X1    g645(.A(G1976), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(G288), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1067), .A2(new_n1068), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G305), .A2(G1981), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n582), .A2(new_n518), .ZN(new_n1075));
  INV_X1    g650(.A(G1981), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n581), .A4(new_n580), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1077), .A2(KEYINPUT114), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(KEYINPUT114), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1074), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT49), .B(new_n1074), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1067), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1070), .A2(new_n1073), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(G303), .A2(G8), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT55), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1038), .A2(new_n1040), .A3(new_n1039), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n807), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT113), .B(G2090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1043), .A2(new_n1044), .A3(new_n1040), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1066), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1085), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT115), .B1(new_n1093), .B2(new_n1088), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1040), .B1(new_n1010), .B2(new_n1042), .ZN(new_n1097));
  NOR3_X1   g672(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1099), .A2(new_n1091), .B1(new_n1089), .B2(new_n807), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1096), .B(new_n1087), .C1(new_n1100), .C2(new_n1066), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1094), .A2(new_n1095), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n1103));
  INV_X1    g678(.A(G1966), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1089), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G2084), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1043), .A2(new_n1044), .A3(new_n1106), .A4(new_n1040), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1066), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(G168), .A2(new_n1066), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1103), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1109), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1099), .A2(new_n1106), .B1(new_n1089), .B2(new_n1104), .ZN(new_n1112));
  OAI211_X1 g687(.A(KEYINPUT51), .B(new_n1111), .C1(new_n1112), .C2(new_n1066), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1112), .A2(new_n1111), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1056), .A2(G171), .ZN(new_n1117));
  AOI21_X1  g692(.A(G301), .B1(new_n1047), .B2(new_n1061), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1065), .A2(new_n1102), .A3(new_n1115), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1089), .B2(G1996), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1060), .A2(KEYINPUT120), .A3(new_n993), .A4(new_n1038), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1010), .A2(new_n1040), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(new_n751), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1122), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n559), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT59), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n603), .A2(new_n604), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1099), .A2(G1348), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1124), .A2(G2067), .ZN(new_n1133));
  OAI211_X1 g708(.A(KEYINPUT60), .B(new_n1131), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n795), .B2(new_n1045), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1131), .A2(KEYINPUT60), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1131), .A2(KEYINPUT60), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT56), .B(G2072), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1060), .A2(new_n1038), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(G1956), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1045), .A2(KEYINPUT118), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT118), .B1(new_n1045), .B2(new_n1143), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1142), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n573), .B(KEYINPUT57), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1140), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1147), .B(new_n1142), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1139), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(KEYINPUT119), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1143), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1045), .A2(KEYINPUT118), .A3(new_n1143), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1158), .A2(new_n1159), .A3(new_n1147), .A4(new_n1142), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1152), .A2(new_n1153), .A3(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1130), .B(new_n1151), .C1(new_n1161), .C2(KEYINPUT61), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1131), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1153), .B1(new_n1163), .B2(new_n1135), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1164), .A2(new_n1152), .A3(new_n1160), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1120), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1102), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1115), .A2(KEYINPUT62), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .A4(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1168), .A2(new_n1170), .A3(new_n1118), .ZN(new_n1171));
  NOR4_X1   g746(.A1(new_n1112), .A2(KEYINPUT116), .A3(new_n1066), .A4(G286), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT116), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1108), .B2(G168), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1175), .A2(KEYINPUT63), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1167), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1087), .A2(KEYINPUT117), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1093), .B(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1085), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(KEYINPUT63), .B1(new_n1181), .B2(new_n1175), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1100), .A2(new_n1066), .A3(new_n1087), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1084), .A2(new_n1071), .A3(new_n816), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1184), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1183), .A2(new_n1180), .B1(new_n1185), .B2(new_n1067), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1182), .A2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1166), .A2(new_n1177), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(G290), .A2(G1986), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT111), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1016), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1014), .B1(new_n999), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1036), .B1(new_n1188), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g768(.A1(G227), .A2(new_n463), .ZN(new_n1195));
  NOR3_X1   g769(.A1(new_n707), .A2(new_n708), .A3(new_n1195), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n666), .A2(new_n889), .A3(new_n1196), .ZN(new_n1197));
  NOR2_X1   g771(.A1(new_n989), .A2(new_n1197), .ZN(G308));
  OR2_X1    g772(.A1(new_n989), .A2(new_n1197), .ZN(G225));
endmodule


