

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U548 ( .A1(n714), .A2(n938), .ZN(n515) );
  AND2_X1 U549 ( .A1(n968), .A2(n818), .ZN(n516) );
  NOR2_X1 U550 ( .A1(n806), .A2(n516), .ZN(n517) );
  INV_X1 U551 ( .A(KEYINPUT64), .ZN(n690) );
  INV_X1 U552 ( .A(n727), .ZN(n714) );
  INV_X1 U553 ( .A(KEYINPUT99), .ZN(n757) );
  INV_X1 U554 ( .A(KEYINPUT6), .ZN(n525) );
  OR2_X1 U555 ( .A1(n772), .A2(n771), .ZN(n807) );
  NOR2_X1 U556 ( .A1(G651), .A2(G543), .ZN(n646) );
  XNOR2_X1 U557 ( .A(n525), .B(KEYINPUT76), .ZN(n526) );
  XOR2_X1 U558 ( .A(KEYINPUT65), .B(n518), .Z(n645) );
  XNOR2_X1 U559 ( .A(n527), .B(n526), .ZN(n535) );
  XNOR2_X1 U560 ( .A(KEYINPUT8), .B(KEYINPUT77), .ZN(n537) );
  XOR2_X1 U561 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  NOR2_X1 U562 ( .A1(G651), .A2(n628), .ZN(n518) );
  NAND2_X1 U563 ( .A1(n645), .A2(G51), .ZN(n519) );
  XNOR2_X1 U564 ( .A(KEYINPUT75), .B(n519), .ZN(n524) );
  INV_X1 U565 ( .A(G651), .ZN(n528) );
  NOR2_X1 U566 ( .A1(G543), .A2(n528), .ZN(n521) );
  XNOR2_X1 U567 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n520) );
  XNOR2_X1 U568 ( .A(n521), .B(n520), .ZN(n649) );
  NAND2_X1 U569 ( .A1(n649), .A2(G63), .ZN(n522) );
  XOR2_X1 U570 ( .A(n522), .B(KEYINPUT74), .Z(n523) );
  NOR2_X1 U571 ( .A1(n524), .A2(n523), .ZN(n527) );
  NOR2_X1 U572 ( .A1(n628), .A2(n528), .ZN(n644) );
  NAND2_X1 U573 ( .A1(n644), .A2(G76), .ZN(n529) );
  XNOR2_X1 U574 ( .A(KEYINPUT73), .B(n529), .ZN(n532) );
  NAND2_X1 U575 ( .A1(n646), .A2(G89), .ZN(n530) );
  XOR2_X1 U576 ( .A(KEYINPUT4), .B(n530), .Z(n531) );
  NOR2_X1 U577 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U578 ( .A(KEYINPUT5), .B(n533), .ZN(n534) );
  NOR2_X1 U579 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U580 ( .A(KEYINPUT7), .B(n536), .Z(G168) );
  XNOR2_X1 U581 ( .A(G168), .B(n537), .ZN(G286) );
  AND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n882) );
  NAND2_X1 U583 ( .A1(n882), .A2(G113), .ZN(n546) );
  NOR2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n538) );
  XOR2_X2 U585 ( .A(KEYINPUT17), .B(n538), .Z(n877) );
  NAND2_X1 U586 ( .A1(G137), .A2(n877), .ZN(n540) );
  INV_X1 U587 ( .A(G2105), .ZN(n541) );
  NOR2_X1 U588 ( .A1(G2104), .A2(n541), .ZN(n881) );
  NAND2_X1 U589 ( .A1(G125), .A2(n881), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n544) );
  AND2_X1 U591 ( .A1(n541), .A2(G2104), .ZN(n878) );
  NAND2_X1 U592 ( .A1(G101), .A2(n878), .ZN(n542) );
  XNOR2_X1 U593 ( .A(KEYINPUT23), .B(n542), .ZN(n543) );
  NOR2_X1 U594 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U595 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X2 U596 ( .A(KEYINPUT66), .B(n547), .Z(G160) );
  XNOR2_X1 U597 ( .A(G2446), .B(G2443), .ZN(n557) );
  XOR2_X1 U598 ( .A(G2430), .B(KEYINPUT103), .Z(n549) );
  XNOR2_X1 U599 ( .A(G2454), .B(G2435), .ZN(n548) );
  XNOR2_X1 U600 ( .A(n549), .B(n548), .ZN(n553) );
  XOR2_X1 U601 ( .A(G2438), .B(G2427), .Z(n551) );
  XNOR2_X1 U602 ( .A(G1348), .B(G1341), .ZN(n550) );
  XNOR2_X1 U603 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U604 ( .A(n553), .B(n552), .Z(n555) );
  XNOR2_X1 U605 ( .A(KEYINPUT102), .B(G2451), .ZN(n554) );
  XNOR2_X1 U606 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U607 ( .A(n557), .B(n556), .ZN(n558) );
  AND2_X1 U608 ( .A1(n558), .A2(G14), .ZN(G401) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U610 ( .A(G132), .ZN(G219) );
  INV_X1 U611 ( .A(G82), .ZN(G220) );
  INV_X1 U612 ( .A(G108), .ZN(G238) );
  NAND2_X1 U613 ( .A1(G90), .A2(n646), .ZN(n560) );
  NAND2_X1 U614 ( .A1(G77), .A2(n644), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U616 ( .A(KEYINPUT9), .B(n561), .ZN(n565) );
  NAND2_X1 U617 ( .A1(n645), .A2(G52), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G64), .A2(n649), .ZN(n562) );
  AND2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n565), .A2(n564), .ZN(G301) );
  INV_X1 U621 ( .A(G301), .ZN(G171) );
  NAND2_X1 U622 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U623 ( .A(n566), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U624 ( .A(G223), .ZN(n823) );
  NAND2_X1 U625 ( .A1(n823), .A2(G567), .ZN(n567) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  NAND2_X1 U627 ( .A1(n649), .A2(G56), .ZN(n568) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(n568), .Z(n574) );
  NAND2_X1 U629 ( .A1(n646), .A2(G81), .ZN(n569) );
  XNOR2_X1 U630 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G68), .A2(n644), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT13), .B(n572), .Z(n573) );
  NOR2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U635 ( .A(n575), .B(KEYINPUT70), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G43), .A2(n645), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n971) );
  XNOR2_X1 U638 ( .A(G860), .B(KEYINPUT71), .ZN(n597) );
  OR2_X1 U639 ( .A1(n971), .A2(n597), .ZN(G153) );
  NAND2_X1 U640 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U641 ( .A1(G79), .A2(n644), .ZN(n584) );
  NAND2_X1 U642 ( .A1(G66), .A2(n649), .ZN(n579) );
  NAND2_X1 U643 ( .A1(G92), .A2(n646), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n645), .A2(G54), .ZN(n580) );
  XOR2_X1 U646 ( .A(KEYINPUT72), .B(n580), .Z(n581) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT15), .ZN(n900) );
  INV_X1 U650 ( .A(n900), .ZN(n956) );
  INV_X1 U651 ( .A(G868), .ZN(n664) );
  NAND2_X1 U652 ( .A1(n956), .A2(n664), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U654 ( .A1(G53), .A2(n645), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G65), .A2(n649), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U657 ( .A1(G91), .A2(n646), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G78), .A2(n644), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n961) );
  INV_X1 U661 ( .A(n961), .ZN(G299) );
  NOR2_X1 U662 ( .A1(G286), .A2(n664), .ZN(n595) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U665 ( .A(KEYINPUT78), .B(n596), .ZN(G297) );
  NAND2_X1 U666 ( .A1(n597), .A2(G559), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n598), .A2(n900), .ZN(n599) );
  XNOR2_X1 U668 ( .A(n599), .B(KEYINPUT16), .ZN(n600) );
  XOR2_X1 U669 ( .A(KEYINPUT79), .B(n600), .Z(G148) );
  NOR2_X1 U670 ( .A1(G868), .A2(n971), .ZN(n603) );
  NAND2_X1 U671 ( .A1(G868), .A2(n900), .ZN(n601) );
  NOR2_X1 U672 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U673 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U674 ( .A1(n881), .A2(G123), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n604), .B(KEYINPUT18), .ZN(n606) );
  NAND2_X1 U676 ( .A1(G111), .A2(n882), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G135), .A2(n877), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G99), .A2(n878), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n993) );
  XNOR2_X1 U682 ( .A(n993), .B(G2096), .ZN(n612) );
  INV_X1 U683 ( .A(G2100), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(G156) );
  NAND2_X1 U685 ( .A1(n645), .A2(G50), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n613), .B(KEYINPUT84), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G62), .A2(n649), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U689 ( .A(KEYINPUT85), .B(n616), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G88), .A2(n646), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G75), .A2(n644), .ZN(n617) );
  AND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(G303) );
  INV_X1 U694 ( .A(G303), .ZN(G166) );
  NAND2_X1 U695 ( .A1(G61), .A2(n649), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G86), .A2(n646), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n644), .A2(G73), .ZN(n623) );
  XOR2_X1 U699 ( .A(KEYINPUT2), .B(n623), .Z(n624) );
  NOR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n645), .A2(G48), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(G305) );
  NAND2_X1 U703 ( .A1(n628), .A2(G87), .ZN(n633) );
  NAND2_X1 U704 ( .A1(G49), .A2(n645), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U707 ( .A1(n649), .A2(n631), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U709 ( .A(KEYINPUT83), .B(n634), .Z(G288) );
  NAND2_X1 U710 ( .A1(n645), .A2(G47), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(KEYINPUT68), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G60), .A2(n649), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U714 ( .A(KEYINPUT69), .B(n638), .ZN(n642) );
  NAND2_X1 U715 ( .A1(G85), .A2(n646), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G72), .A2(n644), .ZN(n639) );
  AND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n642), .A2(n641), .ZN(G290) );
  NAND2_X1 U719 ( .A1(G559), .A2(n900), .ZN(n643) );
  XOR2_X1 U720 ( .A(n971), .B(n643), .Z(n829) );
  XOR2_X1 U721 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n657) );
  NAND2_X1 U722 ( .A1(G80), .A2(n644), .ZN(n654) );
  NAND2_X1 U723 ( .A1(G55), .A2(n645), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G93), .A2(n646), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U726 ( .A1(G67), .A2(n649), .ZN(n650) );
  XNOR2_X1 U727 ( .A(KEYINPUT81), .B(n650), .ZN(n651) );
  NOR2_X1 U728 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U729 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n655), .B(KEYINPUT82), .ZN(n832) );
  XNOR2_X1 U731 ( .A(KEYINPUT87), .B(n832), .ZN(n656) );
  XNOR2_X1 U732 ( .A(n657), .B(n656), .ZN(n660) );
  XNOR2_X1 U733 ( .A(G166), .B(G305), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n658), .B(G288), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n660), .B(n659), .ZN(n662) );
  XNOR2_X1 U736 ( .A(G290), .B(n961), .ZN(n661) );
  XNOR2_X1 U737 ( .A(n662), .B(n661), .ZN(n899) );
  XNOR2_X1 U738 ( .A(n829), .B(n899), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n663), .A2(G868), .ZN(n666) );
  NAND2_X1 U740 ( .A1(n664), .A2(n832), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2084), .A2(G2078), .ZN(n667) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U746 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U748 ( .A1(G69), .A2(G120), .ZN(n671) );
  XNOR2_X1 U749 ( .A(KEYINPUT88), .B(n671), .ZN(n672) );
  NOR2_X1 U750 ( .A1(G238), .A2(n672), .ZN(n673) );
  NAND2_X1 U751 ( .A1(G57), .A2(n673), .ZN(n833) );
  NAND2_X1 U752 ( .A1(G567), .A2(n833), .ZN(n678) );
  NOR2_X1 U753 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U755 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U756 ( .A1(G96), .A2(n676), .ZN(n834) );
  NAND2_X1 U757 ( .A1(G2106), .A2(n834), .ZN(n677) );
  NAND2_X1 U758 ( .A1(n678), .A2(n677), .ZN(n854) );
  NAND2_X1 U759 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U760 ( .A1(n854), .A2(n679), .ZN(n828) );
  NAND2_X1 U761 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U762 ( .A1(G138), .A2(n877), .ZN(n681) );
  NAND2_X1 U763 ( .A1(G102), .A2(n878), .ZN(n680) );
  NAND2_X1 U764 ( .A1(n681), .A2(n680), .ZN(n685) );
  NAND2_X1 U765 ( .A1(G126), .A2(n881), .ZN(n683) );
  NAND2_X1 U766 ( .A1(G114), .A2(n882), .ZN(n682) );
  NAND2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U768 ( .A1(n685), .A2(n684), .ZN(G164) );
  NAND2_X1 U769 ( .A1(G40), .A2(G160), .ZN(n790) );
  INV_X1 U770 ( .A(n790), .ZN(n686) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n791) );
  NAND2_X1 U772 ( .A1(n686), .A2(n791), .ZN(n727) );
  XOR2_X1 U773 ( .A(G1996), .B(KEYINPUT97), .Z(n913) );
  NAND2_X1 U774 ( .A1(n714), .A2(n913), .ZN(n687) );
  XNOR2_X1 U775 ( .A(n687), .B(KEYINPUT26), .ZN(n688) );
  INV_X1 U776 ( .A(G1341), .ZN(n938) );
  NAND2_X1 U777 ( .A1(n688), .A2(n515), .ZN(n689) );
  NOR2_X1 U778 ( .A1(n971), .A2(n689), .ZN(n691) );
  XNOR2_X1 U779 ( .A(n691), .B(n690), .ZN(n695) );
  AND2_X1 U780 ( .A1(n727), .A2(G1348), .ZN(n693) );
  XNOR2_X1 U781 ( .A(KEYINPUT95), .B(n727), .ZN(n700) );
  AND2_X1 U782 ( .A1(n700), .A2(G2067), .ZN(n692) );
  NOR2_X1 U783 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n900), .A2(n696), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n698) );
  OR2_X1 U786 ( .A1(n900), .A2(n696), .ZN(n697) );
  NAND2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n705) );
  NAND2_X1 U788 ( .A1(n700), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U789 ( .A(n699), .B(KEYINPUT27), .ZN(n703) );
  INV_X1 U790 ( .A(G1956), .ZN(n701) );
  BUF_X1 U791 ( .A(n700), .Z(n712) );
  NOR2_X1 U792 ( .A1(n701), .A2(n712), .ZN(n702) );
  NOR2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U794 ( .A1(n961), .A2(n706), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n709) );
  OR2_X1 U796 ( .A1(n961), .A2(n706), .ZN(n707) );
  XNOR2_X1 U797 ( .A(n707), .B(KEYINPUT28), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n711) );
  INV_X1 U799 ( .A(KEYINPUT29), .ZN(n710) );
  XNOR2_X1 U800 ( .A(n711), .B(n710), .ZN(n718) );
  XNOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .ZN(n912) );
  NAND2_X1 U802 ( .A1(n712), .A2(n912), .ZN(n713) );
  XNOR2_X1 U803 ( .A(n713), .B(KEYINPUT96), .ZN(n716) );
  OR2_X1 U804 ( .A1(G1961), .A2(n714), .ZN(n715) );
  NAND2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U806 ( .A1(n719), .A2(G171), .ZN(n717) );
  NAND2_X1 U807 ( .A1(n718), .A2(n717), .ZN(n741) );
  NOR2_X1 U808 ( .A1(G171), .A2(n719), .ZN(n724) );
  NAND2_X1 U809 ( .A1(G8), .A2(n727), .ZN(n770) );
  NOR2_X1 U810 ( .A1(G1966), .A2(n770), .ZN(n743) );
  NOR2_X1 U811 ( .A1(G2084), .A2(n727), .ZN(n739) );
  NOR2_X1 U812 ( .A1(n743), .A2(n739), .ZN(n720) );
  NAND2_X1 U813 ( .A1(G8), .A2(n720), .ZN(n721) );
  XNOR2_X1 U814 ( .A(KEYINPUT30), .B(n721), .ZN(n722) );
  NOR2_X1 U815 ( .A1(G168), .A2(n722), .ZN(n723) );
  NOR2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n726) );
  XOR2_X1 U817 ( .A(KEYINPUT31), .B(KEYINPUT98), .Z(n725) );
  XNOR2_X1 U818 ( .A(n726), .B(n725), .ZN(n740) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n770), .ZN(n729) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U822 ( .A1(n730), .A2(G303), .ZN(n732) );
  AND2_X1 U823 ( .A1(n740), .A2(n732), .ZN(n731) );
  NAND2_X1 U824 ( .A1(n741), .A2(n731), .ZN(n737) );
  INV_X1 U825 ( .A(n732), .ZN(n733) );
  NOR2_X1 U826 ( .A1(n733), .A2(G286), .ZN(n735) );
  INV_X1 U827 ( .A(G8), .ZN(n734) );
  NOR2_X1 U828 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U830 ( .A(n738), .B(KEYINPUT32), .ZN(n747) );
  NAND2_X1 U831 ( .A1(G8), .A2(n739), .ZN(n745) );
  AND2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n762) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n753) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n753), .A2(n748), .ZN(n960) );
  NAND2_X1 U839 ( .A1(n762), .A2(n960), .ZN(n749) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n959) );
  NAND2_X1 U841 ( .A1(n749), .A2(n959), .ZN(n750) );
  NOR2_X1 U842 ( .A1(KEYINPUT33), .A2(n750), .ZN(n751) );
  INV_X1 U843 ( .A(n770), .ZN(n752) );
  NAND2_X1 U844 ( .A1(n751), .A2(n752), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U846 ( .A1(n754), .A2(KEYINPUT33), .ZN(n755) );
  NAND2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n758) );
  XNOR2_X1 U848 ( .A(n758), .B(n757), .ZN(n759) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n975) );
  NAND2_X1 U850 ( .A1(n759), .A2(n975), .ZN(n766) );
  NOR2_X1 U851 ( .A1(G2090), .A2(G303), .ZN(n760) );
  XNOR2_X1 U852 ( .A(n760), .B(KEYINPUT100), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n761), .A2(G8), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U855 ( .A1(n764), .A2(n770), .ZN(n765) );
  NAND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n772) );
  NOR2_X1 U857 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XOR2_X1 U858 ( .A(n767), .B(KEYINPUT24), .Z(n768) );
  XNOR2_X1 U859 ( .A(KEYINPUT94), .B(n768), .ZN(n769) );
  NOR2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n877), .A2(G131), .ZN(n773) );
  XOR2_X1 U862 ( .A(KEYINPUT91), .B(n773), .Z(n775) );
  NAND2_X1 U863 ( .A1(n878), .A2(G95), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U865 ( .A(KEYINPUT92), .B(n776), .Z(n780) );
  NAND2_X1 U866 ( .A1(G119), .A2(n881), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G107), .A2(n882), .ZN(n777) );
  AND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n892) );
  AND2_X1 U870 ( .A1(n892), .A2(G1991), .ZN(n789) );
  NAND2_X1 U871 ( .A1(G141), .A2(n877), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G129), .A2(n881), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n878), .A2(G105), .ZN(n783) );
  XOR2_X1 U875 ( .A(KEYINPUT38), .B(n783), .Z(n784) );
  NOR2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n882), .A2(G117), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n893) );
  AND2_X1 U879 ( .A1(n893), .A2(G1996), .ZN(n788) );
  NOR2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n1004) );
  NOR2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U882 ( .A(KEYINPUT89), .B(n792), .Z(n818) );
  INV_X1 U883 ( .A(n818), .ZN(n793) );
  NOR2_X1 U884 ( .A1(n1004), .A2(n793), .ZN(n810) );
  INV_X1 U885 ( .A(n810), .ZN(n804) );
  NAND2_X1 U886 ( .A1(G140), .A2(n877), .ZN(n795) );
  NAND2_X1 U887 ( .A1(G104), .A2(n878), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n796), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G128), .A2(n881), .ZN(n798) );
  NAND2_X1 U891 ( .A1(G116), .A2(n882), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U893 ( .A(KEYINPUT35), .B(n799), .Z(n800) );
  XNOR2_X1 U894 ( .A(KEYINPUT90), .B(n800), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U896 ( .A(KEYINPUT36), .B(n803), .ZN(n896) );
  XNOR2_X1 U897 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  NOR2_X1 U898 ( .A1(n896), .A2(n816), .ZN(n985) );
  NAND2_X1 U899 ( .A1(n818), .A2(n985), .ZN(n814) );
  NAND2_X1 U900 ( .A1(n804), .A2(n814), .ZN(n805) );
  XOR2_X1 U901 ( .A(KEYINPUT93), .B(n805), .Z(n806) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n968) );
  NAND2_X1 U903 ( .A1(n807), .A2(n517), .ZN(n821) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n893), .ZN(n1001) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n892), .ZN(n997) );
  NOR2_X1 U907 ( .A1(n808), .A2(n997), .ZN(n809) );
  NOR2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U909 ( .A1(n1001), .A2(n811), .ZN(n813) );
  XOR2_X1 U910 ( .A(KEYINPUT39), .B(KEYINPUT101), .Z(n812) );
  XNOR2_X1 U911 ( .A(n813), .B(n812), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n896), .A2(n816), .ZN(n984) );
  NAND2_X1 U914 ( .A1(n817), .A2(n984), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U917 ( .A(KEYINPUT40), .B(n822), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n823), .ZN(G217) );
  INV_X1 U919 ( .A(G661), .ZN(n825) );
  NAND2_X1 U920 ( .A1(G2), .A2(G15), .ZN(n824) );
  NOR2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U922 ( .A(KEYINPUT104), .B(n826), .Z(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U924 ( .A1(n828), .A2(n827), .ZN(G188) );
  XNOR2_X1 U925 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  XOR2_X1 U927 ( .A(n829), .B(KEYINPUT80), .Z(n830) );
  NOR2_X1 U928 ( .A1(G860), .A2(n830), .ZN(n831) );
  XOR2_X1 U929 ( .A(n832), .B(n831), .Z(G145) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G69), .ZN(G235) );
  NOR2_X1 U932 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XOR2_X1 U934 ( .A(KEYINPUT43), .B(G2678), .Z(n836) );
  XNOR2_X1 U935 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U937 ( .A(KEYINPUT42), .B(G2090), .Z(n838) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U940 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2096), .B(G2100), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n844) );
  XOR2_X1 U943 ( .A(G2084), .B(G2078), .Z(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1956), .B(G1961), .Z(n846) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1966), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U948 ( .A(n847), .B(G2474), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1971), .B(G1976), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1981), .Z(n851) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U955 ( .A(KEYINPUT106), .B(n854), .Z(G319) );
  NAND2_X1 U956 ( .A1(G112), .A2(n882), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G136), .A2(n877), .ZN(n856) );
  NAND2_X1 U958 ( .A1(G100), .A2(n878), .ZN(n855) );
  NAND2_X1 U959 ( .A1(n856), .A2(n855), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n881), .A2(G124), .ZN(n857) );
  XOR2_X1 U961 ( .A(KEYINPUT44), .B(n857), .Z(n858) );
  NOR2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n862), .B(KEYINPUT109), .ZN(G162) );
  XOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n864) );
  XNOR2_X1 U966 ( .A(G164), .B(KEYINPUT112), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n993), .B(n865), .ZN(n867) );
  XNOR2_X1 U969 ( .A(G160), .B(G162), .ZN(n866) );
  XNOR2_X1 U970 ( .A(n867), .B(n866), .ZN(n891) );
  NAND2_X1 U971 ( .A1(n878), .A2(G106), .ZN(n868) );
  XOR2_X1 U972 ( .A(KEYINPUT111), .B(n868), .Z(n870) );
  NAND2_X1 U973 ( .A1(n877), .A2(G142), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U975 ( .A(n871), .B(KEYINPUT45), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G130), .A2(n881), .ZN(n873) );
  NAND2_X1 U977 ( .A1(G118), .A2(n882), .ZN(n872) );
  NAND2_X1 U978 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U979 ( .A(KEYINPUT110), .B(n874), .Z(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n889) );
  NAND2_X1 U981 ( .A1(G139), .A2(n877), .ZN(n880) );
  NAND2_X1 U982 ( .A1(G103), .A2(n878), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G127), .A2(n881), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G115), .A2(n882), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U987 ( .A(KEYINPUT47), .B(n885), .ZN(n886) );
  XNOR2_X1 U988 ( .A(KEYINPUT113), .B(n886), .ZN(n887) );
  NOR2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n987) );
  XNOR2_X1 U990 ( .A(n889), .B(n987), .ZN(n890) );
  XOR2_X1 U991 ( .A(n891), .B(n890), .Z(n895) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U994 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U995 ( .A1(G37), .A2(n898), .ZN(G395) );
  XOR2_X1 U996 ( .A(n899), .B(G286), .Z(n902) );
  XNOR2_X1 U997 ( .A(G171), .B(n900), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U999 ( .A(n903), .B(n971), .Z(n904) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n904), .ZN(G397) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n905) );
  XOR2_X1 U1002 ( .A(KEYINPUT49), .B(n905), .Z(n906) );
  NAND2_X1 U1003 ( .A1(n906), .A2(G319), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(G401), .A2(n907), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(KEYINPUT114), .B(n908), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1010 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n1026) );
  XOR2_X1 U1011 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n1008) );
  XOR2_X1 U1012 ( .A(n1008), .B(KEYINPUT118), .Z(n930) );
  XNOR2_X1 U1013 ( .A(G2090), .B(G35), .ZN(n925) );
  XOR2_X1 U1014 ( .A(G25), .B(G1991), .Z(n911) );
  NAND2_X1 U1015 ( .A1(n911), .A2(G28), .ZN(n922) );
  XNOR2_X1 U1016 ( .A(G27), .B(n912), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n913), .B(G32), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(G2067), .B(G26), .ZN(n915) );
  XNOR2_X1 U1019 ( .A(G2072), .B(G33), .ZN(n914) );
  NOR2_X1 U1020 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1021 ( .A(KEYINPUT117), .B(n916), .ZN(n917) );
  NOR2_X1 U1022 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1023 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1025 ( .A(KEYINPUT53), .B(n923), .ZN(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n928) );
  XOR2_X1 U1027 ( .A(G2084), .B(G34), .Z(n926) );
  XNOR2_X1 U1028 ( .A(KEYINPUT54), .B(n926), .ZN(n927) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n930), .B(n929), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(G29), .A2(n931), .ZN(n1024) );
  XOR2_X1 U1032 ( .A(G1986), .B(G24), .Z(n935) );
  XNOR2_X1 U1033 ( .A(G1971), .B(G22), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(G23), .B(G1976), .ZN(n932) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(n937), .B(n936), .ZN(n953) );
  XNOR2_X1 U1039 ( .A(G19), .B(n938), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G1956), .B(G20), .ZN(n940) );
  XNOR2_X1 U1041 ( .A(G6), .B(G1981), .ZN(n939) );
  NOR2_X1 U1042 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1044 ( .A(KEYINPUT59), .B(G1348), .Z(n943) );
  XNOR2_X1 U1045 ( .A(G4), .B(n943), .ZN(n944) );
  NOR2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1047 ( .A(KEYINPUT60), .B(n946), .ZN(n948) );
  XOR2_X1 U1048 ( .A(G1961), .B(G5), .Z(n947) );
  NAND2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(G21), .B(G1966), .ZN(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(KEYINPUT124), .B(n951), .ZN(n952) );
  NAND2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1054 ( .A(KEYINPUT61), .B(n954), .ZN(n1013) );
  NOR2_X1 U1055 ( .A1(KEYINPUT123), .A2(n1013), .ZN(n982) );
  XNOR2_X1 U1056 ( .A(G171), .B(KEYINPUT120), .ZN(n955) );
  XOR2_X1 U1057 ( .A(n955), .B(G1961), .Z(n958) );
  XNOR2_X1 U1058 ( .A(G1348), .B(n956), .ZN(n957) );
  NOR2_X1 U1059 ( .A1(n958), .A2(n957), .ZN(n970) );
  NAND2_X1 U1060 ( .A1(n960), .A2(n959), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(n961), .B(G1956), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(G1971), .A2(G303), .ZN(n962) );
  NAND2_X1 U1063 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1065 ( .A(KEYINPUT121), .B(n966), .ZN(n967) );
  NOR2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(G1341), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1070 ( .A(KEYINPUT122), .B(n974), .Z(n980) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G168), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(n977), .B(KEYINPUT119), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(KEYINPUT57), .B(n978), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n1011) );
  NOR2_X1 U1076 ( .A1(KEYINPUT56), .A2(n1011), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(G16), .A2(n983), .ZN(n1021) );
  INV_X1 U1079 ( .A(n984), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n999) );
  XNOR2_X1 U1081 ( .A(G2084), .B(G160), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(n987), .B(G2072), .ZN(n990) );
  XOR2_X1 U1083 ( .A(G164), .B(G2078), .Z(n988) );
  XNOR2_X1 U1084 ( .A(KEYINPUT115), .B(n988), .ZN(n989) );
  NAND2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1086 ( .A(KEYINPUT50), .B(n991), .ZN(n992) );
  NOR2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1006) );
  XOR2_X1 U1091 ( .A(G2090), .B(G162), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1093 ( .A(KEYINPUT51), .B(n1002), .Z(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT52), .B(n1007), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(G29), .A2(n1010), .ZN(n1019) );
  INV_X1 U1099 ( .A(n1011), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(KEYINPUT56), .A2(n1012), .ZN(n1016) );
  INV_X1 U1101 ( .A(n1013), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(KEYINPUT123), .A2(n1014), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(G16), .A2(n1017), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(G11), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(n1026), .B(n1025), .ZN(n1027) );
  XNOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1027), .ZN(G150) );
  INV_X1 U1111 ( .A(G150), .ZN(G311) );
endmodule

