

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U558 ( .A1(n636), .A2(n542), .ZN(n655) );
  NOR2_X1 U559 ( .A1(G543), .A2(G651), .ZN(n650) );
  AND2_X1 U560 ( .A1(n816), .A2(n832), .ZN(n524) );
  NOR2_X1 U561 ( .A1(n782), .A2(n772), .ZN(n525) );
  NOR2_X1 U562 ( .A1(n703), .A2(n702), .ZN(n705) );
  XNOR2_X1 U563 ( .A(n725), .B(KEYINPUT97), .ZN(n726) );
  XNOR2_X1 U564 ( .A(n727), .B(n726), .ZN(n728) );
  AND2_X1 U565 ( .A1(n797), .A2(n690), .ZN(n706) );
  INV_X1 U566 ( .A(n706), .ZN(n736) );
  INV_X1 U567 ( .A(KEYINPUT88), .ZN(n550) );
  NOR2_X1 U568 ( .A1(n817), .A2(n524), .ZN(n818) );
  NOR2_X1 U569 ( .A1(n636), .A2(G651), .ZN(n659) );
  NOR2_X1 U570 ( .A1(n575), .A2(n574), .ZN(n1000) );
  NOR2_X1 U571 ( .A1(n536), .A2(n535), .ZN(G160) );
  NOR2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  XNOR2_X1 U573 ( .A(n526), .B(KEYINPUT65), .ZN(n528) );
  XNOR2_X1 U574 ( .A(KEYINPUT66), .B(KEYINPUT17), .ZN(n527) );
  XNOR2_X1 U575 ( .A(n528), .B(n527), .ZN(n547) );
  NAND2_X1 U576 ( .A1(G137), .A2(n547), .ZN(n531) );
  INV_X1 U577 ( .A(G2105), .ZN(n532) );
  AND2_X1 U578 ( .A1(n532), .A2(G2104), .ZN(n879) );
  NAND2_X1 U579 ( .A1(G101), .A2(n879), .ZN(n529) );
  XOR2_X1 U580 ( .A(KEYINPUT23), .B(n529), .Z(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n536) );
  AND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n884) );
  NAND2_X1 U583 ( .A1(G113), .A2(n884), .ZN(n534) );
  NOR2_X1 U584 ( .A1(G2104), .A2(n532), .ZN(n882) );
  NAND2_X1 U585 ( .A1(G125), .A2(n882), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n636) );
  NAND2_X1 U588 ( .A1(n659), .A2(G47), .ZN(n541) );
  INV_X1 U589 ( .A(G651), .ZN(n542) );
  NOR2_X1 U590 ( .A1(G543), .A2(n542), .ZN(n538) );
  XNOR2_X1 U591 ( .A(KEYINPUT68), .B(KEYINPUT1), .ZN(n537) );
  XNOR2_X1 U592 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U593 ( .A(KEYINPUT67), .B(n539), .ZN(n651) );
  NAND2_X1 U594 ( .A1(G60), .A2(n651), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n546) );
  NAND2_X1 U596 ( .A1(G85), .A2(n650), .ZN(n544) );
  NAND2_X1 U597 ( .A1(G72), .A2(n655), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U599 ( .A1(n546), .A2(n545), .ZN(G290) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U601 ( .A(G57), .ZN(G237) );
  INV_X1 U602 ( .A(G132), .ZN(G219) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  NAND2_X1 U604 ( .A1(G138), .A2(n547), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n879), .A2(G102), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U607 ( .A(n551), .B(n550), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n882), .A2(G126), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n553), .A2(n552), .ZN(n556) );
  NAND2_X1 U610 ( .A1(G114), .A2(n884), .ZN(n554) );
  XNOR2_X1 U611 ( .A(KEYINPUT87), .B(n554), .ZN(n555) );
  NOR2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n689) );
  BUF_X1 U613 ( .A(n689), .Z(G164) );
  NAND2_X1 U614 ( .A1(n659), .A2(G52), .ZN(n558) );
  NAND2_X1 U615 ( .A1(G64), .A2(n651), .ZN(n557) );
  NAND2_X1 U616 ( .A1(n558), .A2(n557), .ZN(n563) );
  NAND2_X1 U617 ( .A1(G90), .A2(n650), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G77), .A2(n655), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U621 ( .A1(n563), .A2(n562), .ZN(G171) );
  NAND2_X1 U622 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U623 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U624 ( .A(G223), .ZN(n837) );
  NAND2_X1 U625 ( .A1(n837), .A2(G567), .ZN(n565) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(n565), .Z(G234) );
  NAND2_X1 U627 ( .A1(G56), .A2(n651), .ZN(n566) );
  XNOR2_X1 U628 ( .A(n566), .B(KEYINPUT14), .ZN(n568) );
  NAND2_X1 U629 ( .A1(G43), .A2(n659), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n575) );
  NAND2_X1 U631 ( .A1(G68), .A2(n655), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n650), .A2(G81), .ZN(n569) );
  XNOR2_X1 U633 ( .A(n569), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(KEYINPUT13), .ZN(n573) );
  XNOR2_X1 U636 ( .A(KEYINPUT69), .B(n573), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n1000), .A2(G860), .ZN(G153) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(n659), .A2(G54), .ZN(n582) );
  NAND2_X1 U640 ( .A1(G92), .A2(n650), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G79), .A2(n655), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n651), .A2(G66), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT70), .B(n578), .Z(n579) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT15), .B(n583), .Z(n712) );
  INV_X1 U648 ( .A(n712), .ZN(n988) );
  NOR2_X1 U649 ( .A1(n988), .A2(G868), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n584), .B(KEYINPUT71), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U653 ( .A1(G76), .A2(n655), .ZN(n591) );
  XOR2_X1 U654 ( .A(KEYINPUT4), .B(KEYINPUT73), .Z(n588) );
  NAND2_X1 U655 ( .A1(G89), .A2(n650), .ZN(n587) );
  XNOR2_X1 U656 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U657 ( .A(KEYINPUT72), .B(n589), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U659 ( .A(n592), .B(KEYINPUT74), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n593), .B(KEYINPUT5), .ZN(n598) );
  NAND2_X1 U661 ( .A1(n659), .A2(G51), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G63), .A2(n651), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U664 ( .A(KEYINPUT6), .B(n596), .Z(n597) );
  NAND2_X1 U665 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U666 ( .A(n599), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U667 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U668 ( .A1(n659), .A2(G53), .ZN(n601) );
  NAND2_X1 U669 ( .A1(G65), .A2(n651), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U671 ( .A1(G91), .A2(n650), .ZN(n603) );
  NAND2_X1 U672 ( .A1(G78), .A2(n655), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n985) );
  INV_X1 U675 ( .A(n985), .ZN(G299) );
  INV_X1 U676 ( .A(G868), .ZN(n611) );
  NOR2_X1 U677 ( .A1(G286), .A2(n611), .ZN(n607) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n606) );
  NOR2_X1 U679 ( .A1(n607), .A2(n606), .ZN(G297) );
  INV_X1 U680 ( .A(G559), .ZN(n612) );
  NOR2_X1 U681 ( .A1(G860), .A2(n612), .ZN(n608) );
  XNOR2_X1 U682 ( .A(KEYINPUT75), .B(n608), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n609), .A2(n988), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  AND2_X1 U685 ( .A1(n611), .A2(n1000), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G868), .A2(n612), .ZN(n613) );
  NOR2_X1 U687 ( .A1(n613), .A2(n712), .ZN(n614) );
  NOR2_X1 U688 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U689 ( .A1(n882), .A2(G123), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n616), .B(KEYINPUT18), .ZN(n618) );
  BUF_X1 U691 ( .A(n547), .Z(n889) );
  NAND2_X1 U692 ( .A1(G135), .A2(n889), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U694 ( .A(KEYINPUT76), .B(n619), .ZN(n623) );
  NAND2_X1 U695 ( .A1(G99), .A2(n879), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G111), .A2(n884), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n928) );
  XNOR2_X1 U699 ( .A(n928), .B(G2096), .ZN(n625) );
  INV_X1 U700 ( .A(G2100), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(G156) );
  XOR2_X1 U702 ( .A(n1000), .B(KEYINPUT77), .Z(n627) );
  NAND2_X1 U703 ( .A1(G559), .A2(n988), .ZN(n626) );
  XOR2_X1 U704 ( .A(n627), .B(n626), .Z(n670) );
  NOR2_X1 U705 ( .A1(n670), .A2(G860), .ZN(n635) );
  NAND2_X1 U706 ( .A1(G93), .A2(n650), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G80), .A2(n655), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G55), .A2(n659), .ZN(n630) );
  XNOR2_X1 U710 ( .A(n630), .B(KEYINPUT78), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G67), .A2(n651), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n664) );
  XNOR2_X1 U714 ( .A(n635), .B(n664), .ZN(G145) );
  NAND2_X1 U715 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G87), .A2(n636), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U718 ( .A1(n651), .A2(n639), .ZN(n642) );
  NAND2_X1 U719 ( .A1(G49), .A2(n659), .ZN(n640) );
  XOR2_X1 U720 ( .A(KEYINPUT79), .B(n640), .Z(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U722 ( .A1(n659), .A2(G50), .ZN(n644) );
  NAND2_X1 U723 ( .A1(G62), .A2(n651), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G75), .A2(n655), .ZN(n645) );
  XNOR2_X1 U726 ( .A(KEYINPUT81), .B(n645), .ZN(n646) );
  NOR2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n650), .A2(G88), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(G303) );
  INV_X1 U730 ( .A(G303), .ZN(G166) );
  NAND2_X1 U731 ( .A1(n650), .A2(G86), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G61), .A2(n651), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U734 ( .A(KEYINPUT80), .B(n654), .ZN(n658) );
  NAND2_X1 U735 ( .A1(n655), .A2(G73), .ZN(n656) );
  XOR2_X1 U736 ( .A(KEYINPUT2), .B(n656), .Z(n657) );
  NOR2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U738 ( .A1(n659), .A2(G48), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(G305) );
  NOR2_X1 U740 ( .A1(G868), .A2(n664), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n662), .B(KEYINPUT83), .ZN(n673) );
  XNOR2_X1 U742 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n663) );
  XNOR2_X1 U743 ( .A(n663), .B(G288), .ZN(n669) );
  XNOR2_X1 U744 ( .A(G166), .B(n664), .ZN(n666) );
  XNOR2_X1 U745 ( .A(G290), .B(n985), .ZN(n665) );
  XNOR2_X1 U746 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U747 ( .A(n667), .B(G305), .Z(n668) );
  XNOR2_X1 U748 ( .A(n669), .B(n668), .ZN(n910) );
  XOR2_X1 U749 ( .A(n670), .B(n910), .Z(n671) );
  NAND2_X1 U750 ( .A1(G868), .A2(n671), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U754 ( .A1(n675), .A2(G2090), .ZN(n676) );
  XNOR2_X1 U755 ( .A(n676), .B(KEYINPUT84), .ZN(n677) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U757 ( .A1(G2072), .A2(n678), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U759 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n679) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n679), .Z(n680) );
  NOR2_X1 U762 ( .A1(G218), .A2(n680), .ZN(n681) );
  XOR2_X1 U763 ( .A(KEYINPUT85), .B(n681), .Z(n682) );
  NAND2_X1 U764 ( .A1(G96), .A2(n682), .ZN(n841) );
  NAND2_X1 U765 ( .A1(n841), .A2(G2106), .ZN(n686) );
  NAND2_X1 U766 ( .A1(G69), .A2(G120), .ZN(n683) );
  NOR2_X1 U767 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U768 ( .A1(G108), .A2(n684), .ZN(n842) );
  NAND2_X1 U769 ( .A1(n842), .A2(G567), .ZN(n685) );
  NAND2_X1 U770 ( .A1(n686), .A2(n685), .ZN(n843) );
  NOR2_X1 U771 ( .A1(n687), .A2(n843), .ZN(n688) );
  XNOR2_X1 U772 ( .A(n688), .B(KEYINPUT86), .ZN(n840) );
  NAND2_X1 U773 ( .A1(G36), .A2(n840), .ZN(G176) );
  NOR2_X1 U774 ( .A1(n689), .A2(G1384), .ZN(n797) );
  NAND2_X1 U775 ( .A1(G160), .A2(G40), .ZN(n796) );
  INV_X1 U776 ( .A(n796), .ZN(n690) );
  INV_X1 U777 ( .A(G1961), .ZN(n1009) );
  NAND2_X1 U778 ( .A1(n736), .A2(n1009), .ZN(n692) );
  XNOR2_X1 U779 ( .A(G2078), .B(KEYINPUT25), .ZN(n957) );
  NAND2_X1 U780 ( .A1(n706), .A2(n957), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n692), .A2(n691), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n729), .A2(G171), .ZN(n723) );
  NAND2_X1 U783 ( .A1(G2072), .A2(n706), .ZN(n693) );
  XOR2_X1 U784 ( .A(KEYINPUT93), .B(n693), .Z(n694) );
  XNOR2_X1 U785 ( .A(KEYINPUT27), .B(n694), .ZN(n696) );
  INV_X1 U786 ( .A(G1956), .ZN(n1015) );
  NOR2_X1 U787 ( .A1(n706), .A2(n1015), .ZN(n695) );
  NOR2_X1 U788 ( .A1(n696), .A2(n695), .ZN(n716) );
  NOR2_X1 U789 ( .A1(n985), .A2(n716), .ZN(n697) );
  XOR2_X1 U790 ( .A(n697), .B(KEYINPUT28), .Z(n720) );
  INV_X1 U791 ( .A(G1341), .ZN(n698) );
  OR2_X1 U792 ( .A1(n706), .A2(n698), .ZN(n699) );
  XNOR2_X1 U793 ( .A(n699), .B(KEYINPUT94), .ZN(n700) );
  NAND2_X1 U794 ( .A1(n700), .A2(n1000), .ZN(n703) );
  NAND2_X1 U795 ( .A1(G1996), .A2(n706), .ZN(n701) );
  XOR2_X1 U796 ( .A(KEYINPUT26), .B(n701), .Z(n702) );
  INV_X1 U797 ( .A(KEYINPUT64), .ZN(n704) );
  XNOR2_X1 U798 ( .A(n705), .B(n704), .ZN(n713) );
  OR2_X1 U799 ( .A1(n712), .A2(n713), .ZN(n711) );
  AND2_X1 U800 ( .A1(n706), .A2(G2067), .ZN(n707) );
  XNOR2_X1 U801 ( .A(n707), .B(KEYINPUT95), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n736), .A2(G1348), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U804 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U805 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n985), .A2(n716), .ZN(n717) );
  NAND2_X1 U808 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U809 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U810 ( .A(KEYINPUT29), .B(n721), .Z(n722) );
  NAND2_X1 U811 ( .A1(n723), .A2(n722), .ZN(n734) );
  NAND2_X1 U812 ( .A1(G8), .A2(n736), .ZN(n782) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n782), .ZN(n747) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n736), .ZN(n744) );
  NOR2_X1 U815 ( .A1(n747), .A2(n744), .ZN(n724) );
  NAND2_X1 U816 ( .A1(G8), .A2(n724), .ZN(n727) );
  XOR2_X1 U817 ( .A(KEYINPUT30), .B(KEYINPUT96), .Z(n725) );
  NOR2_X1 U818 ( .A1(G168), .A2(n728), .ZN(n731) );
  NOR2_X1 U819 ( .A1(G171), .A2(n729), .ZN(n730) );
  NOR2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U821 ( .A(KEYINPUT31), .B(n732), .Z(n733) );
  NAND2_X1 U822 ( .A1(n734), .A2(n733), .ZN(n745) );
  NAND2_X1 U823 ( .A1(G286), .A2(n745), .ZN(n735) );
  XNOR2_X1 U824 ( .A(n735), .B(KEYINPUT98), .ZN(n741) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n782), .ZN(n738) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U828 ( .A1(n739), .A2(G303), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U830 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U831 ( .A(n743), .B(KEYINPUT32), .ZN(n766) );
  NAND2_X1 U832 ( .A1(G8), .A2(n744), .ZN(n749) );
  INV_X1 U833 ( .A(n745), .ZN(n746) );
  NOR2_X1 U834 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U835 ( .A1(n749), .A2(n748), .ZN(n757) );
  NAND2_X1 U836 ( .A1(n766), .A2(n757), .ZN(n753) );
  NOR2_X1 U837 ( .A1(G2090), .A2(G303), .ZN(n750) );
  NAND2_X1 U838 ( .A1(G8), .A2(n750), .ZN(n751) );
  XNOR2_X1 U839 ( .A(n751), .B(KEYINPUT102), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n755) );
  INV_X1 U841 ( .A(KEYINPUT103), .ZN(n754) );
  XNOR2_X1 U842 ( .A(n755), .B(n754), .ZN(n756) );
  NAND2_X1 U843 ( .A1(n756), .A2(n782), .ZN(n779) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n990) );
  AND2_X1 U845 ( .A1(n757), .A2(n990), .ZN(n759) );
  INV_X1 U846 ( .A(n782), .ZN(n758) );
  AND2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n764) );
  XOR2_X1 U848 ( .A(G1981), .B(G305), .Z(n982) );
  NOR2_X1 U849 ( .A1(G288), .A2(G1976), .ZN(n760) );
  XNOR2_X1 U850 ( .A(n760), .B(KEYINPUT99), .ZN(n767) );
  NOR2_X1 U851 ( .A1(n782), .A2(n767), .ZN(n761) );
  NAND2_X1 U852 ( .A1(KEYINPUT33), .A2(n761), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n982), .A2(n762), .ZN(n774) );
  INV_X1 U854 ( .A(n774), .ZN(n763) );
  AND2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n776) );
  INV_X1 U857 ( .A(n990), .ZN(n771) );
  INV_X1 U858 ( .A(n767), .ZN(n769) );
  NOR2_X1 U859 ( .A1(G1971), .A2(G303), .ZN(n768) );
  NOR2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n998) );
  XNOR2_X1 U861 ( .A(KEYINPUT100), .B(n998), .ZN(n770) );
  OR2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U863 ( .A1(KEYINPUT33), .A2(n525), .ZN(n773) );
  OR2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U866 ( .A(n777), .B(KEYINPUT101), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n785) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n780) );
  XOR2_X1 U869 ( .A(n780), .B(KEYINPUT24), .Z(n781) );
  XNOR2_X1 U870 ( .A(KEYINPUT92), .B(n781), .ZN(n783) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  INV_X1 U873 ( .A(n786), .ZN(n819) );
  NAND2_X1 U874 ( .A1(n879), .A2(G104), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G140), .A2(n889), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U877 ( .A(KEYINPUT34), .B(n789), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G116), .A2(n884), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G128), .A2(n882), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U881 ( .A(KEYINPUT35), .B(n792), .Z(n793) );
  NOR2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U883 ( .A(KEYINPUT36), .B(n795), .ZN(n905) );
  XNOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NOR2_X1 U885 ( .A1(n905), .A2(n820), .ZN(n932) );
  NOR2_X1 U886 ( .A1(n797), .A2(n796), .ZN(n832) );
  NAND2_X1 U887 ( .A1(n932), .A2(n832), .ZN(n798) );
  XOR2_X1 U888 ( .A(KEYINPUT89), .B(n798), .Z(n829) );
  INV_X1 U889 ( .A(n829), .ZN(n817) );
  NAND2_X1 U890 ( .A1(G129), .A2(n882), .ZN(n799) );
  XNOR2_X1 U891 ( .A(n799), .B(KEYINPUT90), .ZN(n803) );
  XOR2_X1 U892 ( .A(KEYINPUT91), .B(KEYINPUT38), .Z(n801) );
  NAND2_X1 U893 ( .A1(G105), .A2(n879), .ZN(n800) );
  XNOR2_X1 U894 ( .A(n801), .B(n800), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n807) );
  NAND2_X1 U896 ( .A1(n884), .A2(G117), .ZN(n805) );
  NAND2_X1 U897 ( .A1(G141), .A2(n889), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n899) );
  INV_X1 U900 ( .A(G1996), .ZN(n958) );
  NOR2_X1 U901 ( .A1(n899), .A2(n958), .ZN(n815) );
  NAND2_X1 U902 ( .A1(n882), .A2(G119), .ZN(n809) );
  NAND2_X1 U903 ( .A1(G131), .A2(n889), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n813) );
  NAND2_X1 U905 ( .A1(G95), .A2(n879), .ZN(n811) );
  NAND2_X1 U906 ( .A1(G107), .A2(n884), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n896) );
  INV_X1 U909 ( .A(G1991), .ZN(n955) );
  NOR2_X1 U910 ( .A1(n896), .A2(n955), .ZN(n814) );
  NOR2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n824) );
  XOR2_X1 U912 ( .A(G1986), .B(G290), .Z(n986) );
  NAND2_X1 U913 ( .A1(n824), .A2(n986), .ZN(n816) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n835) );
  NAND2_X1 U915 ( .A1(n905), .A2(n820), .ZN(n935) );
  AND2_X1 U916 ( .A1(n958), .A2(n899), .ZN(n938) );
  AND2_X1 U917 ( .A1(n955), .A2(n896), .ZN(n821) );
  XOR2_X1 U918 ( .A(KEYINPUT105), .B(n821), .Z(n929) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n822) );
  XNOR2_X1 U920 ( .A(KEYINPUT104), .B(n822), .ZN(n823) );
  NOR2_X1 U921 ( .A1(n929), .A2(n823), .ZN(n825) );
  INV_X1 U922 ( .A(n824), .ZN(n934) );
  NOR2_X1 U923 ( .A1(n825), .A2(n934), .ZN(n826) );
  NOR2_X1 U924 ( .A1(n938), .A2(n826), .ZN(n827) );
  XNOR2_X1 U925 ( .A(KEYINPUT39), .B(n827), .ZN(n828) );
  XNOR2_X1 U926 ( .A(n828), .B(KEYINPUT106), .ZN(n830) );
  NAND2_X1 U927 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n935), .A2(n831), .ZN(n833) );
  NAND2_X1 U929 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U930 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n836), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U934 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U938 ( .A(G120), .ZN(G236) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  NOR2_X1 U941 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  INV_X1 U943 ( .A(n843), .ZN(G319) );
  XOR2_X1 U944 ( .A(KEYINPUT42), .B(G2090), .Z(n845) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2084), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U947 ( .A(n846), .B(G2100), .Z(n848) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U950 ( .A(G2096), .B(KEYINPUT43), .Z(n850) );
  XNOR2_X1 U951 ( .A(G2678), .B(KEYINPUT107), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U953 ( .A(n852), .B(n851), .Z(G227) );
  XNOR2_X1 U954 ( .A(G1991), .B(G2474), .ZN(n862) );
  XOR2_X1 U955 ( .A(G1956), .B(G1961), .Z(n854) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1986), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U958 ( .A(G1976), .B(G1981), .Z(n856) );
  XNOR2_X1 U959 ( .A(G1966), .B(G1971), .ZN(n855) );
  XNOR2_X1 U960 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U961 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U962 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U965 ( .A1(G100), .A2(n879), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G112), .A2(n884), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n882), .A2(G124), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G136), .A2(n889), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U972 ( .A(KEYINPUT109), .B(n868), .Z(n869) );
  NOR2_X1 U973 ( .A1(n870), .A2(n869), .ZN(G162) );
  XNOR2_X1 U974 ( .A(G162), .B(n928), .ZN(n904) );
  NAND2_X1 U975 ( .A1(n879), .A2(G106), .ZN(n872) );
  NAND2_X1 U976 ( .A1(G142), .A2(n889), .ZN(n871) );
  NAND2_X1 U977 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U978 ( .A(n873), .B(KEYINPUT45), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G118), .A2(n884), .ZN(n875) );
  NAND2_X1 U980 ( .A1(G130), .A2(n882), .ZN(n874) );
  NAND2_X1 U981 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U982 ( .A(KEYINPUT110), .B(n876), .Z(n877) );
  NAND2_X1 U983 ( .A1(n878), .A2(n877), .ZN(n894) );
  NAND2_X1 U984 ( .A1(n879), .A2(G103), .ZN(n880) );
  XNOR2_X1 U985 ( .A(KEYINPUT111), .B(n880), .ZN(n893) );
  XOR2_X1 U986 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n881) );
  XNOR2_X1 U987 ( .A(KEYINPUT47), .B(n881), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n882), .A2(G127), .ZN(n883) );
  XNOR2_X1 U989 ( .A(n883), .B(KEYINPUT112), .ZN(n886) );
  NAND2_X1 U990 ( .A1(G115), .A2(n884), .ZN(n885) );
  NAND2_X1 U991 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U992 ( .A(n888), .B(n887), .ZN(n891) );
  NAND2_X1 U993 ( .A1(G139), .A2(n889), .ZN(n890) );
  NAND2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n892) );
  NOR2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n945) );
  XNOR2_X1 U996 ( .A(n894), .B(n945), .ZN(n895) );
  XOR2_X1 U997 ( .A(n895), .B(KEYINPUT46), .Z(n898) );
  XNOR2_X1 U998 ( .A(n896), .B(KEYINPUT48), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n900) );
  XOR2_X1 U1000 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U1001 ( .A(G164), .B(G160), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n906), .B(n905), .Z(n907) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n907), .ZN(G395) );
  XOR2_X1 U1006 ( .A(G286), .B(n1000), .Z(n909) );
  XNOR2_X1 U1007 ( .A(G171), .B(n988), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n912), .ZN(G397) );
  XOR2_X1 U1011 ( .A(G2451), .B(G2430), .Z(n914) );
  XNOR2_X1 U1012 ( .A(G2438), .B(G2443), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n920) );
  XOR2_X1 U1014 ( .A(G2435), .B(G2454), .Z(n916) );
  XNOR2_X1 U1015 ( .A(G1348), .B(G1341), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n916), .B(n915), .ZN(n918) );
  XOR2_X1 U1017 ( .A(G2446), .B(G2427), .Z(n917) );
  XNOR2_X1 U1018 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1019 ( .A(n920), .B(n919), .Z(n921) );
  NAND2_X1 U1020 ( .A1(G14), .A2(n921), .ZN(n927) );
  NAND2_X1 U1021 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(G108), .ZN(G238) );
  INV_X1 U1029 ( .A(n927), .ZN(G401) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(KEYINPUT115), .B(n930), .ZN(n931) );
  NOR2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n944) );
  XOR2_X1 U1033 ( .A(G160), .B(G2084), .Z(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1038 ( .A(KEYINPUT116), .B(n939), .Z(n940) );
  XOR2_X1 U1039 ( .A(KEYINPUT51), .B(n940), .Z(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(G2072), .B(n945), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(G164), .B(G2078), .ZN(n946) );
  NAND2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1045 ( .A(KEYINPUT117), .B(n948), .Z(n949) );
  XNOR2_X1 U1046 ( .A(KEYINPUT50), .B(n949), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n952), .ZN(n953) );
  XOR2_X1 U1049 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n976) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n976), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n954), .A2(G29), .ZN(n1040) );
  XNOR2_X1 U1052 ( .A(G25), .B(n955), .ZN(n956) );
  NAND2_X1 U1053 ( .A1(n956), .A2(G28), .ZN(n963) );
  XOR2_X1 U1054 ( .A(n957), .B(G27), .Z(n960) );
  XOR2_X1 U1055 ( .A(n958), .B(G32), .Z(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1057 ( .A(KEYINPUT120), .B(n961), .Z(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(G2067), .B(G26), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(G33), .B(G2072), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n968), .B(KEYINPUT53), .ZN(n975) );
  XOR2_X1 U1064 ( .A(KEYINPUT121), .B(G34), .Z(n970) );
  XNOR2_X1 U1065 ( .A(G2084), .B(KEYINPUT54), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(n970), .B(n969), .ZN(n973) );
  XOR2_X1 U1067 ( .A(KEYINPUT119), .B(G2090), .Z(n971) );
  XNOR2_X1 U1068 ( .A(G35), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(n977), .B(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(KEYINPUT122), .B(n978), .ZN(n980) );
  INV_X1 U1073 ( .A(G29), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n981), .A2(G11), .ZN(n1038) );
  XNOR2_X1 U1076 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G168), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(KEYINPUT57), .B(n984), .ZN(n1006) );
  XNOR2_X1 U1080 ( .A(n985), .B(G1956), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(G1348), .B(n988), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(G1971), .A2(G303), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(G1961), .B(G301), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(KEYINPUT123), .B(n999), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(n1000), .B(G1341), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1001), .B(KEYINPUT124), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(KEYINPUT125), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1036) );
  INV_X1 U1097 ( .A(G16), .ZN(n1034) );
  XNOR2_X1 U1098 ( .A(G5), .B(n1009), .ZN(n1023) );
  XNOR2_X1 U1099 ( .A(G1348), .B(KEYINPUT59), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(G4), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G1341), .B(G19), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(G6), .B(G1981), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(KEYINPUT126), .B(n1015), .Z(n1016) );
  XNOR2_X1 U1106 ( .A(G20), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1108 ( .A(KEYINPUT60), .B(n1019), .Z(n1021) );
  XNOR2_X1 U1109 ( .A(G1966), .B(G21), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1031) );
  XNOR2_X1 U1112 ( .A(G1971), .B(G22), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(G23), .B(G1976), .ZN(n1024) );
  NOR2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(G1986), .B(KEYINPUT127), .ZN(n1026) );
  XNOR2_X1 U1116 ( .A(n1026), .B(G24), .ZN(n1027) );
  NAND2_X1 U1117 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1118 ( .A(KEYINPUT58), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1119 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1120 ( .A(KEYINPUT61), .B(n1032), .ZN(n1033) );
  NAND2_X1 U1121 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1124 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1041), .Z(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

