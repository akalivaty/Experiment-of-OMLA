//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n203), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n208), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  NOR2_X1   g0019(.A1(new_n208), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n203), .A2(new_n205), .ZN(new_n226));
  INV_X1    g0026(.A(G50), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n222), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G58), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT66), .B(G50), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G97), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n223), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n224), .B1(new_n226), .B2(new_n227), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G150), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n224), .A2(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n249), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n249), .B1(new_n257), .B2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n256), .B(new_n259), .C1(G50), .C2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT9), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(KEYINPUT69), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(KEYINPUT69), .ZN(new_n264));
  XOR2_X1   g0064(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G1), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT67), .B(G45), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G226), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G1), .A3(G13), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n269), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n276), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n277), .A2(G33), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G222), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(G223), .A3(G1698), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n287), .B(new_n288), .C1(new_n210), .C2(new_n285), .ZN(new_n289));
  INV_X1    g0089(.A(new_n272), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n275), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G190), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n265), .B(new_n292), .C1(new_n293), .C2(new_n291), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n261), .C1(G169), .C2(new_n291), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n251), .A2(G50), .ZN(new_n301));
  OAI221_X1 g0101(.A(new_n301), .B1(new_n224), .B2(G68), .C1(new_n210), .C2(new_n254), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n302), .A2(new_n249), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT11), .ZN(new_n304));
  INV_X1    g0104(.A(new_n260), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n202), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(KEYINPUT12), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(KEYINPUT12), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n307), .A2(new_n308), .B1(G68), .B2(new_n258), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n303), .A2(KEYINPUT11), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n300), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n311), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n313), .A2(KEYINPUT72), .A3(new_n304), .A4(new_n309), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT13), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT68), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT68), .B1(new_n282), .B2(new_n283), .ZN(new_n319));
  OAI211_X1 g0119(.A(G232), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(G226), .B(new_n286), .C1(new_n318), .C2(new_n319), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n321), .C1(new_n279), .C2(new_n212), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n290), .ZN(new_n323));
  INV_X1    g0123(.A(G238), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n269), .B1(new_n324), .B2(new_n274), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n317), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  AOI211_X1 g0127(.A(KEYINPUT13), .B(new_n325), .C1(new_n322), .C2(new_n290), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n316), .B1(new_n329), .B2(G200), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n325), .B1(new_n322), .B2(new_n290), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT70), .B1(new_n333), .B2(new_n317), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n333), .A2(KEYINPUT70), .A3(new_n317), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT71), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n332), .B(KEYINPUT71), .C1(new_n334), .C2(new_n335), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n330), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(KEYINPUT73), .B2(KEYINPUT14), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n327), .B2(new_n328), .ZN(new_n344));
  NOR2_X1   g0144(.A1(KEYINPUT73), .A2(KEYINPUT14), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n345), .B(new_n343), .C1(new_n327), .C2(new_n328), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n323), .A2(new_n326), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n296), .B1(new_n349), .B2(KEYINPUT13), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n335), .B2(new_n334), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n347), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT74), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT74), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n347), .A2(new_n351), .A3(new_n354), .A4(new_n348), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n315), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n285), .A2(G232), .A3(new_n286), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n285), .A2(G238), .A3(G1698), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n318), .A2(new_n319), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G107), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n290), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n269), .B1(new_n211), .B2(new_n274), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n342), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n363), .B1(new_n361), .B2(new_n290), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n296), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n258), .A2(G77), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(G77), .B2(new_n260), .ZN(new_n370));
  INV_X1    g0170(.A(new_n253), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT15), .B(G87), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n254), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n370), .B1(new_n249), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n366), .A2(new_n368), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n367), .A2(G190), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(new_n375), .C1(new_n293), .C2(new_n367), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NOR4_X1   g0180(.A1(new_n299), .A2(new_n341), .A3(new_n356), .A4(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n272), .A2(G232), .A3(new_n273), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT78), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT78), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n272), .A2(new_n273), .A3(new_n384), .A4(G232), .ZN(new_n385));
  AND3_X1   g0185(.A1(new_n383), .A2(new_n385), .A3(new_n269), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT75), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(new_n279), .A3(KEYINPUT3), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT75), .B1(new_n277), .B2(G33), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(new_n278), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n270), .A2(G1698), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(G223), .B2(G1698), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n387), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n290), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT79), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n386), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n388), .B1(new_n279), .B2(KEYINPUT3), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n282), .ZN(new_n399));
  NOR2_X1   g0199(.A1(G223), .A2(G1698), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n270), .B2(G1698), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n401), .A3(new_n389), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n272), .B1(new_n402), .B2(new_n387), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n383), .A2(new_n385), .A3(new_n269), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT79), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n397), .A2(new_n405), .A3(new_n342), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n386), .A2(new_n395), .A3(new_n296), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n371), .A2(new_n305), .ZN(new_n410));
  INV_X1    g0210(.A(new_n258), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n411), .B2(new_n371), .ZN(new_n412));
  INV_X1    g0212(.A(new_n249), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n201), .A2(new_n202), .ZN(new_n414));
  OAI21_X1  g0214(.A(G20), .B1(new_n226), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n251), .A2(G159), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n391), .A2(new_n224), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n202), .B1(new_n418), .B2(KEYINPUT7), .ZN(new_n419));
  AOI21_X1  g0219(.A(G20), .B1(new_n399), .B2(new_n389), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT7), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n417), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n413), .B1(new_n423), .B2(KEYINPUT16), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT16), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n281), .A2(new_n224), .A3(new_n284), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n421), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT3), .B(G33), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n421), .A2(G20), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n428), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(KEYINPUT76), .B(new_n430), .C1(new_n278), .C2(new_n280), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n202), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n425), .B1(new_n435), .B2(new_n417), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n412), .B1(new_n424), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT77), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI211_X1 g0239(.A(KEYINPUT77), .B(new_n412), .C1(new_n424), .C2(new_n436), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n409), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n397), .A2(new_n405), .A3(new_n293), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n386), .A2(new_n395), .A3(new_n331), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n437), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT17), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT17), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n437), .A2(new_n447), .A3(new_n444), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n441), .A2(KEYINPUT18), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n412), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT7), .B1(new_n359), .B2(new_n224), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n432), .A2(new_n433), .ZN(new_n452));
  OAI21_X1  g0252(.A(G68), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n415), .A2(new_n416), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT16), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(G68), .B1(new_n420), .B2(new_n421), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n418), .A2(KEYINPUT7), .ZN(new_n457));
  OAI211_X1 g0257(.A(KEYINPUT16), .B(new_n454), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n249), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n450), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT77), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n437), .A2(new_n438), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT18), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n409), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n449), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n466), .B(KEYINPUT80), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n381), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n399), .A2(G244), .A3(new_n389), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(new_n286), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n286), .A2(G238), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n391), .A2(new_n471), .B1(new_n279), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n290), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n257), .A2(G45), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n272), .A2(G250), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT82), .ZN(new_n477));
  INV_X1    g0277(.A(G45), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G1), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G274), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n477), .B1(new_n476), .B2(new_n480), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(G169), .B1(new_n474), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n474), .A2(new_n483), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n296), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n224), .A2(G68), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n254), .A2(new_n212), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n391), .A2(new_n487), .B1(KEYINPUT19), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n490), .A2(KEYINPUT83), .A3(new_n224), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT83), .B1(new_n490), .B2(new_n224), .ZN(new_n492));
  NOR3_X1   g0292(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n249), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n373), .A2(new_n305), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n257), .A2(G33), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n260), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n413), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n495), .B(new_n496), .C1(new_n373), .C2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT84), .ZN(new_n501));
  INV_X1    g0301(.A(G87), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n498), .A2(KEYINPUT84), .A3(new_n413), .A4(G87), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(new_n495), .A3(new_n496), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n474), .A2(new_n483), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(G200), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n485), .A2(G190), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n486), .A2(new_n500), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n469), .B2(G1698), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n211), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n285), .A2(new_n286), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G283), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n512), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n290), .ZN(new_n518));
  XNOR2_X1  g0318(.A(KEYINPUT5), .B(G41), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n290), .B1(new_n519), .B2(new_n479), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G257), .ZN(new_n521));
  XOR2_X1   g0321(.A(KEYINPUT5), .B(G41), .Z(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT81), .B1(new_n522), .B2(new_n480), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT81), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n519), .A2(new_n524), .A3(G274), .A4(new_n479), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n518), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n342), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n527), .B1(new_n517), .B2(new_n290), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n296), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT6), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n245), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(KEYINPUT6), .A3(G97), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G20), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n251), .A2(G77), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n426), .A2(new_n421), .B1(new_n432), .B2(new_n433), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n538), .B(new_n539), .C1(new_n540), .C2(new_n535), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n249), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n305), .A2(new_n212), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n499), .B2(new_n212), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n530), .A2(new_n532), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n531), .A2(G190), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n541), .B2(new_n249), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n549), .C1(new_n293), .C2(new_n531), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n510), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n305), .A2(KEYINPUT25), .A3(new_n535), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT25), .B1(new_n305), .B2(new_n535), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n552), .A2(new_n553), .B1(new_n499), .B2(new_n535), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT22), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n224), .A2(G87), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n359), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(KEYINPUT22), .A2(G87), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n391), .A2(new_n558), .B1(new_n279), .B2(new_n472), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n224), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n224), .A2(G107), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n561), .B(KEYINPUT23), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n557), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n413), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n557), .A2(new_n560), .A3(KEYINPUT24), .A4(new_n562), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n554), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n213), .A2(G1698), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G250), .B2(G1698), .ZN(new_n569));
  INV_X1    g0369(.A(G294), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n391), .A2(new_n569), .B1(new_n279), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n290), .B1(new_n520), .B2(G264), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n526), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT87), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n574), .A3(G169), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n573), .B2(G169), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n573), .A2(new_n296), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n567), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n573), .A2(new_n293), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G190), .B2(new_n573), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n565), .A2(new_n566), .ZN(new_n582));
  INV_X1    g0382(.A(new_n554), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n520), .A2(G270), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n526), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n281), .A2(G303), .A3(new_n284), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n213), .A2(new_n286), .ZN(new_n589));
  OR2_X1    g0389(.A1(new_n286), .A2(G264), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n399), .A2(new_n389), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n272), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT85), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n591), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n290), .ZN(new_n595));
  AOI22_X1  g0395(.A1(G270), .A2(new_n520), .B1(new_n523), .B2(new_n525), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT85), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n593), .A2(new_n598), .A3(G190), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n293), .B1(new_n593), .B2(new_n598), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n248), .A2(new_n223), .B1(G20), .B2(new_n472), .ZN(new_n601));
  AOI21_X1  g0401(.A(G20), .B1(G33), .B2(G283), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n279), .A2(G97), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT86), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n604), .B1(new_n602), .B2(new_n603), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n607), .B(new_n608), .ZN(new_n609));
  MUX2_X1   g0409(.A(new_n260), .B(new_n499), .S(G116), .Z(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n599), .A2(new_n600), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n593), .A2(new_n598), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n342), .B1(new_n609), .B2(new_n610), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(KEYINPUT21), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n587), .A2(new_n592), .A3(new_n296), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT21), .B1(new_n613), .B2(new_n614), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n612), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n551), .A2(new_n585), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n468), .A2(new_n621), .ZN(G372));
  INV_X1    g0422(.A(new_n468), .ZN(new_n623));
  INV_X1    g0423(.A(new_n547), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(KEYINPUT26), .A3(new_n510), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n486), .A2(new_n500), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n508), .A2(new_n509), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n626), .B1(new_n629), .B2(new_n547), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n625), .A2(new_n630), .B1(new_n500), .B2(new_n486), .ZN(new_n631));
  INV_X1    g0431(.A(new_n584), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n618), .A2(new_n619), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n551), .B(new_n632), .C1(new_n579), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n623), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n446), .A2(new_n448), .ZN(new_n637));
  INV_X1    g0437(.A(new_n356), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n367), .A2(new_n296), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n376), .B1(new_n367), .B2(G169), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT88), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT88), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n366), .A2(new_n642), .A3(new_n368), .A4(new_n376), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n340), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n637), .B1(new_n638), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n460), .A2(new_n409), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT18), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n295), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n649), .A2(new_n298), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n636), .A2(new_n650), .ZN(G369));
  INV_X1    g0451(.A(G13), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(G20), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n257), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n611), .A2(new_n659), .ZN(new_n660));
  MUX2_X1   g0460(.A(new_n633), .B(new_n620), .S(new_n660), .Z(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT89), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT90), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n661), .A2(KEYINPUT89), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n661), .A2(KEYINPUT89), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(KEYINPUT90), .A3(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n659), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n585), .B1(new_n567), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n579), .A2(new_n659), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n668), .A2(G330), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n585), .A2(new_n633), .A3(new_n669), .ZN(new_n675));
  INV_X1    g0475(.A(new_n579), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n659), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(KEYINPUT92), .ZN(new_n680));
  INV_X1    g0480(.A(new_n220), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT91), .B1(new_n681), .B2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n681), .A2(KEYINPUT91), .A3(G41), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n493), .A2(new_n472), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n685), .A2(new_n257), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n228), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n680), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n680), .B2(new_n687), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT28), .Z(new_n691));
  AOI21_X1  g0491(.A(new_n659), .B1(new_n631), .B2(new_n634), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT93), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(KEYINPUT93), .A2(KEYINPUT29), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n692), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n551), .A2(new_n585), .A3(new_n620), .A4(new_n669), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n474), .A2(new_n483), .A3(new_n572), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n531), .A2(new_n702), .A3(new_n616), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(G179), .B1(new_n572), .B2(new_n526), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n529), .A2(new_n507), .A3(new_n613), .A4(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n531), .A2(new_n702), .A3(KEYINPUT30), .A4(new_n616), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n701), .B1(new_n709), .B2(new_n659), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n700), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(new_n701), .A3(new_n659), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n711), .A2(G330), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n699), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n691), .B1(new_n716), .B2(G1), .ZN(G364));
  NAND3_X1  g0517(.A1(new_n664), .A2(G330), .A3(new_n667), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n257), .B1(new_n653), .B2(G45), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n685), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G330), .B2(new_n668), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT94), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(G13), .A2(G33), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n662), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n223), .B1(G20), .B2(new_n342), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n224), .A2(G190), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n734), .A2(G179), .A3(G200), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n735), .A2(KEYINPUT96), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(KEYINPUT96), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G329), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n331), .A2(G179), .A3(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n224), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G294), .ZN(new_n744));
  NOR4_X1   g0544(.A1(new_n224), .A2(new_n296), .A3(new_n331), .A4(G200), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G322), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n224), .A2(new_n331), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n293), .A2(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G303), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n746), .A2(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n285), .ZN(new_n753));
  XOR2_X1   g0553(.A(KEYINPUT33), .B(G317), .Z(new_n754));
  NOR2_X1   g0554(.A1(new_n296), .A2(new_n293), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n733), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n748), .A2(new_n755), .ZN(new_n758));
  INV_X1    g0558(.A(G326), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n733), .A2(new_n749), .ZN(new_n760));
  INV_X1    g0560(.A(G283), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n734), .A2(new_n296), .A3(G200), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n757), .B(new_n762), .C1(G311), .C2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n740), .A2(new_n744), .A3(new_n753), .A4(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n763), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n766), .A2(new_n210), .B1(new_n535), .B2(new_n760), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n746), .A2(new_n201), .B1(new_n750), .B2(new_n502), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n735), .A2(G159), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT32), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n770), .A2(KEYINPUT32), .B1(G97), .B2(new_n743), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n758), .A2(new_n227), .B1(new_n756), .B2(new_n202), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n359), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n769), .A2(new_n771), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n732), .B1(new_n765), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n729), .A2(new_n731), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n285), .A2(new_n220), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT95), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n780), .A2(G355), .B1(new_n472), .B2(new_n681), .ZN(new_n781));
  INV_X1    g0581(.A(new_n391), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n681), .ZN(new_n783));
  INV_X1    g0583(.A(new_n268), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n228), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n783), .B(new_n785), .C1(new_n243), .C2(new_n478), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n778), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n776), .A2(new_n722), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n730), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n724), .A2(new_n725), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n726), .A2(new_n789), .A3(new_n790), .ZN(G396));
  NAND2_X1  g0591(.A1(new_n376), .A2(new_n659), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n641), .B2(new_n643), .ZN(new_n793));
  AND3_X1   g0593(.A1(new_n377), .A2(new_n379), .A3(new_n792), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n692), .B(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n721), .B1(new_n796), .B2(new_n713), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n797), .A2(KEYINPUT98), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(KEYINPUT98), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(new_n713), .C2(new_n796), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n731), .A2(new_n727), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n722), .B1(new_n210), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n760), .A2(new_n202), .ZN(new_n803));
  INV_X1    g0603(.A(new_n750), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(G50), .B2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n805), .B(new_n782), .C1(new_n201), .C2(new_n742), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n739), .B2(G132), .ZN(new_n807));
  INV_X1    g0607(.A(new_n756), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G150), .A2(new_n808), .B1(new_n745), .B2(G143), .ZN(new_n809));
  INV_X1    g0609(.A(G137), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(new_n810), .B2(new_n758), .C1(new_n811), .C2(new_n766), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT34), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n359), .B1(new_n502), .B2(new_n760), .C1(new_n751), .C2(new_n758), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n763), .A2(G116), .B1(new_n808), .B2(G283), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n535), .B2(new_n750), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n814), .B(new_n816), .C1(new_n739), .C2(G311), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n743), .A2(G97), .B1(G294), .B2(new_n745), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n807), .A2(new_n813), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n795), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n802), .B1(new_n732), .B2(new_n820), .C1(new_n821), .C2(new_n728), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n800), .A2(new_n822), .ZN(G384));
  OAI211_X1 g0623(.A(new_n228), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(G50), .B2(new_n202), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n825), .A2(G1), .A3(new_n652), .ZN(new_n826));
  OAI211_X1 g0626(.A(G116), .B(new_n225), .C1(new_n537), .C2(KEYINPUT35), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT99), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n827), .A2(new_n828), .B1(KEYINPUT35), .B2(new_n537), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  XNOR2_X1  g0630(.A(KEYINPUT100), .B(KEYINPUT36), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n826), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n830), .B2(new_n831), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n423), .A2(KEYINPUT16), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n450), .B1(new_n459), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n657), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n466), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n409), .A2(new_n835), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n840), .A2(new_n445), .A3(new_n837), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n841), .A2(KEYINPUT37), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT37), .B1(new_n437), .B2(new_n444), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n441), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT101), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n463), .A2(new_n845), .A3(new_n836), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n836), .B1(new_n439), .B2(new_n440), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT101), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n844), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n839), .B(KEYINPUT38), .C1(new_n842), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n846), .ZN(new_n852));
  INV_X1    g0652(.A(new_n844), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n842), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n837), .B1(new_n449), .B2(new_n465), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n442), .A2(new_n443), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT102), .B1(new_n460), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT102), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n437), .A2(new_n861), .A3(new_n444), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n647), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT103), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT103), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n860), .A2(new_n865), .A3(new_n862), .A4(new_n647), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n845), .B1(new_n463), .B2(new_n836), .ZN(new_n867));
  AOI211_X1 g0667(.A(KEYINPUT101), .B(new_n657), .C1(new_n461), .C2(new_n462), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n864), .B(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n849), .B1(new_n869), .B2(KEYINPUT37), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n648), .A2(new_n637), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(new_n852), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n851), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n874), .A3(new_n850), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n858), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n356), .A2(new_n669), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n648), .A2(new_n657), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n315), .A2(new_n669), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n356), .A2(new_n341), .A3(new_n880), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n315), .B(new_n669), .C1(new_n353), .C2(new_n355), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n377), .A2(new_n659), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n692), .B2(new_n821), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n857), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n879), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n878), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n381), .A2(new_n467), .A3(new_n698), .A4(new_n696), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n650), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n889), .B(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n894));
  INV_X1    g0694(.A(new_n849), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n872), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n850), .B1(new_n896), .B2(KEYINPUT38), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n711), .A2(new_n712), .A3(new_n821), .ZN(new_n898));
  INV_X1    g0698(.A(new_n880), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n638), .A2(new_n340), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n882), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n893), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n857), .A2(new_n902), .A3(new_n893), .ZN(new_n904));
  OAI21_X1  g0704(.A(G330), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n381), .A2(new_n467), .A3(new_n713), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n857), .A2(new_n902), .A3(new_n893), .ZN(new_n908));
  INV_X1    g0708(.A(new_n712), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n909), .B(new_n795), .C1(new_n700), .C2(new_n710), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n881), .B2(new_n882), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n873), .B2(new_n850), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n908), .B1(new_n912), .B2(new_n893), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n913), .A2(new_n623), .A3(new_n711), .A4(new_n712), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n892), .A2(new_n915), .B1(new_n257), .B2(new_n653), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n892), .A2(new_n915), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n833), .B1(new_n916), .B2(new_n917), .ZN(G367));
  OAI211_X1 g0718(.A(new_n547), .B(new_n550), .C1(new_n549), .C2(new_n669), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n547), .B2(new_n669), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT104), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT105), .B1(new_n921), .B2(new_n675), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT104), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n920), .B(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT105), .ZN(new_n925));
  INV_X1    g0725(.A(new_n675), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n922), .A2(KEYINPUT42), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n547), .B1(new_n921), .B2(new_n676), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n669), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n506), .A2(new_n659), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n510), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n627), .B2(new_n932), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT42), .B1(new_n922), .B2(new_n927), .ZN(new_n936));
  OR3_X1    g0736(.A1(new_n931), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT106), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n935), .B(new_n940), .C1(new_n931), .C2(new_n936), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n937), .B2(KEYINPUT106), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n939), .A2(new_n942), .B1(new_n674), .B2(new_n921), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n937), .A2(KEYINPUT106), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n674), .A2(new_n921), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n944), .A2(new_n945), .A3(new_n938), .A4(new_n941), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n685), .B(KEYINPUT41), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n633), .A2(new_n669), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n926), .B1(new_n672), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n668), .A2(G330), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n718), .A2(new_n949), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n715), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT45), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n921), .B2(new_n677), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n924), .A2(KEYINPUT45), .A3(new_n678), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT44), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n924), .B2(new_n678), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n921), .A2(KEYINPUT44), .A3(new_n677), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n674), .B1(new_n963), .B2(KEYINPUT107), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n718), .A2(new_n672), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT107), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(new_n966), .A3(new_n962), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n953), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n947), .B1(new_n968), .B2(new_n716), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n943), .B(new_n946), .C1(new_n969), .C2(new_n720), .ZN(new_n970));
  INV_X1    g0770(.A(new_n783), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n777), .B1(new_n220), .B2(new_n373), .C1(new_n971), .C2(new_n238), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n721), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n750), .A2(new_n472), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G107), .B2(new_n743), .ZN(new_n976));
  INV_X1    g0776(.A(new_n760), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G294), .A2(new_n808), .B1(new_n977), .B2(G97), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G283), .A2(new_n763), .B1(new_n735), .B2(G317), .ZN(new_n979));
  INV_X1    g0779(.A(G311), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n746), .A2(new_n751), .B1(new_n758), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n782), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n976), .A2(new_n978), .A3(new_n979), .A4(new_n982), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n766), .A2(new_n227), .B1(new_n811), .B2(new_n756), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT110), .ZN(new_n985));
  INV_X1    g0785(.A(new_n735), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n986), .A2(new_n810), .B1(new_n201), .B2(new_n750), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n984), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n977), .A2(G77), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n285), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT109), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n988), .B(new_n991), .C1(new_n985), .C2(new_n987), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n748), .A2(new_n755), .A3(G143), .ZN(new_n993));
  INV_X1    g0793(.A(G150), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n993), .B1(new_n202), .B2(new_n742), .C1(new_n746), .C2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT108), .Z(new_n996));
  OAI21_X1  g0796(.A(new_n983), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT47), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n732), .B1(new_n997), .B2(new_n998), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n973), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n729), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1001), .B1(new_n934), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n970), .A2(new_n1003), .ZN(G387));
  INV_X1    g0804(.A(new_n685), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n953), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n951), .A2(new_n952), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1006), .B1(new_n716), .B2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n780), .A2(new_n686), .B1(new_n535), .B2(new_n681), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n478), .B1(new_n202), .B2(new_n210), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n371), .A2(new_n227), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n686), .B(new_n1010), .C1(new_n1011), .C2(KEYINPUT50), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n971), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n235), .B2(new_n784), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n1009), .A2(KEYINPUT111), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT111), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1016), .A2(new_n778), .A3(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n763), .A2(G68), .B1(new_n808), .B2(new_n371), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT112), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n986), .A2(new_n994), .B1(new_n212), .B2(new_n760), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n742), .A2(new_n373), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1021), .A2(new_n391), .A3(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n758), .A2(new_n811), .B1(new_n750), .B2(new_n210), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G50), .B2(new_n745), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1020), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n735), .A2(G326), .B1(new_n977), .B2(G116), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G311), .A2(new_n808), .B1(new_n745), .B2(G317), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n747), .B2(new_n758), .C1(new_n751), .C2(new_n766), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT48), .Z(new_n1030));
  OAI22_X1  g0830(.A1(new_n742), .A2(new_n761), .B1(new_n750), .B2(new_n570), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n391), .B(new_n1027), .C1(new_n1032), .C2(KEYINPUT49), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1032), .A2(KEYINPUT49), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1026), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n731), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n721), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1018), .B(new_n1037), .C1(new_n672), .C2(new_n729), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n1007), .B2(new_n720), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1008), .A2(new_n1039), .ZN(G393));
  XNOR2_X1  g0840(.A(new_n965), .B(new_n963), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n720), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n777), .B1(new_n212), .B2(new_n220), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n246), .B2(new_n783), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n722), .A2(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n782), .B1(new_n202), .B2(new_n750), .C1(new_n502), .C2(new_n760), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n735), .A2(G143), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n227), .B2(new_n756), .C1(new_n766), .C2(new_n253), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1046), .B(new_n1048), .C1(G77), .C2(new_n743), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n746), .A2(new_n811), .B1(new_n758), .B2(new_n994), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT51), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n756), .A2(new_n751), .B1(new_n760), .B2(new_n535), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n285), .B(new_n1052), .C1(G116), .C2(new_n743), .ZN(new_n1053));
  INV_X1    g0853(.A(G317), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n746), .A2(new_n980), .B1(new_n758), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT52), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n763), .A2(G294), .B1(new_n804), .B2(G283), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n747), .B2(new_n986), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1049), .A2(new_n1051), .B1(new_n1053), .B2(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1045), .B1(new_n732), .B2(new_n1062), .C1(new_n924), .C2(new_n1002), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n685), .B1(new_n1041), .B2(new_n953), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n968), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1042), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(G390));
  OAI21_X1  g0866(.A(new_n877), .B1(new_n883), .B2(new_n885), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n858), .A2(new_n875), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n713), .A2(new_n821), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(new_n883), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n886), .A2(new_n897), .A3(new_n877), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1070), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1072), .A2(new_n1073), .A3(new_n719), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT114), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n650), .A2(new_n890), .A3(new_n906), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n821), .A2(KEYINPUT113), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n883), .A2(new_n885), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n886), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n713), .A3(new_n821), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n886), .A2(new_n1069), .A3(new_n1080), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1076), .A2(new_n1078), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1078), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n1073), .B2(new_n1072), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1085), .A2(new_n1087), .A3(new_n685), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n876), .A2(new_n727), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n722), .B1(new_n253), .B2(new_n801), .ZN(new_n1090));
  INV_X1    g0890(.A(G132), .ZN(new_n1091));
  INV_X1    g0891(.A(G128), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n746), .A2(new_n1091), .B1(new_n758), .B2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n739), .A2(G125), .B1(new_n1093), .B2(KEYINPUT115), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n750), .A2(new_n994), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT53), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(KEYINPUT115), .C2(new_n1093), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n359), .B1(G159), .B2(new_n743), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT54), .B(G143), .Z(new_n1099));
  AOI22_X1  g0899(.A1(new_n763), .A2(new_n1099), .B1(new_n808), .B2(G137), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(new_n227), .C2(new_n760), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n803), .B1(G87), .B2(new_n804), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1102), .B(new_n359), .C1(new_n210), .C2(new_n742), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n758), .A2(new_n761), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G97), .B2(new_n763), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G107), .A2(new_n808), .B1(new_n745), .B2(G116), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(new_n738), .C2(new_n570), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1097), .A2(new_n1101), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n731), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1089), .B(new_n1090), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1075), .A2(new_n1088), .A3(new_n1112), .ZN(G378));
  NAND2_X1  g0913(.A1(new_n261), .A2(new_n836), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n299), .B(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n905), .A2(KEYINPUT122), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT122), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n913), .A2(new_n1119), .A3(G330), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1117), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1119), .B1(new_n913), .B2(G330), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1117), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n1121), .A2(new_n889), .A3(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n878), .A2(new_n888), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n913), .A2(new_n1119), .A3(G330), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1123), .B1(new_n1127), .B2(new_n1122), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1118), .A2(new_n1117), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n720), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1123), .A2(new_n727), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n801), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n721), .B1(G50), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n782), .A2(G41), .ZN(new_n1135));
  INV_X1    g0935(.A(G41), .ZN(new_n1136));
  AOI211_X1 g0936(.A(G50), .B(new_n1135), .C1(new_n279), .C2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT117), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n758), .A2(new_n472), .B1(new_n750), .B2(new_n210), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n746), .A2(new_n535), .B1(new_n760), .B2(new_n201), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(G68), .C2(new_n743), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1141), .B(new_n1135), .C1(new_n761), .C2(new_n738), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n766), .A2(new_n373), .B1(new_n212), .B2(new_n756), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT118), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1138), .B1(new_n1145), .B2(KEYINPUT58), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n804), .A2(new_n1099), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT119), .Z(new_n1148));
  NOR2_X1   g0948(.A1(new_n742), .A2(new_n994), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n766), .A2(new_n810), .B1(new_n1091), .B2(new_n756), .ZN(new_n1150));
  INV_X1    g0950(.A(G125), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n746), .A2(new_n1092), .B1(new_n758), .B2(new_n1151), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n279), .B(new_n1136), .C1(new_n760), .C2(new_n811), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G124), .B2(new_n735), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1146), .B1(KEYINPUT58), .B2(new_n1145), .C1(new_n1155), .C2(new_n1159), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1160), .A2(KEYINPUT121), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n732), .B1(new_n1160), .B2(KEYINPUT121), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1134), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1132), .A2(new_n1163), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1131), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1077), .B1(new_n1076), .B2(new_n1084), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT57), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT123), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n889), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT123), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1169), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1128), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1166), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n685), .B1(new_n1176), .B2(KEYINPUT57), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1165), .B1(new_n1174), .B2(new_n1177), .ZN(G375));
  INV_X1    g0978(.A(new_n947), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1082), .A2(new_n1077), .A3(new_n1083), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1086), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n989), .B1(new_n472), .B2(new_n756), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1182), .A2(new_n285), .A3(new_n1022), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n766), .A2(new_n535), .B1(new_n212), .B2(new_n750), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n746), .A2(new_n761), .B1(new_n758), .B2(new_n570), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n739), .C2(G303), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n746), .A2(new_n810), .B1(new_n758), .B2(new_n1091), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n808), .A2(new_n1099), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n766), .B2(new_n994), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(new_n739), .C2(G128), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n750), .A2(new_n811), .B1(new_n760), .B2(new_n201), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n391), .B(new_n1191), .C1(G50), .C2(new_n743), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1183), .A2(new_n1186), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n721), .B1(G68), .B2(new_n1133), .C1(new_n1193), .C2(new_n732), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n883), .B2(new_n727), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n1084), .B2(new_n720), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1181), .A2(new_n1196), .ZN(G381));
  INV_X1    g0997(.A(KEYINPUT124), .ZN(new_n1198));
  AOI21_X1  g0998(.A(G378), .B1(G375), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1198), .B2(G375), .ZN(new_n1200));
  INV_X1    g1000(.A(G390), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(G393), .A2(G396), .ZN(new_n1202));
  INV_X1    g1002(.A(G384), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(G381), .ZN(new_n1205));
  OR3_X1    g1005(.A1(new_n1200), .A2(G387), .A3(new_n1205), .ZN(G407));
  OAI211_X1 g1006(.A(G407), .B(G213), .C1(G343), .C2(new_n1200), .ZN(G409));
  OAI211_X1 g1007(.A(G378), .B(new_n1165), .C1(new_n1174), .C2(new_n1177), .ZN(new_n1208));
  INV_X1    g1008(.A(G378), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n719), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1166), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1179), .B(new_n1211), .C1(new_n1125), .C2(new_n1130), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1164), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1209), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1208), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT60), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1180), .A2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1082), .A2(new_n1077), .A3(KEYINPUT60), .A4(new_n1083), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1217), .A2(new_n1086), .A3(new_n685), .A4(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(G384), .A3(new_n1196), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(G384), .B1(new_n1219), .B2(new_n1196), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(G213), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(G343), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1215), .A2(new_n1223), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT62), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT61), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1225), .B1(new_n1208), .B2(new_n1214), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT62), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n1223), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT125), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1221), .A2(new_n1233), .A3(new_n1222), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1225), .A2(G2897), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1223), .A2(KEYINPUT125), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1233), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1236), .B1(new_n1239), .B2(new_n1235), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT123), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1130), .A2(new_n1170), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n720), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1164), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G378), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1131), .A2(new_n1164), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1211), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1005), .B1(new_n1248), .B2(new_n1167), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1168), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1247), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1246), .B1(G378), .B2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1240), .B1(new_n1252), .B2(new_n1225), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1228), .A2(new_n1229), .A3(new_n1232), .A4(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G390), .B1(new_n970), .B2(new_n1003), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1258), .A2(new_n1202), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n970), .A2(new_n1003), .A3(G390), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1257), .A2(new_n1259), .B1(new_n1261), .B2(new_n1255), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1259), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1255), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1256), .A4(new_n1260), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1254), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1222), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT125), .B1(new_n1269), .B2(new_n1220), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1235), .B1(new_n1270), .B2(new_n1234), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1235), .B2(new_n1234), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1268), .B(new_n1229), .C1(new_n1230), .C2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1227), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT127), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1227), .B2(new_n1275), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1230), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1223), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1274), .A2(new_n1276), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1267), .A2(new_n1280), .ZN(G405));
  INV_X1    g1081(.A(new_n1208), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1251), .A2(G378), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1266), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1282), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1268), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1284), .A2(new_n1223), .A3(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1223), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(G402));
endmodule


