//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990;
  INV_X1    g000(.A(G230gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208));
  INV_X1    g007(.A(G85gat), .ZN(new_n209));
  INV_X1    g008(.A(G92gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(KEYINPUT8), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G99gat), .B(G106gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT96), .B(G64gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G57gat), .ZN(new_n216));
  INV_X1    g015(.A(G64gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n216), .B(KEYINPUT97), .C1(G57gat), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G71gat), .A2(G78gat), .ZN(new_n219));
  INV_X1    g018(.A(G71gat), .ZN(new_n220));
  INV_X1    g019(.A(G78gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT9), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n219), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n218), .B(new_n224), .C1(KEYINPUT97), .C2(new_n216), .ZN(new_n225));
  XNOR2_X1  g024(.A(G57gat), .B(G64gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n219), .B(new_n222), .C1(new_n226), .C2(new_n223), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n214), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT10), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n212), .B(new_n213), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n227), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(new_n229), .A3(new_n228), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n204), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n228), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(new_n204), .ZN(new_n237));
  XNOR2_X1  g036(.A(G120gat), .B(G148gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(G176gat), .B(G204gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n238), .B(new_n239), .Z(new_n240));
  OR2_X1    g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n235), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n204), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n243), .A3(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT21), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n232), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G231gat), .A2(G233gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G127gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G8gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(G15gat), .B(G22gat), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n253), .A2(G1gat), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n254), .B2(KEYINPUT94), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT16), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n253), .B1(new_n256), .B2(G1gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n255), .B(new_n258), .Z(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n232), .B2(new_n246), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n251), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n262));
  INV_X1    g061(.A(G155gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G183gat), .B(G211gat), .Z(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n261), .A2(new_n266), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G43gat), .B(G50gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT15), .ZN(new_n271));
  NOR2_X1   g070(.A1(G29gat), .A2(G36gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT14), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G29gat), .ZN(new_n275));
  INV_X1    g074(.A(G36gat), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT93), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OR3_X1    g076(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT93), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(KEYINPUT15), .A3(new_n270), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT17), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(new_n214), .ZN(new_n286));
  NAND2_X1  g085(.A1(G232gat), .A2(G233gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT98), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G190gat), .B(G218gat), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n289), .A2(KEYINPUT41), .B1(KEYINPUT101), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n283), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(new_n231), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n286), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n290), .A2(KEYINPUT101), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n289), .A2(KEYINPUT41), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n297), .B(KEYINPUT99), .Z(new_n298));
  XNOR2_X1  g097(.A(G134gat), .B(G162gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n300), .A2(KEYINPUT102), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n300), .B(KEYINPUT102), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n269), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT64), .ZN(new_n310));
  INV_X1    g109(.A(G169gat), .ZN(new_n311));
  INV_X1    g110(.A(G176gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n314), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n311), .A2(new_n312), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT67), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n316), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT27), .B(G183gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329));
  AOI21_X1  g128(.A(G190gat), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n327), .B(new_n330), .C1(new_n328), .C2(new_n329), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n328), .A2(new_n329), .ZN(new_n332));
  INV_X1    g131(.A(G183gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT27), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT27), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G183gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(KEYINPUT66), .B2(KEYINPUT28), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n325), .A2(new_n326), .A3(new_n331), .A4(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT25), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n317), .A2(KEYINPUT23), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n342), .B1(new_n343), .B2(new_n320), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n313), .A2(KEYINPUT23), .A3(new_n315), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(G183gat), .B2(G190gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT24), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n326), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT65), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT65), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n348), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n346), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n323), .B1(KEYINPUT23), .B2(new_n317), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT23), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  AND2_X1   g159(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(G190gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n350), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT25), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n341), .B1(new_n356), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n309), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n326), .A2(KEYINPUT65), .A3(new_n349), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT65), .B1(new_n326), .B2(new_n349), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n362), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(new_n345), .A3(new_n344), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n343), .A2(new_n320), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n323), .A2(KEYINPUT23), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n347), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n375), .A2(new_n353), .A3(new_n360), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n342), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n371), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n308), .B1(new_n378), .B2(new_n341), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n367), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G211gat), .B(G218gat), .Z(new_n381));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n382));
  XOR2_X1   g181(.A(G197gat), .B(G204gat), .Z(new_n383));
  AOI21_X1  g182(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OR2_X1    g184(.A1(G197gat), .A2(G204gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(G197gat), .A2(G204gat), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT77), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n381), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  AOI211_X1 g189(.A(new_n382), .B(new_n384), .C1(new_n386), .C2(new_n387), .ZN(new_n391));
  INV_X1    g190(.A(new_n381), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n395), .ZN(new_n396));
  XOR2_X1   g195(.A(G8gat), .B(G36gat), .Z(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT81), .ZN(new_n398));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n379), .A2(KEYINPUT80), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n365), .A2(new_n309), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT79), .B(KEYINPUT29), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n404), .B1(new_n378), .B2(new_n341), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n402), .B1(new_n405), .B2(new_n309), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n401), .B1(new_n406), .B2(KEYINPUT80), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT78), .B1(new_n390), .B2(new_n393), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n388), .A2(KEYINPUT77), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n392), .B1(new_n409), .B2(new_n391), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n389), .A2(new_n381), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n396), .B(new_n400), .C1(new_n407), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT89), .B1(new_n380), .B2(new_n395), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT89), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n418), .B(new_n394), .C1(new_n367), .C2(new_n379), .ZN(new_n419));
  INV_X1    g218(.A(new_n401), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n365), .A2(new_n403), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n379), .B1(new_n421), .B2(new_n308), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n414), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n417), .B(new_n419), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT38), .B1(new_n426), .B2(KEYINPUT37), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n424), .A2(new_n425), .B1(new_n395), .B2(new_n380), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT37), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n400), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n416), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G1gat), .B(G29gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT0), .ZN(new_n433));
  XNOR2_X1  g232(.A(G57gat), .B(G85gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  NAND2_X1  g234(.A1(G225gat), .A2(G233gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT83), .B(G162gat), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT2), .B1(new_n439), .B2(new_n263), .ZN(new_n440));
  INV_X1    g239(.A(G141gat), .ZN(new_n441));
  INV_X1    g240(.A(G148gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(G162gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(G155gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n263), .A2(G162gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(G141gat), .A2(G148gat), .ZN(new_n447));
  AND4_X1   g246(.A1(new_n443), .A2(new_n445), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT2), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n443), .A2(new_n449), .A3(new_n447), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n446), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n440), .A2(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT3), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n438), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n451), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n444), .A2(KEYINPUT83), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(G162gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n449), .B1(new_n459), .B2(G155gat), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n443), .A2(new_n445), .A3(new_n446), .A4(new_n447), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n455), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(KEYINPUT84), .A3(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n454), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G120gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G113gat), .ZN(new_n466));
  INV_X1    g265(.A(G113gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G120gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT1), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G134gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G127gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n250), .A2(G134gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT68), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n473), .B2(new_n474), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT69), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(new_n465), .B2(G113gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n467), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n466), .A3(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n482), .A2(new_n470), .A3(new_n473), .A4(new_n474), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n455), .B(new_n453), .C1(new_n460), .C2(new_n461), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI211_X1 g285(.A(KEYINPUT5), .B(new_n437), .C1(new_n464), .C2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT4), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n484), .A2(new_n462), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT70), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT1), .B1(new_n466), .B2(new_n468), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n250), .A2(G134gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n472), .A2(G127gat), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT68), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n473), .A2(new_n474), .A3(new_n470), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT69), .B1(new_n467), .B2(G120gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n467), .A2(G120gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n500), .B2(new_n481), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n490), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n478), .A2(KEYINPUT70), .A3(new_n483), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n452), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n489), .B1(new_n488), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n505), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n452), .A2(new_n438), .A3(new_n453), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT84), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n486), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT4), .A4(new_n452), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n488), .B1(new_n484), .B2(new_n462), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n509), .A2(new_n436), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT5), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n484), .B(new_n462), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(new_n437), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n435), .B1(new_n506), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT85), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT6), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n517), .B2(KEYINPUT6), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n428), .A2(new_n429), .ZN(new_n522));
  INV_X1    g321(.A(new_n400), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n396), .B1(new_n407), .B2(new_n414), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(KEYINPUT37), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT38), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n487), .A2(new_n505), .B1(new_n512), .B2(new_n515), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(new_n435), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT6), .B1(new_n528), .B2(new_n435), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n506), .A2(new_n516), .ZN(new_n531));
  INV_X1    g330(.A(new_n435), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(KEYINPUT88), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n431), .A2(new_n521), .A3(new_n526), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G228gat), .A2(G233gat), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n403), .B1(new_n390), .B2(new_n393), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n452), .B1(new_n537), .B2(new_n453), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n485), .A2(new_n403), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n394), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT29), .B1(new_n410), .B2(new_n412), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n462), .B1(new_n542), .B2(KEYINPUT3), .ZN(new_n543));
  INV_X1    g342(.A(new_n536), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n408), .A2(new_n413), .A3(new_n539), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G22gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n541), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT86), .ZN(new_n549));
  XNOR2_X1  g348(.A(G78gat), .B(G106gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT31), .B(G50gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n541), .A2(new_n546), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G22gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n548), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n549), .A2(new_n555), .A3(new_n548), .A4(new_n552), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT82), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n415), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT30), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n428), .A2(new_n400), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n415), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n529), .A2(new_n533), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n505), .A2(new_n509), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n437), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n514), .A2(new_n437), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(KEYINPUT39), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n435), .B1(new_n569), .B2(KEYINPUT39), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT40), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n569), .A2(KEYINPUT39), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT40), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n575), .A2(new_n576), .A3(new_n435), .A4(new_n571), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n566), .A2(new_n567), .A3(new_n578), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n535), .A2(new_n559), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581));
  XNOR2_X1  g380(.A(G15gat), .B(G43gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT72), .ZN(new_n583));
  XNOR2_X1  g382(.A(G71gat), .B(G99gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G227gat), .A2(G233gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AND4_X1   g386(.A1(new_n502), .A2(new_n378), .A3(new_n503), .A4(new_n341), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n378), .A2(new_n341), .B1(new_n502), .B2(new_n503), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n585), .B1(new_n590), .B2(KEYINPUT32), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(KEYINPUT71), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT71), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n502), .A2(new_n503), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n365), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n378), .A2(new_n502), .A3(new_n503), .A4(new_n341), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n586), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n594), .B1(new_n598), .B2(KEYINPUT33), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n591), .A2(new_n593), .A3(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n590), .B(KEYINPUT32), .C1(new_n592), .C2(new_n585), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(new_n586), .A3(new_n597), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT73), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n604), .B1(new_n602), .B2(new_n603), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n600), .A2(new_n601), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n600), .B2(new_n601), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n581), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT76), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT75), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n602), .A2(new_n603), .ZN(new_n614));
  INV_X1    g413(.A(new_n604), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI211_X1 g417(.A(new_n613), .B(new_n618), .C1(new_n601), .C2(new_n600), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n601), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n607), .B1(new_n620), .B2(KEYINPUT75), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT36), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(KEYINPUT76), .B(new_n581), .C1(new_n608), .C2(new_n609), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n612), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n559), .ZN(new_n625));
  INV_X1    g424(.A(new_n517), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n530), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n531), .A2(KEYINPUT6), .A3(new_n532), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT85), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT6), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n625), .B1(new_n631), .B2(new_n566), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT87), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n580), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n624), .A2(new_n632), .A3(KEYINPUT87), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT90), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n534), .A2(new_n630), .A3(new_n629), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT35), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n608), .A2(new_n609), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .A4(new_n559), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n637), .B1(new_n641), .B2(new_n566), .ZN(new_n642));
  INV_X1    g441(.A(new_n640), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n643), .A2(new_n625), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT35), .B1(new_n521), .B2(new_n534), .ZN(new_n645));
  INV_X1    g444(.A(new_n566), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT90), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n559), .B1(new_n619), .B2(new_n621), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT91), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n631), .A2(new_n566), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n559), .B(KEYINPUT91), .C1(new_n619), .C2(new_n621), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT35), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n635), .A2(new_n636), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  MUX2_X1   g455(.A(new_n292), .B(new_n285), .S(new_n259), .Z(new_n657));
  NAND2_X1  g456(.A1(G229gat), .A2(G233gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(KEYINPUT18), .A3(new_n658), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n259), .B(new_n292), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n658), .B(KEYINPUT13), .Z(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G113gat), .B(G141gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(G169gat), .B(G197gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT12), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n661), .A2(new_n662), .A3(new_n665), .A4(new_n672), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT95), .B1(new_n656), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n633), .A2(new_n634), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n535), .A2(new_n559), .A3(new_n579), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n636), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n648), .A2(new_n655), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT95), .ZN(new_n683));
  INV_X1    g482(.A(new_n676), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n245), .B(new_n307), .C1(new_n677), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n631), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT103), .B(G1gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1324gat));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  NAND3_X1  g489(.A1(new_n686), .A2(new_n566), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n252), .B1(new_n686), .B2(new_n566), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT42), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(KEYINPUT42), .B2(new_n692), .ZN(G1325gat));
  INV_X1    g494(.A(new_n686), .ZN(new_n696));
  OAI21_X1  g495(.A(G15gat), .B1(new_n696), .B2(new_n624), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n643), .A2(G15gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n696), .B2(new_n698), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n686), .A2(new_n625), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  NOR3_X1   g501(.A1(new_n269), .A2(new_n306), .A3(new_n245), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n677), .B2(new_n685), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n275), .A3(new_n631), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(KEYINPUT45), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n706), .A2(KEYINPUT45), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n624), .A2(new_n632), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n648), .A2(new_n655), .B1(new_n710), .B2(new_n679), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n306), .A2(KEYINPUT44), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n709), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  AOI22_X1  g513(.A1(new_n642), .A2(new_n647), .B1(new_n654), .B2(KEYINPUT35), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n633), .A2(new_n580), .ZN(new_n716));
  OAI211_X1 g515(.A(KEYINPUT105), .B(new_n712), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT44), .B1(new_n656), .B2(new_n306), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n269), .B(KEYINPUT104), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n721), .A2(new_n676), .A3(new_n245), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n631), .ZN(new_n724));
  OAI21_X1  g523(.A(G29gat), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n707), .B1(new_n708), .B2(new_n725), .ZN(G1328gat));
  NAND3_X1  g525(.A1(new_n705), .A2(new_n276), .A3(new_n566), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n728));
  OAI21_X1  g527(.A(G36gat), .B1(new_n723), .B2(new_n646), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(G1329gat));
  NOR3_X1   g530(.A1(new_n656), .A2(KEYINPUT95), .A3(new_n676), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n683), .B1(new_n682), .B2(new_n684), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n703), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n643), .ZN(new_n735));
  INV_X1    g534(.A(new_n624), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G43gat), .ZN(new_n737));
  OAI22_X1  g536(.A1(new_n735), .A2(G43gat), .B1(new_n723), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g538(.A(KEYINPUT106), .B(G50gat), .C1(new_n723), .C2(new_n559), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n705), .A2(KEYINPUT107), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n559), .A2(new_n744), .A3(G50gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n740), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n740), .B2(new_n746), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(G1331gat));
  NAND3_X1  g549(.A1(new_n269), .A2(new_n676), .A3(new_n306), .ZN(new_n751));
  INV_X1    g550(.A(new_n245), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n710), .A2(new_n679), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n681), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n724), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT109), .B(G57gat), .Z(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1332gat));
  AOI211_X1 g559(.A(new_n646), .B(new_n757), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1333gat));
  NOR3_X1   g562(.A1(new_n757), .A2(G71gat), .A3(new_n643), .ZN(new_n764));
  INV_X1    g563(.A(new_n757), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n736), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n764), .B1(G71gat), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g567(.A1(new_n757), .A2(new_n559), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(new_n221), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n684), .A2(new_n269), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n245), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n720), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774), .B2(new_n724), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n756), .A2(new_n305), .A3(new_n771), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n778), .A2(new_n209), .A3(new_n631), .A4(new_n245), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n775), .A2(new_n779), .ZN(G1336gat));
  XOR2_X1   g579(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n781));
  NOR3_X1   g580(.A1(new_n752), .A2(G92gat), .A3(new_n646), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n646), .B(new_n772), .C1(new_n718), .C2(new_n719), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n210), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n720), .A2(new_n566), .A3(new_n773), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n782), .B(KEYINPUT110), .Z(new_n787));
  AOI22_X1  g586(.A1(new_n786), .A2(G92gat), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n788), .A2(KEYINPUT111), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n776), .A2(new_n777), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n787), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n784), .B2(new_n210), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n791), .B1(new_n795), .B2(KEYINPUT52), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n785), .B1(new_n790), .B2(new_n796), .ZN(G1337gat));
  NOR3_X1   g596(.A1(new_n752), .A2(G99gat), .A3(new_n643), .ZN(new_n798));
  XOR2_X1   g597(.A(new_n798), .B(KEYINPUT114), .Z(new_n799));
  NAND2_X1  g598(.A1(new_n778), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n774), .A2(new_n624), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(KEYINPUT113), .ZN(new_n802));
  OAI21_X1  g601(.A(G99gat), .B1(new_n801), .B2(KEYINPUT113), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(G1338gat));
  OAI21_X1  g603(.A(G106gat), .B1(new_n774), .B2(new_n559), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT115), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n752), .A2(G106gat), .A3(new_n559), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n778), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n809), .A3(KEYINPUT53), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n805), .B(new_n808), .C1(KEYINPUT115), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1339gat));
  NOR2_X1   g612(.A1(new_n751), .A2(new_n245), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n657), .A2(new_n658), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n663), .A2(new_n664), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n671), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n675), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT116), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n675), .A2(new_n821), .A3(new_n818), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n820), .A2(new_n305), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n230), .A2(new_n234), .A3(new_n204), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n242), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n240), .B1(new_n235), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n828), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n244), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n823), .A2(new_n824), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n305), .A3(new_n822), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT117), .B1(new_n836), .B2(new_n833), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n676), .A2(new_n833), .B1(new_n752), .B2(new_n819), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n835), .A2(new_n837), .B1(new_n306), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n815), .B1(new_n839), .B2(new_n721), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n644), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n724), .A2(new_n566), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(new_n467), .A3(new_n676), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n838), .A2(new_n306), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n824), .B1(new_n823), .B2(new_n834), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n836), .A2(KEYINPUT117), .A3(new_n833), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n721), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n814), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n651), .A2(new_n653), .ZN(new_n851));
  NOR4_X1   g650(.A1(new_n850), .A2(new_n724), .A3(new_n566), .A4(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n684), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n844), .A2(new_n853), .ZN(G1340gat));
  NOR3_X1   g653(.A1(new_n843), .A2(new_n465), .A3(new_n752), .ZN(new_n855));
  AOI21_X1  g654(.A(G120gat), .B1(new_n852), .B2(new_n245), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n843), .B2(new_n849), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n852), .A2(new_n250), .A3(new_n269), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1342gat));
  NAND3_X1  g659(.A1(new_n852), .A2(new_n472), .A3(new_n305), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n843), .B2(new_n306), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n842), .A2(new_n624), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n867), .B1(new_n850), .B2(new_n559), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n559), .A2(new_n867), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n839), .A2(new_n269), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n814), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n866), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n441), .B1(new_n872), .B2(new_n684), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n850), .A2(new_n724), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n624), .A2(new_n625), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n566), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n676), .A2(G141gat), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT118), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n874), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT58), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n840), .B2(new_n625), .ZN(new_n881));
  INV_X1    g680(.A(new_n869), .ZN(new_n882));
  INV_X1    g681(.A(new_n269), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n848), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n884), .B2(new_n815), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n624), .B(new_n842), .C1(new_n881), .C2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G141gat), .B1(new_n886), .B2(new_n676), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  INV_X1    g687(.A(new_n879), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n880), .A2(new_n890), .ZN(G1344gat));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n442), .A3(new_n245), .ZN(new_n894));
  AOI211_X1 g693(.A(KEYINPUT59), .B(new_n442), .C1(new_n872), .C2(new_n245), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n752), .B1(new_n866), .B2(KEYINPUT119), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n850), .A2(new_n882), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n823), .A2(new_n834), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n845), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n883), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n815), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n902), .B2(new_n625), .ZN(new_n903));
  OAI221_X1 g702(.A(new_n897), .B1(KEYINPUT119), .B2(new_n866), .C1(new_n898), .C2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n896), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n894), .B1(new_n895), .B2(new_n905), .ZN(G1345gat));
  AOI21_X1  g705(.A(new_n263), .B1(new_n872), .B2(new_n721), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n892), .A2(G155gat), .A3(new_n883), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT120), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G155gat), .B1(new_n886), .B2(new_n849), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n893), .A2(new_n263), .A3(new_n269), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n913), .ZN(G1346gat));
  AOI21_X1  g713(.A(new_n459), .B1(new_n893), .B2(new_n305), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n306), .A2(new_n439), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n872), .B2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n850), .A2(new_n631), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n851), .A2(new_n646), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(G169gat), .B1(new_n921), .B2(new_n684), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n646), .A2(new_n631), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n841), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n311), .A3(new_n676), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n922), .A2(new_n925), .ZN(G1348gat));
  OAI21_X1  g725(.A(G176gat), .B1(new_n924), .B2(new_n752), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n918), .A2(new_n312), .A3(new_n245), .A4(new_n919), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(KEYINPUT121), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1349gat));
  NAND3_X1  g732(.A1(new_n841), .A2(new_n721), .A3(new_n923), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G183gat), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n269), .A2(new_n327), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n920), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT60), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n920), .A2(new_n938), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n941), .A2(new_n935), .A3(new_n937), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n940), .A2(new_n943), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n921), .A2(new_n338), .A3(new_n305), .ZN(new_n945));
  OAI21_X1  g744(.A(G190gat), .B1(new_n924), .B2(new_n306), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(KEYINPUT61), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(KEYINPUT61), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1351gat));
  NAND2_X1  g748(.A1(new_n902), .A2(new_n625), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n867), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n840), .A2(new_n869), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT123), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n954), .B1(new_n898), .B2(new_n903), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n624), .A2(new_n923), .ZN(new_n956));
  INV_X1    g755(.A(G197gat), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n676), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n953), .A2(new_n955), .A3(new_n956), .A4(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n875), .A2(new_n646), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n918), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n961), .B2(new_n676), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n959), .A2(new_n962), .ZN(G1352gat));
  XNOR2_X1  g762(.A(KEYINPUT124), .B(G204gat), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n752), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n752), .A2(new_n964), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n918), .A2(new_n960), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n968), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n968), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n966), .A2(new_n972), .A3(new_n973), .ZN(G1353gat));
  INV_X1    g773(.A(G211gat), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n918), .A2(new_n975), .A3(new_n269), .A4(new_n960), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n956), .A2(new_n269), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n977), .B1(new_n951), .B2(new_n952), .ZN(new_n978));
  OAI21_X1  g777(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT63), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NOR4_X1   g783(.A1(new_n978), .A2(new_n981), .A3(new_n982), .A4(new_n975), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n976), .B1(new_n984), .B2(new_n985), .ZN(G1354gat));
  INV_X1    g785(.A(G218gat), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n306), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n953), .A2(new_n955), .A3(new_n956), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n987), .B1(new_n961), .B2(new_n306), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n989), .A2(new_n990), .ZN(G1355gat));
endmodule


