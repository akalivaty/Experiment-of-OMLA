

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U548 ( .A(KEYINPUT31), .ZN(n687) );
  XOR2_X1 U549 ( .A(n679), .B(KEYINPUT92), .Z(n754) );
  XOR2_X1 U550 ( .A(n532), .B(KEYINPUT1), .Z(n635) );
  NOR2_X1 U551 ( .A1(G651), .A2(n628), .ZN(n642) );
  NOR2_X1 U552 ( .A1(n522), .A2(n521), .ZN(G160) );
  INV_X1 U553 ( .A(G2105), .ZN(n513) );
  XNOR2_X1 U554 ( .A(G2104), .B(KEYINPUT66), .ZN(n512) );
  NAND2_X1 U555 ( .A1(n513), .A2(n512), .ZN(n510) );
  XNOR2_X2 U556 ( .A(KEYINPUT67), .B(n510), .ZN(n880) );
  NAND2_X1 U557 ( .A1(n880), .A2(G101), .ZN(n511) );
  XOR2_X1 U558 ( .A(n511), .B(KEYINPUT23), .Z(n515) );
  NOR2_X1 U559 ( .A1(n513), .A2(n512), .ZN(n882) );
  NAND2_X1 U560 ( .A1(n882), .A2(G125), .ZN(n514) );
  NAND2_X1 U561 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U562 ( .A(n516), .B(KEYINPUT68), .ZN(n522) );
  AND2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  NAND2_X1 U564 ( .A1(n884), .A2(G113), .ZN(n519) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XOR2_X1 U566 ( .A(KEYINPUT17), .B(n517), .Z(n889) );
  NAND2_X1 U567 ( .A1(n889), .A2(G137), .ZN(n518) );
  NAND2_X1 U568 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U569 ( .A(KEYINPUT69), .B(n520), .Z(n521) );
  XOR2_X1 U570 ( .A(G2443), .B(G2446), .Z(n524) );
  XNOR2_X1 U571 ( .A(G2427), .B(G2451), .ZN(n523) );
  XNOR2_X1 U572 ( .A(n524), .B(n523), .ZN(n530) );
  XOR2_X1 U573 ( .A(G2430), .B(G2454), .Z(n526) );
  XNOR2_X1 U574 ( .A(G1348), .B(G1341), .ZN(n525) );
  XNOR2_X1 U575 ( .A(n526), .B(n525), .ZN(n528) );
  XOR2_X1 U576 ( .A(G2435), .B(G2438), .Z(n527) );
  XNOR2_X1 U577 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U578 ( .A(n530), .B(n529), .Z(n531) );
  AND2_X1 U579 ( .A1(G14), .A2(n531), .ZN(G401) );
  XOR2_X1 U580 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  NAND2_X1 U581 ( .A1(G52), .A2(n642), .ZN(n534) );
  INV_X1 U582 ( .A(G651), .ZN(n535) );
  NOR2_X1 U583 ( .A1(n535), .A2(G543), .ZN(n532) );
  NAND2_X1 U584 ( .A1(G64), .A2(n635), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n540) );
  NOR2_X1 U586 ( .A1(n628), .A2(n535), .ZN(n638) );
  NAND2_X1 U587 ( .A1(G77), .A2(n638), .ZN(n537) );
  NOR2_X1 U588 ( .A1(G543), .A2(G651), .ZN(n634) );
  NAND2_X1 U589 ( .A1(G90), .A2(n634), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U591 ( .A(KEYINPUT9), .B(n538), .Z(n539) );
  NOR2_X1 U592 ( .A1(n540), .A2(n539), .ZN(G171) );
  AND2_X1 U593 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U594 ( .A(G57), .ZN(G237) );
  INV_X1 U595 ( .A(G108), .ZN(G238) );
  INV_X1 U596 ( .A(G69), .ZN(G235) );
  INV_X1 U597 ( .A(G132), .ZN(G219) );
  INV_X1 U598 ( .A(G82), .ZN(G220) );
  NAND2_X1 U599 ( .A1(G51), .A2(n642), .ZN(n542) );
  NAND2_X1 U600 ( .A1(G63), .A2(n635), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U602 ( .A(KEYINPUT6), .B(n543), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G89), .A2(n634), .ZN(n544) );
  XNOR2_X1 U604 ( .A(n544), .B(KEYINPUT4), .ZN(n545) );
  XNOR2_X1 U605 ( .A(n545), .B(KEYINPUT76), .ZN(n547) );
  NAND2_X1 U606 ( .A1(G76), .A2(n638), .ZN(n546) );
  NAND2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U608 ( .A(n548), .B(KEYINPUT5), .Z(n549) );
  NOR2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U610 ( .A(KEYINPUT7), .B(n551), .Z(n552) );
  XOR2_X1 U611 ( .A(KEYINPUT77), .B(n552), .Z(G168) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(n553) );
  XNOR2_X1 U613 ( .A(KEYINPUT78), .B(n553), .ZN(G286) );
  NAND2_X1 U614 ( .A1(G7), .A2(G661), .ZN(n554) );
  XOR2_X1 U615 ( .A(n554), .B(KEYINPUT10), .Z(n828) );
  NAND2_X1 U616 ( .A1(n828), .A2(G567), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT11), .B(n555), .Z(G234) );
  XOR2_X1 U618 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n557) );
  NAND2_X1 U619 ( .A1(G56), .A2(n635), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n557), .B(n556), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n634), .A2(G81), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n558), .B(KEYINPUT12), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G68), .A2(n638), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n561), .B(KEYINPUT13), .ZN(n562) );
  XNOR2_X1 U626 ( .A(KEYINPUT73), .B(n562), .ZN(n563) );
  NOR2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U628 ( .A(KEYINPUT74), .B(n565), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G43), .A2(n642), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n997) );
  INV_X1 U631 ( .A(n997), .ZN(n902) );
  NAND2_X1 U632 ( .A1(n902), .A2(G860), .ZN(G153) );
  INV_X1 U633 ( .A(G171), .ZN(G301) );
  NAND2_X1 U634 ( .A1(G868), .A2(G301), .ZN(n577) );
  NAND2_X1 U635 ( .A1(G66), .A2(n635), .ZN(n574) );
  NAND2_X1 U636 ( .A1(G79), .A2(n638), .ZN(n569) );
  NAND2_X1 U637 ( .A1(G92), .A2(n634), .ZN(n568) );
  NAND2_X1 U638 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U639 ( .A1(G54), .A2(n642), .ZN(n570) );
  XNOR2_X1 U640 ( .A(KEYINPUT75), .B(n570), .ZN(n571) );
  NOR2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U643 ( .A(n575), .B(KEYINPUT15), .Z(n992) );
  INV_X1 U644 ( .A(G868), .ZN(n652) );
  NAND2_X1 U645 ( .A1(n992), .A2(n652), .ZN(n576) );
  NAND2_X1 U646 ( .A1(n577), .A2(n576), .ZN(G284) );
  NAND2_X1 U647 ( .A1(G91), .A2(n634), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G65), .A2(n635), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G78), .A2(n638), .ZN(n580) );
  XNOR2_X1 U651 ( .A(KEYINPUT71), .B(n580), .ZN(n581) );
  NOR2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n642), .A2(G53), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n584), .A2(n583), .ZN(G299) );
  XOR2_X1 U655 ( .A(KEYINPUT79), .B(n652), .Z(n585) );
  NOR2_X1 U656 ( .A1(G286), .A2(n585), .ZN(n587) );
  NOR2_X1 U657 ( .A1(G868), .A2(G299), .ZN(n586) );
  NOR2_X1 U658 ( .A1(n587), .A2(n586), .ZN(G297) );
  INV_X1 U659 ( .A(G860), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n588), .A2(G559), .ZN(n589) );
  INV_X1 U661 ( .A(n992), .ZN(n609) );
  NAND2_X1 U662 ( .A1(n589), .A2(n609), .ZN(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U664 ( .A1(n609), .A2(G868), .ZN(n591) );
  NOR2_X1 U665 ( .A1(G559), .A2(n591), .ZN(n593) );
  NOR2_X1 U666 ( .A1(G868), .A2(n997), .ZN(n592) );
  NOR2_X1 U667 ( .A1(n593), .A2(n592), .ZN(G282) );
  NAND2_X1 U668 ( .A1(G111), .A2(n884), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G135), .A2(n889), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G123), .A2(n882), .ZN(n596) );
  XNOR2_X1 U672 ( .A(n596), .B(KEYINPUT18), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n880), .A2(G99), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n952) );
  XNOR2_X1 U676 ( .A(n952), .B(G2096), .ZN(n601) );
  INV_X1 U677 ( .A(G2100), .ZN(n841) );
  NAND2_X1 U678 ( .A1(n601), .A2(n841), .ZN(G156) );
  NAND2_X1 U679 ( .A1(G80), .A2(n638), .ZN(n603) );
  NAND2_X1 U680 ( .A1(G93), .A2(n634), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n608) );
  NAND2_X1 U682 ( .A1(G55), .A2(n642), .ZN(n605) );
  NAND2_X1 U683 ( .A1(G67), .A2(n635), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U685 ( .A(KEYINPUT81), .B(n606), .Z(n607) );
  OR2_X1 U686 ( .A1(n608), .A2(n607), .ZN(n653) );
  NAND2_X1 U687 ( .A1(G559), .A2(n609), .ZN(n610) );
  XNOR2_X1 U688 ( .A(n997), .B(n610), .ZN(n650) );
  XNOR2_X1 U689 ( .A(KEYINPUT80), .B(n650), .ZN(n611) );
  NOR2_X1 U690 ( .A1(G860), .A2(n611), .ZN(n612) );
  XOR2_X1 U691 ( .A(n653), .B(n612), .Z(G145) );
  NAND2_X1 U692 ( .A1(G75), .A2(n638), .ZN(n614) );
  NAND2_X1 U693 ( .A1(G88), .A2(n634), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G50), .A2(n642), .ZN(n616) );
  NAND2_X1 U696 ( .A1(G62), .A2(n635), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U698 ( .A1(n618), .A2(n617), .ZN(G166) );
  INV_X1 U699 ( .A(G166), .ZN(G303) );
  NAND2_X1 U700 ( .A1(G85), .A2(n634), .ZN(n620) );
  NAND2_X1 U701 ( .A1(G60), .A2(n635), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n638), .A2(G72), .ZN(n621) );
  XOR2_X1 U704 ( .A(KEYINPUT70), .B(n621), .Z(n622) );
  NOR2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n642), .A2(G47), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(G290) );
  NAND2_X1 U708 ( .A1(G49), .A2(n642), .ZN(n627) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n628), .A2(G87), .ZN(n629) );
  XOR2_X1 U712 ( .A(KEYINPUT82), .B(n629), .Z(n630) );
  NOR2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n633) );
  INV_X1 U714 ( .A(n635), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U716 ( .A1(G86), .A2(n634), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G61), .A2(n635), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G73), .A2(n638), .ZN(n639) );
  XOR2_X1 U720 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U721 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n642), .A2(G48), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(G305) );
  XOR2_X1 U724 ( .A(G303), .B(KEYINPUT19), .Z(n649) );
  XOR2_X1 U725 ( .A(n653), .B(G299), .Z(n645) );
  XNOR2_X1 U726 ( .A(n645), .B(G290), .ZN(n646) );
  XNOR2_X1 U727 ( .A(n646), .B(G288), .ZN(n647) );
  XNOR2_X1 U728 ( .A(n647), .B(G305), .ZN(n648) );
  XNOR2_X1 U729 ( .A(n649), .B(n648), .ZN(n901) );
  XOR2_X1 U730 ( .A(n901), .B(n650), .Z(n651) );
  NAND2_X1 U731 ( .A1(G868), .A2(n651), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(G295) );
  NAND2_X1 U734 ( .A1(G2078), .A2(G2084), .ZN(n656) );
  XOR2_X1 U735 ( .A(KEYINPUT20), .B(n656), .Z(n657) );
  NAND2_X1 U736 ( .A1(G2090), .A2(n657), .ZN(n658) );
  XNOR2_X1 U737 ( .A(KEYINPUT21), .B(n658), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n659), .A2(G2072), .ZN(n660) );
  XOR2_X1 U739 ( .A(KEYINPUT83), .B(n660), .Z(G158) );
  XNOR2_X1 U740 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U741 ( .A1(G483), .A2(G661), .ZN(n670) );
  NOR2_X1 U742 ( .A1(G220), .A2(G219), .ZN(n661) );
  XOR2_X1 U743 ( .A(KEYINPUT22), .B(n661), .Z(n662) );
  NOR2_X1 U744 ( .A1(G218), .A2(n662), .ZN(n663) );
  NAND2_X1 U745 ( .A1(G96), .A2(n663), .ZN(n833) );
  NAND2_X1 U746 ( .A1(G2106), .A2(n833), .ZN(n664) );
  XNOR2_X1 U747 ( .A(n664), .B(KEYINPUT84), .ZN(n669) );
  NOR2_X1 U748 ( .A1(G235), .A2(G238), .ZN(n665) );
  NAND2_X1 U749 ( .A1(G120), .A2(n665), .ZN(n666) );
  NOR2_X1 U750 ( .A1(n666), .A2(G237), .ZN(n667) );
  XNOR2_X1 U751 ( .A(n667), .B(KEYINPUT85), .ZN(n834) );
  NAND2_X1 U752 ( .A1(G567), .A2(n834), .ZN(n668) );
  NAND2_X1 U753 ( .A1(n669), .A2(n668), .ZN(n856) );
  NOR2_X1 U754 ( .A1(n670), .A2(n856), .ZN(n671) );
  XNOR2_X1 U755 ( .A(n671), .B(KEYINPUT86), .ZN(n832) );
  NAND2_X1 U756 ( .A1(G36), .A2(n832), .ZN(G176) );
  NAND2_X1 U757 ( .A1(G102), .A2(n880), .ZN(n673) );
  NAND2_X1 U758 ( .A1(G138), .A2(n889), .ZN(n672) );
  NAND2_X1 U759 ( .A1(n673), .A2(n672), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G126), .A2(n882), .ZN(n675) );
  NAND2_X1 U761 ( .A1(G114), .A2(n884), .ZN(n674) );
  NAND2_X1 U762 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U763 ( .A1(n677), .A2(n676), .ZN(G164) );
  NAND2_X1 U764 ( .A1(G160), .A2(G40), .ZN(n775) );
  NOR2_X1 U765 ( .A1(G1384), .A2(G164), .ZN(n678) );
  XOR2_X1 U766 ( .A(n678), .B(KEYINPUT64), .Z(n776) );
  NOR2_X4 U767 ( .A1(n775), .A2(n776), .ZN(n703) );
  INV_X1 U768 ( .A(n703), .ZN(n721) );
  NAND2_X1 U769 ( .A1(n721), .A2(G8), .ZN(n679) );
  INV_X1 U770 ( .A(n754), .ZN(n720) );
  NOR2_X1 U771 ( .A1(n720), .A2(G1966), .ZN(n741) );
  NOR2_X1 U772 ( .A1(G2084), .A2(n721), .ZN(n734) );
  NOR2_X1 U773 ( .A1(n741), .A2(n734), .ZN(n680) );
  NAND2_X1 U774 ( .A1(G8), .A2(n680), .ZN(n681) );
  XNOR2_X1 U775 ( .A(KEYINPUT30), .B(n681), .ZN(n682) );
  NOR2_X1 U776 ( .A1(G168), .A2(n682), .ZN(n686) );
  XNOR2_X1 U777 ( .A(G2078), .B(KEYINPUT25), .ZN(n975) );
  NOR2_X1 U778 ( .A1(n721), .A2(n975), .ZN(n684) );
  INV_X1 U779 ( .A(G1961), .ZN(n846) );
  NOR2_X1 U780 ( .A1(n703), .A2(n846), .ZN(n683) );
  NOR2_X1 U781 ( .A1(n684), .A2(n683), .ZN(n689) );
  NOR2_X1 U782 ( .A1(G171), .A2(n689), .ZN(n685) );
  NOR2_X1 U783 ( .A1(n686), .A2(n685), .ZN(n688) );
  XNOR2_X1 U784 ( .A(n688), .B(n687), .ZN(n737) );
  AND2_X1 U785 ( .A1(G171), .A2(n689), .ZN(n690) );
  XOR2_X1 U786 ( .A(KEYINPUT94), .B(n690), .Z(n719) );
  NAND2_X1 U787 ( .A1(n703), .A2(G2072), .ZN(n692) );
  XOR2_X1 U788 ( .A(KEYINPUT95), .B(KEYINPUT27), .Z(n691) );
  XOR2_X1 U789 ( .A(n692), .B(n691), .Z(n695) );
  XOR2_X1 U790 ( .A(KEYINPUT96), .B(G1956), .Z(n917) );
  NOR2_X1 U791 ( .A1(n703), .A2(n917), .ZN(n693) );
  XNOR2_X1 U792 ( .A(KEYINPUT97), .B(n693), .ZN(n694) );
  NAND2_X1 U793 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U794 ( .A1(G299), .A2(n697), .ZN(n696) );
  XNOR2_X1 U795 ( .A(n696), .B(KEYINPUT28), .ZN(n716) );
  NOR2_X1 U796 ( .A1(G299), .A2(n697), .ZN(n698) );
  XNOR2_X1 U797 ( .A(KEYINPUT99), .B(n698), .ZN(n714) );
  NAND2_X1 U798 ( .A1(G2067), .A2(n703), .ZN(n700) );
  NAND2_X1 U799 ( .A1(G1348), .A2(n721), .ZN(n699) );
  NAND2_X1 U800 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U801 ( .A1(n992), .A2(n701), .ZN(n712) );
  OR2_X1 U802 ( .A1(n992), .A2(n701), .ZN(n710) );
  NAND2_X1 U803 ( .A1(G1341), .A2(n721), .ZN(n702) );
  XOR2_X1 U804 ( .A(KEYINPUT98), .B(n702), .Z(n707) );
  XOR2_X1 U805 ( .A(KEYINPUT65), .B(KEYINPUT26), .Z(n705) );
  NAND2_X1 U806 ( .A1(G1996), .A2(n703), .ZN(n704) );
  XOR2_X1 U807 ( .A(n705), .B(n704), .Z(n706) );
  NOR2_X1 U808 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U809 ( .A1(n708), .A2(n902), .ZN(n709) );
  NAND2_X1 U810 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U811 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U812 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U813 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U814 ( .A(KEYINPUT29), .B(n717), .Z(n718) );
  NAND2_X1 U815 ( .A1(n719), .A2(n718), .ZN(n736) );
  INV_X1 U816 ( .A(G8), .ZN(n726) );
  NOR2_X1 U817 ( .A1(n720), .A2(G1971), .ZN(n723) );
  NOR2_X1 U818 ( .A1(G2090), .A2(n721), .ZN(n722) );
  NOR2_X1 U819 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U820 ( .A1(n724), .A2(G303), .ZN(n725) );
  OR2_X1 U821 ( .A1(n726), .A2(n725), .ZN(n728) );
  AND2_X1 U822 ( .A1(n736), .A2(n728), .ZN(n727) );
  NAND2_X1 U823 ( .A1(n737), .A2(n727), .ZN(n732) );
  INV_X1 U824 ( .A(n728), .ZN(n730) );
  AND2_X1 U825 ( .A1(G286), .A2(G8), .ZN(n729) );
  OR2_X1 U826 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U827 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U828 ( .A(KEYINPUT32), .B(n733), .Z(n743) );
  NAND2_X1 U829 ( .A1(G8), .A2(n734), .ZN(n735) );
  XOR2_X1 U830 ( .A(KEYINPUT93), .B(n735), .Z(n739) );
  NAND2_X1 U831 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U833 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U834 ( .A1(n743), .A2(n742), .ZN(n747) );
  NAND2_X1 U835 ( .A1(G166), .A2(G8), .ZN(n744) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n744), .ZN(n745) );
  NOR2_X1 U837 ( .A1(n747), .A2(n745), .ZN(n746) );
  OR2_X1 U838 ( .A1(n746), .A2(n754), .ZN(n774) );
  INV_X1 U839 ( .A(n747), .ZN(n763) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U842 ( .A1(n749), .A2(n748), .ZN(n1007) );
  XNOR2_X1 U843 ( .A(KEYINPUT100), .B(n1007), .ZN(n761) );
  XOR2_X1 U844 ( .A(n749), .B(KEYINPUT101), .Z(n750) );
  NAND2_X1 U845 ( .A1(n750), .A2(n754), .ZN(n753) );
  XNOR2_X1 U846 ( .A(KEYINPUT102), .B(G1981), .ZN(n751) );
  XOR2_X1 U847 ( .A(n751), .B(G305), .Z(n988) );
  AND2_X1 U848 ( .A1(KEYINPUT33), .A2(n988), .ZN(n752) );
  NAND2_X1 U849 ( .A1(n753), .A2(n752), .ZN(n757) );
  INV_X1 U850 ( .A(n757), .ZN(n755) );
  OR2_X1 U851 ( .A1(n755), .A2(n754), .ZN(n767) );
  INV_X1 U852 ( .A(n767), .ZN(n760) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n756) );
  XOR2_X1 U854 ( .A(n756), .B(KEYINPUT24), .Z(n758) );
  AND2_X1 U855 ( .A1(n758), .A2(n757), .ZN(n759) );
  OR2_X1 U856 ( .A1(n760), .A2(n759), .ZN(n764) );
  AND2_X1 U857 ( .A1(n761), .A2(n764), .ZN(n762) );
  NAND2_X1 U858 ( .A1(n763), .A2(n762), .ZN(n772) );
  INV_X1 U859 ( .A(n764), .ZN(n770) );
  NAND2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n1004) );
  NAND2_X1 U861 ( .A1(n1004), .A2(n988), .ZN(n766) );
  OR2_X1 U862 ( .A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(n765) );
  NOR2_X1 U863 ( .A1(n766), .A2(n765), .ZN(n768) );
  AND2_X1 U864 ( .A1(n768), .A2(n767), .ZN(n769) );
  OR2_X1 U865 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U866 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n812) );
  XNOR2_X1 U868 ( .A(G1986), .B(G290), .ZN(n994) );
  INV_X1 U869 ( .A(n775), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n777), .A2(n776), .ZN(n795) );
  INV_X1 U871 ( .A(n795), .ZN(n823) );
  AND2_X1 U872 ( .A1(n994), .A2(n823), .ZN(n810) );
  NAND2_X1 U873 ( .A1(n880), .A2(G95), .ZN(n779) );
  NAND2_X1 U874 ( .A1(n889), .A2(G131), .ZN(n778) );
  NAND2_X1 U875 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U876 ( .A(KEYINPUT90), .B(n780), .Z(n784) );
  NAND2_X1 U877 ( .A1(G119), .A2(n882), .ZN(n782) );
  NAND2_X1 U878 ( .A1(G107), .A2(n884), .ZN(n781) );
  AND2_X1 U879 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U880 ( .A1(n784), .A2(n783), .ZN(n894) );
  AND2_X1 U881 ( .A1(n894), .A2(G1991), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G129), .A2(n882), .ZN(n786) );
  NAND2_X1 U883 ( .A1(G117), .A2(n884), .ZN(n785) );
  NAND2_X1 U884 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U885 ( .A1(n880), .A2(G105), .ZN(n787) );
  XOR2_X1 U886 ( .A(KEYINPUT38), .B(n787), .Z(n788) );
  NOR2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U888 ( .A(KEYINPUT91), .B(n790), .Z(n792) );
  NAND2_X1 U889 ( .A1(n889), .A2(G141), .ZN(n791) );
  NAND2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n897) );
  AND2_X1 U891 ( .A1(n897), .A2(G1996), .ZN(n793) );
  NOR2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n938) );
  NOR2_X1 U893 ( .A1(n938), .A2(n795), .ZN(n815) );
  INV_X1 U894 ( .A(n815), .ZN(n808) );
  XOR2_X1 U895 ( .A(G2067), .B(KEYINPUT37), .Z(n796) );
  XNOR2_X1 U896 ( .A(KEYINPUT87), .B(n796), .ZN(n820) );
  XNOR2_X1 U897 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n807) );
  NAND2_X1 U898 ( .A1(G128), .A2(n882), .ZN(n798) );
  NAND2_X1 U899 ( .A1(G116), .A2(n884), .ZN(n797) );
  NAND2_X1 U900 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U901 ( .A(KEYINPUT35), .B(n799), .ZN(n805) );
  NAND2_X1 U902 ( .A1(G104), .A2(n880), .ZN(n801) );
  NAND2_X1 U903 ( .A1(G140), .A2(n889), .ZN(n800) );
  NAND2_X1 U904 ( .A1(n801), .A2(n800), .ZN(n803) );
  XOR2_X1 U905 ( .A(KEYINPUT34), .B(KEYINPUT88), .Z(n802) );
  XNOR2_X1 U906 ( .A(n803), .B(n802), .ZN(n804) );
  NAND2_X1 U907 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U908 ( .A(n807), .B(n806), .ZN(n876) );
  NOR2_X1 U909 ( .A1(n820), .A2(n876), .ZN(n956) );
  NAND2_X1 U910 ( .A1(n823), .A2(n956), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n808), .A2(n818), .ZN(n809) );
  NOR2_X1 U912 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U913 ( .A1(n812), .A2(n811), .ZN(n826) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n897), .ZN(n946) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n894), .ZN(n953) );
  NOR2_X1 U917 ( .A1(n813), .A2(n953), .ZN(n814) );
  NOR2_X1 U918 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U919 ( .A1(n946), .A2(n816), .ZN(n817) );
  XNOR2_X1 U920 ( .A(KEYINPUT39), .B(n817), .ZN(n819) );
  NAND2_X1 U921 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U922 ( .A1(n820), .A2(n876), .ZN(n954) );
  NAND2_X1 U923 ( .A1(n821), .A2(n954), .ZN(n822) );
  NAND2_X1 U924 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U925 ( .A(KEYINPUT103), .B(n824), .Z(n825) );
  NAND2_X1 U926 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U927 ( .A(KEYINPUT40), .B(n827), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n828), .ZN(G217) );
  INV_X1 U929 ( .A(n828), .ZN(G223) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n829) );
  XOR2_X1 U931 ( .A(KEYINPUT104), .B(n829), .Z(n830) );
  NAND2_X1 U932 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U934 ( .A1(n832), .A2(n831), .ZN(G188) );
  XNOR2_X1 U935 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  XOR2_X1 U936 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  NOR2_X1 U937 ( .A1(n834), .A2(n833), .ZN(G325) );
  XNOR2_X1 U938 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2678), .Z(n836) );
  XNOR2_X1 U941 ( .A(KEYINPUT110), .B(KEYINPUT109), .ZN(n835) );
  XNOR2_X1 U942 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U943 ( .A(KEYINPUT42), .B(G2090), .Z(n838) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n837) );
  XNOR2_X1 U945 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U946 ( .A(n840), .B(n839), .Z(n843) );
  XOR2_X1 U947 ( .A(G2096), .B(n841), .Z(n842) );
  XNOR2_X1 U948 ( .A(n843), .B(n842), .ZN(n845) );
  XOR2_X1 U949 ( .A(G2078), .B(G2084), .Z(n844) );
  XNOR2_X1 U950 ( .A(n845), .B(n844), .ZN(G227) );
  XNOR2_X1 U951 ( .A(n846), .B(G1956), .ZN(n848) );
  XNOR2_X1 U952 ( .A(G1981), .B(G1966), .ZN(n847) );
  XNOR2_X1 U953 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U954 ( .A(n849), .B(G2474), .Z(n851) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U956 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U957 ( .A(KEYINPUT41), .B(G1986), .Z(n853) );
  XNOR2_X1 U958 ( .A(G1976), .B(G1971), .ZN(n852) );
  XNOR2_X1 U959 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U960 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U961 ( .A(KEYINPUT108), .B(n856), .Z(G319) );
  NAND2_X1 U962 ( .A1(G112), .A2(n884), .ZN(n858) );
  NAND2_X1 U963 ( .A1(G136), .A2(n889), .ZN(n857) );
  NAND2_X1 U964 ( .A1(n858), .A2(n857), .ZN(n863) );
  NAND2_X1 U965 ( .A1(G124), .A2(n882), .ZN(n859) );
  XNOR2_X1 U966 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U967 ( .A1(n880), .A2(G100), .ZN(n860) );
  NAND2_X1 U968 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U969 ( .A1(n863), .A2(n862), .ZN(G162) );
  XOR2_X1 U970 ( .A(KEYINPUT48), .B(KEYINPUT115), .Z(n865) );
  XNOR2_X1 U971 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n864) );
  XNOR2_X1 U972 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U973 ( .A(n866), .B(n952), .Z(n868) );
  XNOR2_X1 U974 ( .A(G164), .B(G162), .ZN(n867) );
  XNOR2_X1 U975 ( .A(n868), .B(n867), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G130), .A2(n882), .ZN(n870) );
  NAND2_X1 U977 ( .A1(G118), .A2(n884), .ZN(n869) );
  NAND2_X1 U978 ( .A1(n870), .A2(n869), .ZN(n875) );
  NAND2_X1 U979 ( .A1(G106), .A2(n880), .ZN(n872) );
  NAND2_X1 U980 ( .A1(G142), .A2(n889), .ZN(n871) );
  NAND2_X1 U981 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U982 ( .A(n873), .B(KEYINPUT45), .Z(n874) );
  NOR2_X1 U983 ( .A1(n875), .A2(n874), .ZN(n877) );
  XNOR2_X1 U984 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U985 ( .A(n879), .B(n878), .Z(n896) );
  NAND2_X1 U986 ( .A1(n880), .A2(G103), .ZN(n881) );
  XNOR2_X1 U987 ( .A(KEYINPUT111), .B(n881), .ZN(n893) );
  NAND2_X1 U988 ( .A1(n882), .A2(G127), .ZN(n883) );
  XNOR2_X1 U989 ( .A(n883), .B(KEYINPUT112), .ZN(n886) );
  NAND2_X1 U990 ( .A1(G115), .A2(n884), .ZN(n885) );
  NAND2_X1 U991 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U992 ( .A(KEYINPUT113), .B(n887), .Z(n888) );
  XNOR2_X1 U993 ( .A(n888), .B(KEYINPUT47), .ZN(n891) );
  NAND2_X1 U994 ( .A1(G139), .A2(n889), .ZN(n890) );
  NAND2_X1 U995 ( .A1(n891), .A2(n890), .ZN(n892) );
  NOR2_X1 U996 ( .A1(n893), .A2(n892), .ZN(n941) );
  XOR2_X1 U997 ( .A(n894), .B(n941), .Z(n895) );
  XNOR2_X1 U998 ( .A(n896), .B(n895), .ZN(n899) );
  XOR2_X1 U999 ( .A(G160), .B(n897), .Z(n898) );
  XNOR2_X1 U1000 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n900), .ZN(G395) );
  XNOR2_X1 U1002 ( .A(G286), .B(n901), .ZN(n904) );
  XOR2_X1 U1003 ( .A(n992), .B(n902), .Z(n903) );
  XNOR2_X1 U1004 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(n905), .B(G171), .Z(n906) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n906), .ZN(G397) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n907) );
  XOR2_X1 U1008 ( .A(KEYINPUT49), .B(n907), .Z(n908) );
  NAND2_X1 U1009 ( .A1(n908), .A2(G319), .ZN(n909) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n909), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(KEYINPUT116), .B(n910), .ZN(n912) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1015 ( .A(G5), .B(G1961), .Z(n933) );
  XOR2_X1 U1016 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n924) );
  XNOR2_X1 U1017 ( .A(G1981), .B(G6), .ZN(n914) );
  XNOR2_X1 U1018 ( .A(G1341), .B(G19), .ZN(n913) );
  NOR2_X1 U1019 ( .A1(n914), .A2(n913), .ZN(n922) );
  XOR2_X1 U1020 ( .A(KEYINPUT126), .B(G4), .Z(n916) );
  XNOR2_X1 U1021 ( .A(G1348), .B(KEYINPUT59), .ZN(n915) );
  XNOR2_X1 U1022 ( .A(n916), .B(n915), .ZN(n920) );
  XNOR2_X1 U1023 ( .A(G20), .B(n917), .ZN(n918) );
  XNOR2_X1 U1024 ( .A(KEYINPUT125), .B(n918), .ZN(n919) );
  NOR2_X1 U1025 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1026 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1027 ( .A(n924), .B(n923), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(G1976), .B(G23), .ZN(n926) );
  XNOR2_X1 U1029 ( .A(G1971), .B(G22), .ZN(n925) );
  NOR2_X1 U1030 ( .A1(n926), .A2(n925), .ZN(n928) );
  XOR2_X1 U1031 ( .A(G1986), .B(G24), .Z(n927) );
  NAND2_X1 U1032 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1033 ( .A(KEYINPUT58), .B(n929), .ZN(n930) );
  NOR2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(G21), .B(G1966), .ZN(n934) );
  NOR2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1038 ( .A(KEYINPUT61), .B(n936), .Z(n937) );
  NOR2_X1 U1039 ( .A1(G16), .A2(n937), .ZN(n1019) );
  INV_X1 U1040 ( .A(KEYINPUT55), .ZN(n963) );
  XOR2_X1 U1041 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n961) );
  XNOR2_X1 U1042 ( .A(G160), .B(G2084), .ZN(n939) );
  NAND2_X1 U1043 ( .A1(n939), .A2(n938), .ZN(n951) );
  XOR2_X1 U1044 ( .A(G2072), .B(KEYINPUT117), .Z(n940) );
  XOR2_X1 U1045 ( .A(n941), .B(n940), .Z(n943) );
  XOR2_X1 U1046 ( .A(G164), .B(G2078), .Z(n942) );
  NOR2_X1 U1047 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1048 ( .A(KEYINPUT50), .B(n944), .ZN(n949) );
  XOR2_X1 U1049 ( .A(G2090), .B(G162), .Z(n945) );
  NOR2_X1 U1050 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1051 ( .A(KEYINPUT51), .B(n947), .Z(n948) );
  NAND2_X1 U1052 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1053 ( .A1(n951), .A2(n950), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n953), .A2(n952), .ZN(n955) );
  NAND2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(n961), .B(n960), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1060 ( .A1(n964), .A2(G29), .ZN(n1017) );
  XNOR2_X1 U1061 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(n965), .B(G34), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(G2084), .B(n966), .ZN(n983) );
  XNOR2_X1 U1064 ( .A(G2090), .B(G35), .ZN(n981) );
  XNOR2_X1 U1065 ( .A(G1991), .B(G25), .ZN(n968) );
  XNOR2_X1 U1066 ( .A(G33), .B(G2072), .ZN(n967) );
  NOR2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n974) );
  XOR2_X1 U1068 ( .A(G2067), .B(G26), .Z(n969) );
  NAND2_X1 U1069 ( .A1(n969), .A2(G28), .ZN(n972) );
  XNOR2_X1 U1070 ( .A(G32), .B(G1996), .ZN(n970) );
  XNOR2_X1 U1071 ( .A(KEYINPUT120), .B(n970), .ZN(n971) );
  NOR2_X1 U1072 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1073 ( .A1(n974), .A2(n973), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(G27), .B(n975), .ZN(n976) );
  XNOR2_X1 U1075 ( .A(KEYINPUT119), .B(n976), .ZN(n977) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1077 ( .A(KEYINPUT53), .B(n979), .ZN(n980) );
  NOR2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1080 ( .A(KEYINPUT55), .B(n984), .Z(n986) );
  INV_X1 U1081 ( .A(G29), .ZN(n985) );
  NAND2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1083 ( .A1(G11), .A2(n987), .ZN(n1015) );
  XOR2_X1 U1084 ( .A(G16), .B(KEYINPUT56), .Z(n1012) );
  XNOR2_X1 U1085 ( .A(G1966), .B(G168), .ZN(n989) );
  NAND2_X1 U1086 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1087 ( .A(n990), .B(KEYINPUT122), .ZN(n991) );
  XNOR2_X1 U1088 ( .A(KEYINPUT57), .B(n991), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(G1348), .B(n992), .Z(n996) );
  XNOR2_X1 U1090 ( .A(G1956), .B(G299), .ZN(n993) );
  NOR2_X1 U1091 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1092 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(n997), .B(G1341), .ZN(n998) );
  NOR2_X1 U1094 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1010) );
  XOR2_X1 U1096 ( .A(G301), .B(G1961), .Z(n1002) );
  XNOR2_X1 U1097 ( .A(n1002), .B(KEYINPUT123), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(G1971), .A2(G303), .ZN(n1003) );
  NAND2_X1 U1099 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1100 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1104 ( .A(n1013), .B(KEYINPUT124), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(n1020), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1109 ( .A(G150), .ZN(G311) );
endmodule

