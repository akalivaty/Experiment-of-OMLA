//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT14), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  AND3_X1   g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT84), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G50gat), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(G43gat), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT15), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(G50gat), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT15), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n208), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n208), .A2(new_n218), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n223), .A2(G1gat), .ZN(new_n228));
  OAI21_X1  g027(.A(G8gat), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n226), .B(new_n230), .C1(G1gat), .C2(new_n223), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n219), .A2(new_n233), .A3(new_n220), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n222), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT85), .ZN(new_n236));
  INV_X1    g035(.A(new_n221), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n229), .A2(new_n231), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT85), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n222), .A2(new_n241), .A3(new_n232), .A4(new_n234), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n236), .A2(new_n239), .A3(new_n240), .A4(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT18), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n232), .A2(new_n221), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n240), .B(KEYINPUT13), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT83), .ZN(new_n252));
  XOR2_X1   g051(.A(G169gat), .B(G197gat), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n254), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT12), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n254), .B(new_n255), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT12), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n250), .A2(new_n263), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n219), .A2(new_n233), .A3(new_n220), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n233), .B1(new_n219), .B2(new_n220), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n241), .B1(new_n267), .B2(new_n232), .ZN(new_n268));
  INV_X1    g067(.A(new_n242), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n270), .A2(KEYINPUT18), .A3(new_n239), .A4(new_n240), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT18), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n243), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n271), .A2(new_n249), .A3(new_n273), .A4(new_n262), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n274), .A2(KEYINPUT86), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(KEYINPUT86), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n264), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT87), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT86), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n244), .A2(new_n279), .A3(new_n249), .A4(new_n262), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(KEYINPUT86), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n280), .A2(new_n281), .B1(new_n250), .B2(new_n263), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT87), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT96), .ZN(new_n286));
  NAND2_X1  g085(.A1(G99gat), .A2(G106gat), .ZN(new_n287));
  INV_X1    g086(.A(G85gat), .ZN(new_n288));
  INV_X1    g087(.A(G92gat), .ZN(new_n289));
  AOI22_X1  g088(.A1(KEYINPUT8), .A2(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT7), .ZN(new_n291));
  OAI211_X1 g090(.A(G85gat), .B(G92gat), .C1(new_n291), .C2(KEYINPUT91), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT92), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(KEYINPUT7), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n291), .A2(KEYINPUT91), .A3(KEYINPUT92), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n290), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G99gat), .B(G106gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n301), .B(new_n290), .C1(new_n298), .C2(new_n299), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(KEYINPUT93), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n300), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT93), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n307), .A3(new_n301), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n305), .A2(new_n222), .A3(new_n308), .A4(new_n234), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT94), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT94), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n267), .A2(new_n311), .A3(new_n308), .A4(new_n305), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n303), .A2(KEYINPUT93), .A3(new_n304), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n300), .A2(KEYINPUT93), .A3(new_n302), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n237), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n310), .A2(new_n312), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT95), .ZN(new_n318));
  XNOR2_X1  g117(.A(G190gat), .B(G218gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n318), .B1(new_n317), .B2(new_n319), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n286), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n317), .A2(new_n319), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT95), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(KEYINPUT96), .A3(new_n320), .ZN(new_n326));
  XNOR2_X1  g125(.A(G134gat), .B(G162gat), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n317), .A2(new_n319), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n323), .A2(new_n326), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G127gat), .B(G155gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(G211gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT88), .ZN(new_n334));
  INV_X1    g133(.A(G57gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(G64gat), .ZN(new_n336));
  INV_X1    g135(.A(G64gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(KEYINPUT88), .A3(G57gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n336), .B(new_n338), .C1(G57gat), .C2(new_n337), .ZN(new_n339));
  AND2_X1   g138(.A1(G71gat), .A2(G78gat), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n340), .A2(KEYINPUT9), .ZN(new_n341));
  NOR2_X1   g140(.A1(G71gat), .A2(G78gat), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n339), .B(new_n341), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n340), .A2(new_n342), .ZN(new_n344));
  XNOR2_X1  g143(.A(G57gat), .B(G64gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n343), .A2(KEYINPUT21), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(G183gat), .B1(new_n348), .B2(new_n238), .ZN(new_n349));
  INV_X1    g148(.A(G183gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n343), .A2(KEYINPUT21), .A3(new_n347), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n232), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G231gat), .A2(G233gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n353), .B1(new_n349), .B2(new_n352), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n343), .A2(new_n347), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n355), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n349), .A2(new_n352), .ZN(new_n363));
  INV_X1    g162(.A(new_n353), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n360), .B1(new_n365), .B2(new_n354), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n333), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n361), .B1(new_n355), .B2(new_n356), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n360), .A3(new_n354), .ZN(new_n370));
  INV_X1    g169(.A(new_n333), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n367), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n368), .B1(new_n367), .B2(new_n372), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n325), .A2(new_n320), .A3(new_n330), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n329), .B(KEYINPUT90), .Z(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G230gat), .A2(G233gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n305), .A2(new_n357), .A3(new_n308), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n358), .A2(new_n303), .A3(new_n304), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT98), .ZN(new_n383));
  XNOR2_X1  g182(.A(G120gat), .B(G148gat), .ZN(new_n384));
  INV_X1    g183(.A(G204gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT99), .B(G176gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n386), .B(new_n387), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n379), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n380), .A2(new_n391), .A3(new_n381), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT10), .B(new_n358), .C1(new_n313), .C2(new_n314), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT97), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI211_X1 g195(.A(KEYINPUT97), .B(new_n390), .C1(new_n392), .C2(new_n393), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n383), .B(new_n389), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n388), .B1(new_n394), .B2(new_n382), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n331), .A2(new_n375), .A3(new_n378), .A4(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT31), .B(G50gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(G22gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT2), .ZN(new_n406));
  INV_X1    g205(.A(G148gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(G141gat), .ZN(new_n408));
  INV_X1    g207(.A(G141gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(G148gat), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n406), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G155gat), .B(G162gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT72), .B(G148gat), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n408), .B1(new_n415), .B2(G141gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(KEYINPUT73), .A2(G155gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT2), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n414), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G197gat), .B(G204gat), .ZN(new_n421));
  XOR2_X1   g220(.A(KEYINPUT69), .B(G211gat), .Z(new_n422));
  INV_X1    g221(.A(G218gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n421), .B1(new_n424), .B2(KEYINPUT22), .ZN(new_n425));
  XNOR2_X1  g224(.A(G211gat), .B(G218gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n427), .A2(KEYINPUT29), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n420), .B1(new_n428), .B2(KEYINPUT3), .ZN(new_n429));
  INV_X1    g228(.A(new_n426), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n425), .B(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n420), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT29), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT78), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT78), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n431), .B2(new_n435), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n429), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(G228gat), .A2(G233gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n420), .B1(new_n428), .B2(new_n433), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n436), .A2(new_n441), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G78gat), .B(G106gat), .ZN(new_n446));
  XOR2_X1   g245(.A(new_n446), .B(KEYINPUT77), .Z(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n442), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(new_n442), .B2(new_n445), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n405), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n442), .A2(new_n445), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n447), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n442), .A2(new_n445), .A3(new_n448), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n404), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT68), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT27), .B(G183gat), .ZN(new_n458));
  INV_X1    g257(.A(G190gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT28), .ZN(new_n461));
  INV_X1    g260(.A(G169gat), .ZN(new_n462));
  INV_X1    g261(.A(G176gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT26), .ZN(new_n465));
  OR3_X1    g264(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n465), .B(new_n466), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  NAND2_X1  g266(.A1(G183gat), .A2(G190gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT28), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n458), .A2(new_n469), .A3(new_n459), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n461), .A2(new_n467), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  XOR2_X1   g270(.A(KEYINPUT65), .B(G169gat), .Z(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(KEYINPUT23), .A3(new_n463), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT24), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(G183gat), .A2(G190gat), .ZN(new_n477));
  OR3_X1    g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT25), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT23), .B1(new_n462), .B2(new_n463), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n464), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n473), .A2(new_n478), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n471), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n475), .A2(new_n477), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n476), .A2(KEYINPUT66), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(KEYINPUT66), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT23), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n487), .B(new_n481), .C1(new_n488), .C2(new_n464), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT25), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G134gat), .ZN(new_n492));
  INV_X1    g291(.A(G120gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G113gat), .ZN(new_n494));
  INV_X1    g293(.A(G113gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G120gat), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT67), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT1), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(G127gat), .ZN(new_n500));
  AOI211_X1 g299(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n494), .C2(new_n496), .ZN(new_n501));
  INV_X1    g300(.A(G127gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n492), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(G127gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n502), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(G134gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G227gat), .A2(G233gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n510), .B(KEYINPUT64), .Z(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n483), .A2(new_n490), .A3(new_n507), .A4(new_n504), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT34), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G43gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G71gat), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n517), .B(G99gat), .Z(new_n518));
  AOI21_X1  g317(.A(new_n512), .B1(new_n509), .B2(new_n513), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(KEYINPUT33), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT32), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n520), .A2(new_n522), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n457), .B(new_n515), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n515), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n520), .A2(new_n522), .ZN(new_n528));
  INV_X1    g327(.A(new_n515), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(new_n523), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n530), .A3(KEYINPUT68), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n456), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n532), .A2(KEYINPUT35), .ZN(new_n533));
  XNOR2_X1  g332(.A(G1gat), .B(G29gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(new_n288), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT0), .B(G57gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT75), .ZN(new_n538));
  NAND2_X1  g337(.A1(G225gat), .A2(G233gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n507), .ZN(new_n540));
  AOI21_X1  g339(.A(G134gat), .B1(new_n505), .B2(new_n506), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n420), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n504), .A2(new_n432), .A3(new_n507), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT5), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n538), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n539), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n540), .A2(new_n420), .A3(new_n541), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n432), .B1(new_n504), .B2(new_n507), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(KEYINPUT4), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n420), .A2(KEYINPUT3), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n508), .B(new_n553), .C1(new_n420), .C2(new_n433), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT4), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n543), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n552), .A2(new_n554), .A3(new_n539), .A4(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n546), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT76), .B1(new_n557), .B2(KEYINPUT5), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n546), .A2(new_n551), .A3(KEYINPUT76), .A4(new_n557), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n537), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT6), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n537), .A3(new_n561), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT6), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n563), .B1(new_n566), .B2(new_n562), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT29), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n491), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G226gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT70), .ZN(new_n571));
  INV_X1    g370(.A(new_n570), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n569), .A2(new_n571), .B1(new_n491), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n427), .ZN(new_n574));
  XNOR2_X1  g373(.A(G8gat), .B(G36gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G64gat), .B(G92gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n572), .B1(new_n491), .B2(new_n568), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n571), .B1(new_n483), .B2(new_n490), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n431), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n574), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n581), .A2(KEYINPUT71), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(KEYINPUT71), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n574), .A2(new_n580), .ZN(new_n585));
  INV_X1    g384(.A(new_n577), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI211_X1 g386(.A(KEYINPUT30), .B(new_n577), .C1(new_n574), .C2(new_n580), .ZN(new_n588));
  OAI22_X1  g387(.A1(new_n582), .A2(new_n583), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n567), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n562), .A2(KEYINPUT79), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT79), .ZN(new_n594));
  AOI211_X1 g393(.A(new_n594), .B(new_n537), .C1(new_n560), .C2(new_n561), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n563), .B1(new_n596), .B2(new_n566), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n527), .A2(new_n530), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n456), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n590), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT35), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n533), .A2(new_n592), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(KEYINPUT39), .B(new_n539), .C1(new_n548), .C2(new_n549), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT39), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n537), .B(new_n603), .C1(new_n605), .C2(new_n539), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n606), .A2(KEYINPUT40), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(KEYINPUT40), .ZN(new_n608));
  OAI221_X1 g407(.A(new_n589), .B1(new_n593), .B2(new_n595), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n456), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT37), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n585), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n585), .A2(new_n611), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT38), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n563), .B(new_n615), .C1(new_n596), .C2(new_n566), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n585), .A2(KEYINPUT38), .A3(new_n577), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n573), .A2(new_n431), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT80), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n427), .B1(new_n578), .B2(new_n579), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT80), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n573), .A2(new_n621), .A3(new_n431), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT37), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT81), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT38), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(KEYINPUT81), .A3(KEYINPUT37), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n612), .A4(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n617), .B1(new_n629), .B2(new_n577), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n609), .B(new_n610), .C1(new_n616), .C2(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n598), .A2(KEYINPUT36), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n531), .A2(KEYINPUT36), .A3(new_n526), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n591), .A2(new_n456), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI211_X1 g435(.A(new_n285), .B(new_n402), .C1(new_n602), .C2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n567), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n589), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n224), .A2(new_n230), .ZN(new_n642));
  NOR2_X1   g441(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT42), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(G8gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(KEYINPUT100), .Z(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(G1325gat));
  INV_X1    g447(.A(new_n598), .ZN(new_n649));
  AOI21_X1  g448(.A(G15gat), .B1(new_n637), .B2(new_n649), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n632), .A2(KEYINPUT101), .A3(new_n633), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT101), .B1(new_n632), .B2(new_n633), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n654), .A2(G15gat), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n650), .B1(new_n637), .B2(new_n655), .ZN(G1326gat));
  NAND2_X1  g455(.A1(new_n637), .A2(new_n456), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT43), .B(G22gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  AOI21_X1  g458(.A(new_n285), .B1(new_n602), .B2(new_n636), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n331), .A2(new_n378), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n375), .A2(new_n400), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(new_n202), .A3(new_n638), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT45), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n602), .A2(new_n636), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(KEYINPUT44), .A3(new_n661), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n282), .A2(new_n375), .A3(new_n400), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n331), .A2(new_n378), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n631), .A3(new_n635), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(new_n671), .B2(new_n602), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n668), .B(new_n669), .C1(KEYINPUT44), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT102), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n602), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n661), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n678), .A2(new_n679), .A3(new_n669), .A4(new_n668), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n567), .B1(new_n674), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n666), .B1(new_n202), .B2(new_n681), .ZN(G1328gat));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n664), .A2(new_n683), .A3(new_n203), .A4(new_n589), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n660), .A2(new_n203), .A3(new_n661), .A4(new_n662), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT46), .B1(new_n685), .B2(new_n590), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n590), .B1(new_n674), .B2(new_n680), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(new_n203), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT103), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n687), .B(new_n691), .C1(new_n688), .C2(new_n203), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(G1329gat));
  OAI21_X1  g492(.A(G43gat), .B1(new_n673), .B2(new_n653), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n663), .A2(G43gat), .A3(new_n598), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n696), .A3(KEYINPUT47), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n673), .A2(KEYINPUT102), .ZN(new_n698));
  INV_X1    g497(.A(new_n680), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n654), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n695), .B1(new_n700), .B2(G43gat), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n702));
  OAI21_X1  g501(.A(new_n697), .B1(new_n701), .B2(new_n702), .ZN(G1330gat));
  NAND2_X1  g502(.A1(new_n210), .A2(new_n212), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(new_n673), .B2(new_n610), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n663), .A2(new_n610), .A3(new_n705), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n708), .A3(KEYINPUT48), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n456), .B1(new_n698), .B2(new_n699), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n707), .B1(new_n710), .B2(new_n705), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g511(.A1(new_n331), .A2(new_n375), .A3(new_n378), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n675), .A2(new_n282), .A3(new_n713), .A4(new_n400), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n567), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(new_n335), .ZN(G1332gat));
  NOR2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n716), .A2(new_n717), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(new_n589), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT49), .B(G64gat), .Z(new_n724));
  NOR3_X1   g523(.A1(new_n718), .A2(new_n590), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT106), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n724), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n722), .A2(new_n589), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n718), .A2(new_n590), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n721), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n726), .A2(new_n731), .ZN(G1333gat));
  NOR2_X1   g531(.A1(new_n598), .A2(G71gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n722), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G71gat), .B1(new_n718), .B2(new_n653), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n734), .B2(new_n735), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(G1334gat));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n456), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g540(.A1(new_n678), .A2(new_n668), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n277), .A2(new_n375), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n400), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(KEYINPUT107), .Z(new_n745));
  NOR2_X1   g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G85gat), .B1(new_n747), .B2(new_n567), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n672), .A2(new_n743), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n672), .A2(KEYINPUT51), .A3(new_n743), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n751), .A2(KEYINPUT108), .A3(new_n752), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n567), .A2(G85gat), .A3(new_n401), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n748), .A2(new_n758), .ZN(G1336gat));
  AOI21_X1  g558(.A(new_n289), .B1(new_n746), .B2(new_n589), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n590), .A2(G92gat), .A3(new_n401), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT109), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n751), .B2(new_n752), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT52), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n753), .A2(new_n761), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(KEYINPUT52), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n766), .B2(new_n760), .ZN(G1337gat));
  OAI21_X1  g566(.A(G99gat), .B1(new_n747), .B2(new_n653), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n598), .A2(new_n401), .A3(G99gat), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT110), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n756), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(G1338gat));
  INV_X1    g571(.A(G106gat), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n746), .B2(new_n456), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n456), .A2(new_n773), .A3(new_n400), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n751), .B2(new_n752), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n774), .A2(KEYINPUT53), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT53), .B1(new_n774), .B2(new_n776), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1339gat));
  INV_X1    g578(.A(new_n375), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n392), .A2(new_n393), .A3(new_n390), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT54), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n396), .B2(new_n397), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n785));
  AOI21_X1  g584(.A(new_n389), .B1(new_n394), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n786), .A3(KEYINPUT55), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n398), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n392), .A2(new_n393), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n379), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT97), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n394), .A2(new_n395), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n782), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n786), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n789), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n788), .A2(new_n277), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n247), .A2(new_n248), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n270), .A2(new_n239), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n240), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n257), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n400), .B(new_n801), .C1(new_n275), .C2(new_n276), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n661), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n280), .A2(new_n281), .B1(new_n257), .B2(new_n800), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n661), .A2(new_n804), .A3(new_n788), .A4(new_n796), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n780), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n713), .A2(new_n808), .A3(new_n282), .A4(new_n401), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT111), .B1(new_n402), .B2(new_n277), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n807), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n398), .A3(new_n787), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n802), .B1(new_n814), .B2(new_n282), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n670), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n375), .B1(new_n816), .B2(new_n805), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n809), .A2(new_n810), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT113), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n638), .A3(new_n532), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n823), .A2(new_n590), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n495), .A3(new_n277), .ZN(new_n826));
  INV_X1    g625(.A(new_n285), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n638), .A2(new_n590), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n820), .A2(new_n599), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n833), .A2(KEYINPUT115), .A3(G113gat), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT115), .B1(new_n833), .B2(G113gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n826), .B1(new_n834), .B2(new_n835), .ZN(G1340gat));
  NOR2_X1   g635(.A1(new_n401), .A2(new_n589), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n823), .A2(new_n493), .A3(new_n824), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n400), .B1(new_n831), .B2(new_n832), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n839), .A2(new_n840), .A3(G120gat), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n839), .B2(G120gat), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(G1341gat));
  OAI21_X1  g642(.A(new_n375), .B1(new_n831), .B2(new_n832), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n502), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n825), .A2(new_n375), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(new_n502), .ZN(G1342gat));
  NAND4_X1  g646(.A1(new_n823), .A2(new_n492), .A3(new_n590), .A4(new_n824), .ZN(new_n848));
  OR3_X1    g647(.A1(new_n848), .A2(KEYINPUT56), .A3(new_n670), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n661), .B1(new_n831), .B2(new_n832), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(G134gat), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT56), .B1(new_n848), .B2(new_n670), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(G1343gat));
  NOR2_X1   g652(.A1(new_n654), .A2(new_n610), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n820), .A2(new_n638), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n589), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n409), .A3(new_n827), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n653), .A2(new_n829), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n813), .A2(new_n819), .A3(new_n456), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g661(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n794), .B2(new_n795), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n278), .A2(new_n284), .A3(new_n788), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n802), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n670), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n375), .B1(new_n867), .B2(new_n805), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT57), .B(new_n456), .C1(new_n868), .C2(new_n818), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n859), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(new_n827), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n857), .B(new_n858), .C1(new_n871), .C2(new_n409), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n277), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G141gat), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(new_n857), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n872), .B1(new_n875), .B2(new_n858), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n860), .A2(KEYINPUT57), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n827), .A2(new_n402), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n861), .B(new_n456), .C1(new_n868), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(new_n401), .A3(new_n859), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT59), .B1(new_n881), .B2(new_n407), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n870), .A2(new_n400), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n415), .A2(KEYINPUT59), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n883), .A2(KEYINPUT119), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT119), .B1(new_n883), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n837), .A2(new_n415), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n855), .B2(new_n888), .ZN(G1345gat));
  NAND2_X1  g688(.A1(new_n856), .A2(new_n375), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT120), .ZN(new_n891));
  XOR2_X1   g690(.A(KEYINPUT73), .B(G155gat), .Z(new_n892));
  NOR2_X1   g691(.A1(new_n780), .A2(new_n892), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n891), .A2(new_n892), .B1(new_n870), .B2(new_n893), .ZN(G1346gat));
  AOI21_X1  g693(.A(G162gat), .B1(new_n856), .B2(new_n661), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n661), .A2(G162gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n870), .B2(new_n896), .ZN(G1347gat));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n813), .A2(new_n819), .A3(new_n567), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n813), .A2(new_n819), .A3(KEYINPUT121), .A4(new_n567), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n532), .A2(new_n589), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n898), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT122), .B(new_n904), .C1(new_n901), .C2(new_n902), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n472), .A3(new_n277), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n638), .A2(new_n590), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n813), .A2(new_n819), .A3(new_n599), .A4(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n911), .B(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(new_n827), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n909), .B1(new_n462), .B2(new_n914), .ZN(G1348gat));
  NOR2_X1   g714(.A1(new_n401), .A2(G176gat), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n906), .A2(new_n907), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n463), .B1(new_n913), .B2(new_n400), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n918), .A2(KEYINPUT124), .A3(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n903), .A2(new_n905), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT122), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n904), .B1(new_n901), .B2(new_n902), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n898), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n925), .A3(new_n916), .ZN(new_n926));
  INV_X1    g725(.A(new_n919), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n920), .A2(new_n928), .ZN(G1349gat));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n375), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(G183gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n375), .A2(new_n458), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT125), .B1(new_n924), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT60), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1350gat));
  AOI21_X1  g738(.A(new_n459), .B1(new_n913), .B2(new_n661), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n670), .A2(G190gat), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT126), .B1(new_n908), .B2(new_n943), .ZN(new_n944));
  AND4_X1   g743(.A1(KEYINPUT126), .A2(new_n923), .A3(new_n925), .A4(new_n943), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  AND2_X1   g745(.A1(new_n903), .A2(new_n854), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(new_n589), .ZN(new_n948));
  INV_X1    g747(.A(G197gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n949), .A3(new_n277), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n653), .A2(new_n910), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n880), .A2(new_n285), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n949), .B2(new_n952), .ZN(G1352gat));
  NAND4_X1  g752(.A1(new_n947), .A2(new_n385), .A3(new_n589), .A4(new_n400), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n955));
  INV_X1    g754(.A(new_n880), .ZN(new_n956));
  INV_X1    g755(.A(new_n951), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n400), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G204gat), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n955), .A2(new_n959), .A3(new_n960), .ZN(G1353gat));
  NAND3_X1  g760(.A1(new_n948), .A2(new_n422), .A3(new_n375), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n956), .A2(new_n375), .A3(new_n957), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1354gat));
  NAND4_X1  g765(.A1(new_n947), .A2(new_n423), .A3(new_n589), .A4(new_n661), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n956), .A2(new_n661), .A3(new_n957), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G218gat), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT127), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n967), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1355gat));
endmodule


