//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(new_n460), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(new_n460), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(KEYINPUT65), .A3(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n466), .B1(new_n469), .B2(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n463), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT67), .B1(new_n463), .B2(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n470), .A2(new_n471), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT66), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n464), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI221_X1 g065(.A(new_n478), .B1(new_n482), .B2(new_n483), .C1(new_n484), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n470), .B2(new_n471), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n494), .B(new_n497), .C1(new_n471), .C2(new_n470), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n470), .B2(new_n471), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(KEYINPUT68), .B(new_n500), .C1(new_n470), .C2(new_n471), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n499), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT69), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(G62), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n520), .A2(new_n521), .B1(G75), .B2(G543), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n515), .A2(new_n517), .B1(KEYINPUT5), .B2(new_n514), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(KEYINPUT70), .A3(G62), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n512), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n526), .B1(new_n522), .B2(new_n524), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT71), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT6), .B(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n530), .A2(G543), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n532), .A2(G88), .B1(G50), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n527), .A2(KEYINPUT72), .A3(new_n529), .A4(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n528), .B2(KEYINPUT71), .ZN(new_n537));
  AOI211_X1 g112(.A(new_n512), .B(new_n526), .C1(new_n522), .C2(new_n524), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n535), .A2(new_n539), .ZN(G166));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT7), .Z(new_n542));
  AND3_X1   g117(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT73), .B(G51), .ZN(new_n544));
  AOI211_X1 g119(.A(new_n542), .B(new_n543), .C1(new_n533), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n532), .A2(G89), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  AOI22_X1  g123(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n526), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n530), .A2(G543), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n531), .A2(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n550), .A2(new_n554), .ZN(G171));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n518), .A2(new_n519), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n526), .B1(new_n559), .B2(KEYINPUT74), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n560), .B1(KEYINPUT74), .B2(new_n559), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n532), .A2(G81), .B1(G43), .B2(new_n533), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  NAND3_X1  g145(.A1(new_n523), .A2(G91), .A3(new_n530), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  AND2_X1   g147(.A1(G53), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(KEYINPUT76), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n530), .A2(new_n572), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n530), .A2(new_n573), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n574), .B1(new_n577), .B2(KEYINPUT76), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n530), .A2(new_n572), .A3(new_n573), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n571), .B(new_n576), .C1(new_n578), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n523), .A2(G65), .ZN(new_n582));
  NAND2_X1  g157(.A1(G78), .A2(G543), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n526), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  AND2_X1   g162(.A1(new_n535), .A2(new_n539), .ZN(G303));
  OAI21_X1  g163(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n533), .A2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n523), .A2(G87), .A3(new_n530), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  AOI22_X1  g167(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n526), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  INV_X1    g171(.A(G48), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n531), .A2(new_n596), .B1(new_n597), .B2(new_n553), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G305));
  AOI22_X1  g175(.A1(new_n532), .A2(G85), .B1(G47), .B2(new_n533), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G60), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n557), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(G290));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NOR2_X1   g182(.A1(G301), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n532), .A2(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n557), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(G54), .B2(new_n533), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT78), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n608), .B1(new_n617), .B2(new_n607), .ZN(G284));
  AOI21_X1  g193(.A(new_n608), .B1(new_n617), .B2(new_n607), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n585), .ZN(G280));
  XOR2_X1   g196(.A(G280), .B(KEYINPUT79), .Z(G297));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g203(.A(new_n490), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G135), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT82), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(G111), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(new_n482), .ZN(new_n635));
  AND2_X1   g210(.A1(new_n635), .A2(G123), .ZN(new_n636));
  NOR3_X1   g211(.A1(new_n631), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G2096), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n463), .A2(new_n461), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT81), .B(G2100), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n640), .A3(new_n646), .ZN(G156));
  XOR2_X1   g222(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n648));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  AOI21_X1  g226(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n650), .B2(new_n651), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(G14), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT84), .Z(G401));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2096), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT85), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n677), .A2(new_n679), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n682), .A3(new_n680), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n682), .C2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT94), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G105), .B2(new_n461), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n629), .A2(G141), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n635), .A2(G129), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n704), .B2(G32), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT27), .B(G1996), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT95), .Z(new_n709));
  INV_X1    g284(.A(G2072), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n704), .A2(G33), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT25), .Z(new_n713));
  INV_X1    g288(.A(G139), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n490), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n719));
  OAI22_X1  g294(.A1(new_n717), .A2(new_n718), .B1(new_n460), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n711), .B1(new_n720), .B2(G29), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n709), .B1(new_n710), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n704), .A2(G35), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G162), .B2(new_n704), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT29), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2090), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n727), .A2(G21), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G286), .B2(G16), .ZN(new_n729));
  INV_X1    g304(.A(G1966), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT96), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n510), .A2(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n704), .A2(G27), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G2078), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n737), .B(new_n738), .C1(new_n637), .C2(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n729), .A2(new_n730), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT97), .B(G28), .Z(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n741), .B2(KEYINPUT30), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(KEYINPUT30), .B2(new_n741), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT31), .B(G11), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G2084), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n704), .B1(KEYINPUT24), .B2(G34), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(KEYINPUT24), .B2(G34), .ZN(new_n748));
  INV_X1    g323(.A(G160), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G29), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n745), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n732), .A2(new_n739), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G5), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G171), .B2(G16), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G1961), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n706), .B2(new_n707), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n727), .A2(G20), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT23), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n585), .B2(new_n727), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1956), .ZN(new_n760));
  OAI22_X1  g335(.A1(new_n750), .A2(new_n746), .B1(new_n754), .B2(G1961), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n752), .A2(new_n756), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n722), .A2(new_n726), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G4), .A2(G16), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n617), .B2(G16), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT88), .B(G1348), .Z(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n704), .A2(G26), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT28), .ZN(new_n770));
  OR2_X1    g345(.A1(G104), .A2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n771), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n772));
  INV_X1    g347(.A(G128), .ZN(new_n773));
  INV_X1    g348(.A(G140), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n772), .B1(new_n482), .B2(new_n773), .C1(new_n774), .C2(new_n490), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n770), .B1(new_n776), .B2(new_n704), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT91), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT90), .B(G2067), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n766), .A2(new_n767), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n768), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n721), .A2(new_n710), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n727), .A2(G19), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n564), .B2(new_n727), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT89), .B(G1341), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n786), .B2(new_n787), .ZN(new_n789));
  OR3_X1    g364(.A1(new_n763), .A2(new_n782), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n727), .A2(G23), .ZN(new_n791));
  INV_X1    g366(.A(G288), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n727), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT33), .B(G1976), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n727), .A2(G22), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G166), .B2(new_n727), .ZN(new_n797));
  NOR2_X1   g372(.A1(G6), .A2(G16), .ZN(new_n798));
  INV_X1    g373(.A(G305), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT32), .ZN(new_n801));
  INV_X1    g376(.A(G1981), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  OAI221_X1 g379(.A(new_n795), .B1(G1971), .B2(new_n797), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n797), .A2(G1971), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n805), .A2(KEYINPUT34), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT34), .B1(new_n805), .B2(new_n806), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT87), .B1(G95), .B2(G2105), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NOR3_X1   g385(.A1(KEYINPUT87), .A2(G95), .A3(G2105), .ZN(new_n811));
  OAI221_X1 g386(.A(G2104), .B1(G107), .B2(new_n460), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G119), .ZN(new_n813));
  INV_X1    g388(.A(G131), .ZN(new_n814));
  OAI221_X1 g389(.A(new_n812), .B1(new_n482), .B2(new_n813), .C1(new_n814), .C2(new_n490), .ZN(new_n815));
  MUX2_X1   g390(.A(G25), .B(new_n815), .S(G29), .Z(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  MUX2_X1   g394(.A(G24), .B(G290), .S(G16), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1986), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n807), .A2(new_n808), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT36), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(KEYINPUT36), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n790), .B1(new_n824), .B2(new_n825), .ZN(G311));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n824), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n763), .A2(new_n782), .A3(new_n789), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(G150));
  AOI22_X1  g404(.A1(new_n532), .A2(G93), .B1(G55), .B2(new_n533), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n526), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(new_n564), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n563), .A2(new_n833), .A3(new_n832), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n617), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT99), .ZN(new_n844));
  AOI21_X1  g419(.A(G860), .B1(new_n841), .B2(new_n842), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n832), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G145));
  AOI21_X1  g424(.A(KEYINPUT68), .B1(new_n463), .B2(new_n500), .ZN(new_n850));
  INV_X1    g425(.A(new_n504), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n509), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n498), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n497), .B1(new_n463), .B2(new_n494), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT101), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n496), .A2(new_n856), .A3(new_n498), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n852), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n775), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n720), .A2(new_n702), .ZN(new_n861));
  OR2_X1    g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n863));
  INV_X1    g438(.A(G142), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n490), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(G130), .B2(new_n635), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n720), .A2(new_n702), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n867), .B1(new_n861), .B2(new_n868), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n860), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n859), .A3(new_n869), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n815), .B(new_n643), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n872), .A2(new_n874), .A3(new_n876), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(KEYINPUT102), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(G160), .B(KEYINPUT100), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n491), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n637), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n878), .A2(KEYINPUT102), .A3(new_n883), .A4(new_n879), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g464(.A(new_n625), .B(new_n838), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n616), .A2(G299), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n585), .B1(new_n611), .B2(new_n615), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(KEYINPUT41), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n890), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(new_n894), .B2(new_n890), .ZN(new_n899));
  NOR2_X1   g474(.A1(G303), .A2(G305), .ZN(new_n900));
  XNOR2_X1  g475(.A(G290), .B(G288), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(G166), .A2(new_n799), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n903), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n901), .A2(new_n902), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n900), .B2(new_n904), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n899), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n899), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g490(.A(G868), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n832), .A2(new_n607), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(G295));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n917), .ZN(G331));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  XNOR2_X1  g495(.A(G286), .B(G171), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(new_n837), .A3(new_n836), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n836), .B2(new_n837), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n896), .B(new_n897), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n924), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n893), .A3(new_n922), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n925), .A2(new_n927), .B1(new_n906), .B2(new_n910), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(G37), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n925), .A2(new_n927), .A3(new_n906), .A4(new_n910), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n925), .A2(new_n927), .ZN(new_n933));
  OAI211_X1 g508(.A(KEYINPUT104), .B(new_n886), .C1(new_n933), .C2(new_n911), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n928), .B2(G37), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT43), .B1(new_n933), .B2(new_n911), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n920), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n929), .A2(new_n937), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n934), .A2(new_n936), .A3(new_n930), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n940), .B1(KEYINPUT43), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n939), .B1(new_n942), .B2(new_n920), .ZN(G397));
  AOI21_X1  g518(.A(new_n508), .B1(new_n503), .B2(new_n504), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n496), .A2(new_n856), .A3(new_n498), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n856), .B1(new_n496), .B2(new_n498), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT105), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n855), .A2(new_n857), .ZN(new_n951));
  AOI21_X1  g526(.A(G1384), .B1(new_n951), .B2(new_n944), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n486), .A2(G137), .B1(G101), .B2(new_n461), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT65), .B1(new_n474), .B2(G2105), .ZN(new_n958));
  AOI211_X1 g533(.A(new_n467), .B(new_n460), .C1(new_n472), .C2(new_n473), .ZN(new_n959));
  OAI211_X1 g534(.A(G40), .B(new_n957), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n775), .B(G2067), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT106), .ZN(new_n963));
  INV_X1    g538(.A(G1996), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n702), .B(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n815), .B(new_n817), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(G290), .B(G1986), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n961), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(G286), .A2(G8), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n952), .A2(KEYINPUT45), .ZN(new_n973));
  INV_X1    g548(.A(new_n960), .ZN(new_n974));
  AOI21_X1  g549(.A(G1384), .B1(new_n944), .B2(new_n499), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n730), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n947), .A2(new_n979), .A3(new_n948), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n853), .A2(new_n854), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n948), .B1(new_n852), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(KEYINPUT107), .A3(KEYINPUT50), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n975), .B2(new_n979), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n980), .A2(new_n983), .A3(new_n985), .A4(new_n974), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT112), .B(G2084), .Z(new_n987));
  OAI21_X1  g562(.A(new_n978), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n972), .B1(new_n988), .B2(G8), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT51), .B1(new_n971), .B2(KEYINPUT120), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(G8), .B(new_n990), .C1(new_n988), .C2(G286), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n988), .A2(new_n972), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT121), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n992), .A2(KEYINPUT121), .A3(new_n993), .A4(new_n994), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n1001), .A3(new_n998), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n535), .A2(new_n539), .A3(G8), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n535), .A2(new_n539), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT108), .B(G2090), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n986), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n948), .A2(KEYINPUT45), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n951), .B2(new_n944), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n510), .B2(new_n948), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n960), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(G1971), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT109), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n1016));
  OAI221_X1 g591(.A(new_n1016), .B1(new_n1013), .B2(G1971), .C1(new_n986), .C2(new_n1008), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1007), .A2(G8), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(G40), .B(G160), .C1(new_n982), .C2(KEYINPUT50), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n979), .B1(new_n947), .B2(new_n948), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1019), .A2(new_n1020), .A3(new_n1008), .ZN(new_n1021));
  OAI21_X1  g596(.A(G8), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1005), .A2(new_n1022), .A3(new_n1006), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n947), .A2(G160), .A3(G40), .A4(new_n948), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1024), .A2(G8), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n594), .A2(new_n598), .A3(G1981), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(G1981), .B1(new_n594), .B2(new_n598), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(KEYINPUT49), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT49), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1028), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n1026), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1025), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n589), .A2(new_n590), .A3(G1976), .A4(new_n591), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT110), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(G8), .A3(new_n1024), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1035), .A2(G8), .A3(new_n1024), .A4(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1033), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1033), .A2(new_n1037), .A3(KEYINPUT111), .A4(new_n1040), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1018), .A2(new_n1023), .A3(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT122), .B(G1961), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n986), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n949), .A2(new_n955), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(G2078), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1050), .A2(new_n974), .A3(new_n1052), .A4(new_n976), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1049), .A2(KEYINPUT123), .A3(new_n1053), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n947), .A2(KEYINPUT45), .A3(new_n948), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n982), .A2(new_n955), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1058), .A2(new_n736), .A3(new_n974), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1056), .A2(new_n1057), .B1(new_n1051), .B2(new_n1060), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1046), .A2(G301), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1000), .A2(new_n1002), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1956), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT56), .B(G2072), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1058), .A2(new_n974), .A3(new_n1059), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n581), .B2(new_n584), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1068), .B(new_n1070), .C1(new_n581), .C2(new_n584), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1065), .A2(new_n1067), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G1348), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n986), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G2067), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n952), .A2(new_n1078), .A3(new_n974), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n617), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1074), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1075), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n960), .B1(new_n979), .B2(new_n975), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT50), .B1(new_n858), .B2(G1384), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1956), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1066), .ZN(new_n1090));
  NOR4_X1   g665(.A1(new_n1011), .A2(new_n1012), .A3(new_n960), .A4(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1086), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(KEYINPUT61), .A3(new_n1075), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1075), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g672(.A(KEYINPUT118), .B(KEYINPUT61), .C1(new_n1092), .C2(new_n1075), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1093), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1058), .A2(new_n964), .A3(new_n974), .A4(new_n1059), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT58), .B(G1341), .Z(new_n1102));
  NAND2_X1  g677(.A1(new_n1024), .A2(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1101), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n564), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT59), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1108), .B(new_n564), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT119), .B1(new_n1099), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1075), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1096), .B1(new_n1112), .B2(new_n1082), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT118), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1095), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1093), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1111), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n617), .A2(KEYINPUT60), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n1121), .B(new_n1080), .Z(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(KEYINPUT60), .B2(new_n617), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1085), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n957), .A2(G40), .A3(new_n1052), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1126), .B(new_n1011), .C1(G2105), .C2(new_n474), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1127), .A2(new_n956), .B1(new_n1051), .B2(new_n1060), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n986), .B2(new_n1048), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1049), .A2(KEYINPUT124), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1128), .B(G301), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1061), .B2(G301), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1046), .B1(new_n1125), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1128), .B1(new_n1131), .B2(new_n1130), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1125), .B1(new_n1136), .B2(G171), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1060), .A2(new_n1051), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(G301), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT125), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1143), .B(new_n1140), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1135), .B(new_n1137), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1049), .A2(KEYINPUT123), .A3(new_n1053), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT123), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1141), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1143), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1138), .A2(KEYINPUT125), .A3(new_n1141), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1135), .B1(new_n1152), .B2(new_n1137), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n999), .B(new_n1134), .C1(new_n1146), .C2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1063), .B1(new_n1124), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1033), .A2(new_n1038), .A3(new_n792), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1027), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1025), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1018), .B2(new_n1041), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n988), .A2(G8), .A3(G168), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1161), .A2(new_n1162), .A3(new_n1041), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1018), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1015), .A2(new_n1017), .A3(G8), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1165), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1161), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1018), .A2(new_n1045), .A3(new_n1023), .A4(new_n1168), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1169), .A2(new_n1162), .ZN(new_n1170));
  OAI211_X1 g745(.A(KEYINPUT113), .B(new_n1160), .C1(new_n1167), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT113), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1166), .A2(new_n1164), .B1(new_n1169), .B2(new_n1162), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1172), .B1(new_n1173), .B2(new_n1159), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n970), .B1(new_n1155), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n961), .A2(new_n964), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT46), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n963), .A2(new_n703), .ZN(new_n1179));
  INV_X1    g754(.A(new_n961), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT127), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT47), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n815), .A2(new_n818), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n966), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n776), .A2(new_n1078), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1180), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1180), .A2(G1986), .A3(G290), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n968), .A2(new_n961), .B1(KEYINPUT48), .B2(new_n1190), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1190), .A2(KEYINPUT48), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1189), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1184), .A2(new_n1185), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1176), .A2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g770(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1197), .A2(new_n888), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n1198), .A2(new_n942), .ZN(G308));
  OR2_X1    g773(.A1(new_n1198), .A2(new_n942), .ZN(G225));
endmodule


