//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT68), .B1(new_n187), .B2(G119), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n196), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n203), .A2(KEYINPUT4), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n197), .A2(new_n200), .A3(new_n205), .A4(new_n201), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT78), .ZN(new_n207));
  OAI211_X1 g021(.A(KEYINPUT4), .B(new_n206), .C1(new_n203), .C2(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT78), .B1(new_n202), .B2(G101), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n195), .B(new_n204), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT5), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n190), .A3(G116), .ZN(new_n212));
  OAI211_X1 g026(.A(G113), .B(new_n212), .C1(new_n193), .C2(new_n211), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n193), .A2(new_n194), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n196), .A2(G107), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n199), .A2(G104), .ZN(new_n216));
  OAI21_X1  g030(.A(G101), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n213), .A2(new_n214), .A3(new_n206), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g033(.A(G110), .B(G122), .Z(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n220), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n210), .A2(new_n222), .A3(new_n218), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(KEYINPUT6), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G143), .B(G146), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT0), .A3(G128), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G128), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n226), .B(G125), .C1(new_n225), .C2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT1), .B1(new_n229), .B2(G146), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(G146), .ZN(new_n231));
  INV_X1    g045(.A(G146), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(G143), .ZN(new_n233));
  OAI211_X1 g047(.A(G128), .B(new_n230), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G125), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(G143), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n229), .A2(G146), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n236), .B(new_n237), .C1(KEYINPUT1), .C2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n234), .A2(new_n235), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n228), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G953), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G224), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n241), .B(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n222), .B1(new_n210), .B2(new_n218), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT6), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n245), .A2(KEYINPUT80), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT80), .B1(new_n245), .B2(new_n246), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n224), .B(new_n244), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(G210), .B1(G237), .B2(G902), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n220), .B(KEYINPUT8), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n213), .A2(new_n214), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n206), .A2(new_n217), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n251), .B1(new_n254), .B2(new_n218), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n243), .A2(KEYINPUT7), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n256), .A2(KEYINPUT81), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(KEYINPUT81), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(new_n241), .B2(new_n259), .ZN(new_n260));
  AOI211_X1 g074(.A(KEYINPUT81), .B(new_n256), .C1(new_n228), .C2(new_n240), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n255), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(G902), .B1(new_n262), .B2(new_n223), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n249), .A2(new_n250), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n250), .B1(new_n249), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(G214), .B1(G237), .B2(G902), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G221), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT9), .B(G234), .Z(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT77), .ZN(new_n272));
  INV_X1    g086(.A(G902), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT66), .B(G137), .ZN(new_n275));
  AND2_X1   g089(.A1(KEYINPUT11), .A2(G134), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT67), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G137), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT66), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G137), .ZN(new_n281));
  AND4_X1   g095(.A1(KEYINPUT67), .A2(new_n279), .A3(new_n281), .A4(new_n276), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT11), .ZN(new_n284));
  INV_X1    g098(.A(G134), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(G137), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n278), .A2(G134), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT65), .A3(new_n284), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n285), .A2(G137), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G131), .B1(new_n283), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n279), .A2(new_n281), .A3(new_n276), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n276), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G131), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n288), .A2(new_n290), .B1(new_n285), .B2(G137), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n234), .A2(new_n239), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n253), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n234), .A2(new_n206), .A3(new_n217), .A4(new_n239), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(KEYINPUT12), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT12), .B1(new_n303), .B2(new_n307), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT79), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n306), .B(KEYINPUT10), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n226), .B1(new_n225), .B2(new_n227), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n204), .B(new_n314), .C1(new_n208), .C2(new_n209), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n312), .A2(new_n315), .A3(new_n302), .A4(new_n294), .ZN(new_n316));
  XNOR2_X1  g130(.A(G110), .B(G140), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n242), .A2(G227), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n303), .A2(new_n307), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT12), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(new_n308), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n311), .A2(new_n321), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n312), .A2(new_n315), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n303), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n316), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n319), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G469), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(new_n273), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n316), .B1(new_n309), .B2(new_n310), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n319), .A2(new_n335), .B1(new_n321), .B2(new_n329), .ZN(new_n336));
  OAI21_X1  g150(.A(G469), .B1(new_n336), .B2(G902), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n274), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n269), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G116), .B(G122), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT85), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(new_n199), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT88), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n238), .A2(G143), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT87), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n229), .B2(G128), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n238), .A2(KEYINPUT87), .A3(G143), .ZN(new_n347));
  AOI211_X1 g161(.A(new_n343), .B(new_n344), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n347), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n229), .A2(G128), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT88), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n285), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT86), .B(KEYINPUT13), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n344), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n349), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n353), .A2(new_n344), .ZN(new_n356));
  OAI21_X1  g170(.A(G134), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n342), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n348), .A2(new_n351), .A3(new_n285), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n238), .A2(KEYINPUT87), .A3(G143), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT87), .B1(new_n238), .B2(G143), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n350), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n343), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n349), .A2(KEYINPUT88), .A3(new_n350), .ZN(new_n364));
  AOI21_X1  g178(.A(G134), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT89), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(G134), .A3(new_n364), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT89), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n352), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n187), .A2(G122), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n199), .B1(new_n371), .B2(KEYINPUT14), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(new_n340), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT90), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT90), .ZN(new_n375));
  INV_X1    g189(.A(new_n373), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n375), .B(new_n376), .C1(new_n366), .C2(new_n369), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n358), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n272), .A2(G217), .A3(new_n242), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT91), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n352), .A2(new_n367), .A3(new_n368), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n368), .B1(new_n352), .B2(new_n367), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n373), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n375), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n370), .A2(KEYINPUT90), .A3(new_n373), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n380), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n358), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n381), .A2(new_n273), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT92), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G478), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(KEYINPUT15), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n381), .A2(KEYINPUT92), .A3(new_n389), .A4(new_n273), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G140), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G125), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT74), .B1(new_n398), .B2(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n235), .A2(G140), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n400), .A3(KEYINPUT73), .ZN(new_n401));
  OR3_X1    g215(.A1(new_n397), .A2(KEYINPUT73), .A3(G125), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n399), .B1(new_n403), .B2(KEYINPUT16), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT16), .ZN(new_n405));
  AOI211_X1 g219(.A(KEYINPUT74), .B(new_n405), .C1(new_n401), .C2(new_n402), .ZN(new_n406));
  OAI21_X1  g220(.A(G146), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G237), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n242), .A3(G214), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(new_n229), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G131), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n409), .B(G143), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n300), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT17), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n399), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n397), .A2(KEYINPUT73), .A3(G125), .ZN(new_n417));
  XNOR2_X1  g231(.A(G125), .B(G140), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n417), .B1(new_n418), .B2(KEYINPUT73), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n416), .B1(new_n419), .B2(new_n405), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT74), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n403), .A2(new_n421), .A3(KEYINPUT16), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n232), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n410), .A2(KEYINPUT17), .A3(G131), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n407), .A2(new_n415), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT18), .A2(G131), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n410), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n418), .A2(new_n232), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n403), .B2(new_n232), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(G113), .B(G122), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(new_n196), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(KEYINPUT84), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n425), .A2(new_n430), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(KEYINPUT84), .B2(new_n433), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n273), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G475), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT19), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n418), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT82), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT19), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n418), .A2(new_n444), .A3(new_n440), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n407), .B(KEYINPUT83), .C1(G146), .C2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n232), .B1(new_n420), .B2(new_n422), .ZN(new_n449));
  AND4_X1   g263(.A1(new_n232), .A2(new_n442), .A3(new_n443), .A4(new_n445), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n411), .A2(new_n413), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n433), .B1(new_n427), .B2(new_n429), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n453), .A2(new_n454), .B1(new_n436), .B2(new_n433), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n456));
  NOR2_X1   g270(.A1(G475), .A2(G902), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n456), .B1(new_n455), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n439), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT93), .B(G952), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(G953), .ZN(new_n463));
  NAND2_X1  g277(.A1(G234), .A2(G237), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(G898), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(G902), .A3(G953), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n466), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n390), .A2(new_n394), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n396), .A2(new_n461), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n313), .B1(new_n294), .B2(new_n302), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n289), .B1(new_n275), .B2(G134), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n304), .B1(G131), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n479), .A2(new_n302), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n476), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n314), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n302), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(KEYINPUT30), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(new_n195), .A3(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n488));
  NAND3_X1  g302(.A1(new_n408), .A2(new_n242), .A3(G210), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT26), .B(G101), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n477), .A2(new_n480), .ZN(new_n493));
  INV_X1    g307(.A(new_n195), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n487), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT31), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n487), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n195), .B1(new_n477), .B2(new_n480), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n484), .A2(new_n494), .A3(new_n485), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT28), .B1(new_n493), .B2(new_n494), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n492), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n497), .A2(new_n499), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G472), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n273), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT32), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT32), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n506), .A2(new_n510), .A3(new_n507), .A4(new_n273), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n501), .A2(new_n502), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT28), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n502), .A2(new_n500), .ZN(new_n515));
  INV_X1    g329(.A(new_n492), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n514), .A2(KEYINPUT70), .A3(new_n515), .A4(new_n516), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n487), .A2(new_n502), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT29), .B1(new_n521), .B2(new_n492), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n503), .A2(new_n504), .A3(new_n492), .ZN(new_n524));
  AOI21_X1  g338(.A(G902), .B1(new_n524), .B2(KEYINPUT29), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G472), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n512), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT72), .B1(new_n190), .B2(G128), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT23), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n190), .A2(G128), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT23), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT72), .B(new_n532), .C1(new_n190), .C2(G128), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(G110), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT71), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n190), .B2(G128), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n238), .A2(KEYINPUT71), .A3(G119), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n537), .A2(new_n538), .A3(new_n531), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT24), .B(G110), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n407), .B(new_n428), .C1(new_n535), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT75), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n407), .A2(new_n423), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n534), .A2(G110), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n539), .A2(new_n541), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n544), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  AOI211_X1 g364(.A(KEYINPUT75), .B(new_n548), .C1(new_n407), .C2(new_n423), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n543), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT22), .B(G137), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n242), .A2(G221), .A3(G234), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n553), .B(new_n554), .Z(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n543), .B(new_n555), .C1(new_n550), .C2(new_n551), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n273), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT25), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n557), .A2(KEYINPUT25), .A3(new_n273), .A4(new_n558), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G217), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(G234), .B2(new_n273), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n557), .A2(new_n558), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(G902), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n563), .A2(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT76), .B1(new_n528), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n509), .A2(new_n511), .B1(new_n526), .B2(G472), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT76), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(new_n565), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n567), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n339), .B(new_n474), .C1(new_n569), .C2(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT94), .B(G101), .Z(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(G3));
  NAND2_X1  g392(.A1(new_n568), .A2(new_n338), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n506), .A2(new_n273), .ZN(new_n580));
  NAND2_X1  g394(.A1(KEYINPUT95), .A2(G472), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n580), .B(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT96), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n580), .B(new_n581), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n338), .A4(new_n568), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(KEYINPUT97), .Z(new_n589));
  AOI21_X1  g403(.A(new_n388), .B1(new_n387), .B2(new_n358), .ZN(new_n590));
  INV_X1    g404(.A(new_n358), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n380), .B(new_n591), .C1(new_n385), .C2(new_n386), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT33), .B1(new_n381), .B2(new_n389), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n273), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G478), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n590), .A2(new_n592), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT92), .B1(new_n598), .B2(new_n273), .ZN(new_n599));
  INV_X1    g413(.A(new_n395), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n393), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n593), .B1(new_n590), .B2(new_n592), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n381), .A2(KEYINPUT33), .A3(new_n389), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n393), .B1(new_n606), .B2(new_n273), .ZN(new_n607));
  AOI21_X1  g421(.A(G478), .B1(new_n392), .B2(new_n395), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT98), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n267), .B(new_n471), .C1(new_n264), .C2(new_n265), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n603), .A2(new_n609), .A3(new_n460), .A4(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n589), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT34), .B(G104), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  AOI211_X1 g430(.A(new_n460), .B(new_n610), .C1(new_n472), .C2(new_n396), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n589), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT99), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT35), .B(G107), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  NOR2_X1   g435(.A1(new_n556), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n552), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n567), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n572), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n474), .A2(new_n339), .A3(new_n585), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT37), .B(G110), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT100), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n626), .B(new_n628), .ZN(G12));
  AOI22_X1  g443(.A1(new_n563), .A2(new_n565), .B1(new_n567), .B2(new_n623), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n512), .B2(new_n527), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n339), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(G900), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT101), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n634), .A2(KEYINPUT101), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n469), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n465), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AOI211_X1 g453(.A(new_n460), .B(new_n639), .C1(new_n396), .C2(new_n472), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G128), .ZN(G30));
  XNOR2_X1  g456(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n638), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n338), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n492), .B1(new_n487), .B2(new_n502), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n273), .B1(new_n513), .B2(new_n516), .ZN(new_n649));
  OAI21_X1  g463(.A(G472), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n625), .B1(new_n512), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT103), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n266), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n460), .A2(new_n267), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n396), .B2(new_n472), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n647), .A2(new_n651), .A3(new_n654), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G143), .ZN(G45));
  NAND4_X1  g472(.A1(new_n603), .A2(new_n609), .A3(new_n460), .A4(new_n638), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n633), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G146), .ZN(G48));
  NAND2_X1  g476(.A1(new_n332), .A2(new_n273), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G469), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n334), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n274), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n528), .A2(new_n568), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n612), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT41), .B(G113), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G15));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n460), .B1(new_n396), .B2(new_n472), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n611), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n671), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n574), .B1(new_n512), .B2(new_n527), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n617), .A2(new_n675), .A3(KEYINPUT106), .A4(new_n666), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G116), .ZN(G18));
  NAND2_X1  g492(.A1(new_n666), .A2(new_n269), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n473), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n631), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT107), .B(G119), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G21));
  INV_X1    g497(.A(new_n266), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n684), .A2(new_n656), .A3(new_n471), .A4(new_n666), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n508), .A2(KEYINPUT108), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n580), .A2(G472), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n506), .A2(new_n688), .A3(new_n507), .A4(new_n273), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n574), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G122), .ZN(G24));
  AND2_X1   g507(.A1(new_n603), .A2(new_n609), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n694), .A2(new_n695), .A3(new_n460), .A4(new_n638), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n659), .A2(KEYINPUT110), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n687), .A2(new_n689), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n698), .A2(new_n625), .A3(new_n699), .A4(new_n686), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT109), .B1(new_n690), .B2(new_n630), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n679), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n696), .A2(new_n697), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G125), .ZN(G27));
  NAND2_X1  g518(.A1(new_n249), .A2(new_n263), .ZN(new_n705));
  INV_X1    g519(.A(new_n250), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n249), .A2(new_n250), .A3(new_n263), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n267), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT111), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n707), .A2(new_n711), .A3(new_n267), .A4(new_n708), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n710), .A2(new_n338), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n675), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n696), .A2(new_n697), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n696), .A2(KEYINPUT42), .A3(new_n697), .A4(new_n714), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G131), .ZN(G33));
  NAND3_X1  g534(.A1(new_n675), .A2(new_n640), .A3(new_n713), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  NAND2_X1  g536(.A1(new_n694), .A2(new_n461), .ZN(new_n723));
  NAND2_X1  g537(.A1(KEYINPUT112), .A2(KEYINPUT43), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n694), .A2(new_n461), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n585), .A2(new_n630), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT44), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n274), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n336), .A2(KEYINPUT45), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n336), .A2(KEYINPUT45), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(G469), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(G469), .A2(G902), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT46), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n334), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n736), .A2(new_n737), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n731), .B(new_n644), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n730), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n710), .A2(new_n712), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n728), .A2(KEYINPUT44), .A3(new_n729), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT113), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n728), .A2(new_n746), .A3(KEYINPUT44), .A4(new_n729), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n743), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n742), .B1(new_n748), .B2(KEYINPUT114), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n750));
  AOI211_X1 g564(.A(new_n750), .B(new_n743), .C1(new_n745), .C2(new_n747), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n278), .ZN(G39));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n739), .A2(new_n740), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n754), .B1(new_n755), .B2(new_n274), .ZN(new_n756));
  OAI211_X1 g570(.A(KEYINPUT47), .B(new_n731), .C1(new_n739), .C2(new_n740), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n528), .A2(new_n743), .A3(new_n568), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n660), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  NAND3_X1  g575(.A1(new_n568), .A2(new_n267), .A3(new_n731), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT115), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n665), .B(KEYINPUT49), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n512), .A2(new_n650), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n764), .A2(new_n765), .A3(new_n654), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n763), .A2(new_n766), .A3(new_n461), .A4(new_n694), .ZN(new_n767));
  INV_X1    g581(.A(new_n668), .ZN(new_n768));
  AND4_X1   g582(.A1(new_n472), .A2(new_n396), .A3(new_n461), .A4(new_n638), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n631), .A2(new_n713), .A3(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n721), .A2(new_n770), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n685), .A2(new_n691), .B1(new_n680), .B2(new_n631), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n677), .A2(new_n768), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n697), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n659), .A2(KEYINPUT110), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n700), .A2(new_n701), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n713), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n569), .A2(new_n575), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n474), .A2(new_n339), .ZN(new_n781));
  OAI22_X1  g595(.A1(new_n780), .A2(new_n781), .B1(new_n612), .B2(new_n588), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n584), .A2(new_n617), .A3(new_n587), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n783), .B1(new_n784), .B2(new_n626), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n626), .A3(new_n783), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n782), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n779), .A2(new_n719), .A3(new_n788), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n266), .B(new_n655), .C1(new_n396), .C2(new_n472), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n338), .A2(new_n638), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n651), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n703), .A2(new_n641), .A3(new_n661), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n792), .B(KEYINPUT52), .C1(new_n659), .C2(new_n632), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n703), .A2(new_n797), .A3(new_n641), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT53), .B1(new_n789), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(KEYINPUT117), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n703), .A2(new_n797), .A3(new_n802), .A4(new_n641), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n801), .A2(new_n803), .B1(new_n794), .B2(new_n793), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n779), .A2(new_n719), .A3(KEYINPUT53), .A4(new_n788), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n800), .A2(new_n806), .A3(KEYINPUT54), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n613), .A2(new_n584), .A3(new_n587), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n784), .A2(new_n626), .A3(new_n783), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n576), .B(new_n808), .C1(new_n809), .C2(new_n785), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n778), .A3(new_n773), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n799), .A2(new_n811), .A3(KEYINPUT53), .A4(new_n719), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT118), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n789), .A2(new_n814), .A3(KEYINPUT53), .A4(new_n799), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n779), .A2(new_n719), .A3(new_n788), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n816), .B1(new_n804), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n807), .B1(KEYINPUT54), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n691), .A2(new_n466), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n725), .B2(new_n727), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n654), .A2(new_n267), .A3(new_n274), .A4(new_n665), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n666), .A2(new_n710), .A3(new_n712), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT119), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n728), .A2(new_n466), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n758), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n664), .A2(new_n274), .A3(new_n334), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n743), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n776), .A2(new_n829), .B1(new_n832), .B2(new_n822), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n826), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n765), .A2(new_n574), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n828), .A2(new_n466), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT120), .ZN(new_n837));
  INV_X1    g651(.A(new_n694), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n828), .A2(new_n839), .A3(new_n466), .A4(new_n835), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n837), .A2(new_n461), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n834), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n844), .B1(new_n834), .B2(new_n843), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n838), .A2(new_n461), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n837), .A2(new_n847), .A3(new_n840), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n822), .A2(new_n269), .A3(new_n666), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n463), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n829), .A2(new_n675), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n851), .A2(KEYINPUT48), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(KEYINPUT48), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n820), .A2(new_n845), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(G952), .A2(G953), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n767), .B1(new_n856), .B2(new_n857), .ZN(G75));
  OAI211_X1 g672(.A(G210), .B(G902), .C1(new_n800), .C2(new_n806), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n859), .A2(KEYINPUT122), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(KEYINPUT122), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n224), .B1(new_n247), .B2(new_n248), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(new_n244), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT55), .Z(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n860), .A2(new_n861), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n242), .A2(G952), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n867), .B1(new_n869), .B2(new_n864), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n866), .A2(new_n870), .ZN(G51));
  XOR2_X1   g685(.A(new_n735), .B(KEYINPUT57), .Z(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n804), .A2(new_n805), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n795), .A2(new_n798), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n816), .B1(new_n875), .B2(new_n817), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n873), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n872), .B1(new_n877), .B2(new_n807), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n332), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n874), .A2(new_n876), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(G902), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n881), .A2(new_n734), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n867), .B1(new_n879), .B2(new_n882), .ZN(G54));
  INV_X1    g697(.A(new_n455), .ZN(new_n884));
  NAND2_X1  g698(.A1(KEYINPUT58), .A2(G475), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n884), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n867), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n881), .A2(new_n884), .A3(new_n885), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(G60));
  INV_X1    g704(.A(new_n606), .ZN(new_n891));
  NAND2_X1  g705(.A1(G478), .A2(G902), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT59), .Z(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n820), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n891), .A2(new_n893), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n874), .A2(new_n876), .A3(new_n873), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT54), .B1(new_n800), .B2(new_n806), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n895), .B1(new_n900), .B2(new_n867), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n896), .B1(new_n877), .B2(new_n807), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(KEYINPUT123), .A3(new_n887), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n894), .A2(new_n901), .A3(new_n903), .ZN(G63));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT60), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n880), .A2(new_n623), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n874), .B2(new_n876), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n908), .B(new_n887), .C1(new_n566), .C2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(G66));
  INV_X1    g726(.A(G224), .ZN(new_n913));
  OAI21_X1  g727(.A(G953), .B1(new_n467), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n768), .A2(new_n772), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n788), .A2(new_n677), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n914), .B1(new_n917), .B2(G953), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n862), .B1(G898), .B2(new_n242), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT125), .Z(new_n920));
  XNOR2_X1  g734(.A(new_n918), .B(new_n920), .ZN(G69));
  NAND4_X1  g735(.A1(new_n703), .A2(new_n641), .A3(new_n657), .A4(new_n661), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT62), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n569), .A2(new_n575), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n713), .A2(new_n644), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n924), .B(new_n925), .C1(new_n847), .C2(new_n672), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n923), .A2(new_n760), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n922), .A2(KEYINPUT62), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n749), .B2(new_n751), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n242), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n481), .A2(new_n486), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(new_n446), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(G900), .B2(G953), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n675), .A2(new_n790), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n741), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n760), .A2(new_n721), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n703), .A2(new_n641), .A3(new_n661), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n938), .B(new_n939), .C1(new_n717), .C2(new_n718), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n749), .B2(new_n751), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n935), .B1(new_n941), .B2(G953), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n934), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n242), .B1(G227), .B2(G900), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n944), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n934), .A2(new_n946), .A3(new_n942), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(G72));
  NAND2_X1  g762(.A1(G472), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT63), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT126), .ZN(new_n951));
  INV_X1    g765(.A(new_n917), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n930), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n648), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n521), .A2(new_n516), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n955), .A2(new_n648), .A3(new_n950), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n819), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(new_n887), .A3(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n917), .B(new_n940), .C1(new_n749), .C2(new_n751), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(KEYINPUT127), .A3(new_n951), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n955), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT127), .B1(new_n959), .B2(new_n951), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n958), .A2(new_n963), .ZN(G57));
endmodule


