//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g003(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(KEYINPUT24), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(KEYINPUT24), .B2(new_n210), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n206), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT25), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n214), .B(new_n215), .C1(new_n213), .C2(new_n212), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT25), .B1(new_n212), .B2(new_n206), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT27), .B(G183gat), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT65), .B1(new_n218), .B2(new_n208), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT28), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(new_n202), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n225), .B(new_n210), .C1(new_n224), .C2(new_n223), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n219), .A2(KEYINPUT28), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n220), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n216), .A2(new_n217), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n231));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT66), .B(G113gat), .ZN(new_n233));
  INV_X1    g032(.A(G120gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n234), .A2(G113gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n231), .B(new_n232), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G120gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n239), .A2(new_n232), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n230), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n240), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n216), .A2(new_n243), .A3(new_n229), .A4(new_n217), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n242), .A2(G227gat), .A3(G233gat), .A4(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G15gat), .B(G43gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(G71gat), .ZN(new_n247));
  INV_X1    g046(.A(G99gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT33), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n245), .A2(KEYINPUT32), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT33), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n245), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n245), .A2(KEYINPUT32), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n245), .A2(KEYINPUT67), .A3(new_n254), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n249), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n244), .ZN(new_n262));
  NAND2_X1  g061(.A1(G227gat), .A2(G233gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n266), .A2(KEYINPUT69), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G78gat), .B(G106gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT31), .B(G50gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(G22gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n272), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G228gat), .ZN(new_n276));
  INV_X1    g075(.A(G233gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n282));
  INV_X1    g081(.A(G148gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(G141gat), .ZN(new_n284));
  INV_X1    g083(.A(G141gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(G148gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n282), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G155gat), .ZN(new_n288));
  INV_X1    g087(.A(G162gat), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n281), .B(new_n287), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n279), .A2(new_n282), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(new_n288), .B2(new_n289), .ZN(new_n292));
  OR3_X1    g091(.A1(new_n285), .A2(KEYINPUT75), .A3(G148gat), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT75), .B1(new_n285), .B2(G148gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n292), .B1(new_n295), .B2(new_n284), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT3), .ZN(new_n298));
  XOR2_X1   g097(.A(KEYINPUT71), .B(KEYINPUT22), .Z(new_n299));
  XNOR2_X1  g098(.A(G197gat), .B(G204gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G211gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT72), .B(G218gat), .ZN(new_n304));
  OAI211_X1 g103(.A(G211gat), .B(new_n300), .C1(new_n299), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G218gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(KEYINPUT29), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n298), .B1(new_n309), .B2(KEYINPUT81), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n306), .B(G218gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(KEYINPUT81), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n297), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n290), .A2(new_n296), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n298), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n312), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n308), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT82), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n278), .B1(new_n315), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n309), .A2(new_n297), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n278), .A4(new_n319), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n275), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n275), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n312), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT3), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n316), .B1(new_n331), .B2(new_n313), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n319), .B(KEYINPUT82), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n325), .B(new_n328), .C1(new_n334), .C2(new_n278), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n266), .A2(KEYINPUT69), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(new_n253), .A3(new_n260), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n268), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT85), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT4), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n241), .A2(new_n316), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT4), .B1(new_n243), .B2(new_n297), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n317), .A2(new_n243), .A3(new_n324), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT5), .ZN(new_n348));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n241), .A2(new_n316), .A3(new_n351), .A4(new_n342), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n343), .A2(KEYINPUT76), .A3(new_n344), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n353), .A2(KEYINPUT77), .A3(new_n349), .A4(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n354), .A2(new_n349), .A3(new_n352), .A4(new_n346), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n243), .B(new_n297), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n362), .B2(new_n349), .ZN(new_n363));
  INV_X1    g162(.A(new_n349), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(KEYINPUT78), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n348), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n359), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n367), .B1(new_n359), .B2(new_n366), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n350), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT0), .B(G57gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(G85gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(KEYINPUT6), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT80), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(new_n375), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n374), .B(new_n350), .C1(new_n368), .C2(new_n369), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n370), .A2(new_n382), .A3(KEYINPUT6), .A4(new_n375), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n377), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT30), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n230), .A2(G226gat), .A3(G233gat), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n230), .A2(new_n312), .B1(G226gat), .B2(G233gat), .ZN(new_n387));
  OR3_X1    g186(.A1(new_n386), .A2(new_n387), .A3(new_n308), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n308), .B1(new_n386), .B2(new_n387), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(G64gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(G92gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n393), .B(KEYINPUT73), .Z(new_n394));
  AOI21_X1  g193(.A(new_n385), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(new_n390), .B2(new_n393), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n390), .A2(new_n393), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n385), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n341), .A2(new_n384), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT35), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n399), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n261), .B(new_n266), .ZN(new_n403));
  INV_X1    g202(.A(new_n336), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT35), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n401), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n268), .ZN(new_n409));
  INV_X1    g208(.A(new_n338), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT36), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n403), .B2(KEYINPUT36), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n412), .B1(new_n402), .B2(new_n404), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n347), .A2(new_n349), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT39), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n375), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n361), .A2(new_n364), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(new_n415), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n399), .B1(KEYINPUT40), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n421), .B(new_n378), .C1(KEYINPUT40), .C2(new_n420), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n390), .A2(KEYINPUT37), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n390), .A2(KEYINPUT37), .ZN(new_n426));
  AND4_X1   g225(.A1(new_n394), .A2(new_n423), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(new_n393), .A3(new_n426), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n397), .B1(new_n428), .B2(new_n424), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n377), .A2(new_n381), .A3(new_n383), .A4(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n422), .B(new_n336), .C1(new_n427), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n408), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G176gat), .B(G204gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT98), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(G120gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(new_n283), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G230gat), .A2(G233gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n439), .B(KEYINPUT97), .Z(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AND2_X1   g240(.A1(G71gat), .A2(G78gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(G71gat), .A2(G78gat), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(KEYINPUT9), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G57gat), .B(G64gat), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT92), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G71gat), .A2(G78gat), .ZN(new_n447));
  OR2_X1    g246(.A1(G71gat), .A2(G78gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT9), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G57gat), .B(G64gat), .Z(new_n451));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n446), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n447), .B(new_n448), .C1(new_n445), .C2(new_n449), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G99gat), .A2(G106gat), .ZN(new_n457));
  INV_X1    g256(.A(G85gat), .ZN(new_n458));
  INV_X1    g257(.A(G92gat), .ZN(new_n459));
  AOI22_X1  g258(.A1(KEYINPUT8), .A2(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT7), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n458), .B2(new_n459), .ZN(new_n462));
  NAND3_X1  g261(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G99gat), .B(G106gat), .Z(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n456), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT10), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n464), .A2(new_n465), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n464), .A2(new_n465), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n469), .A2(new_n454), .A3(new_n470), .A4(new_n455), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n467), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(KEYINPUT10), .A3(new_n470), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n456), .A2(KEYINPUT94), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT94), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n454), .A2(new_n475), .A3(new_n455), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n473), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n441), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n467), .A2(new_n471), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n440), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n438), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(KEYINPUT99), .ZN(new_n482));
  INV_X1    g281(.A(new_n473), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n454), .A2(new_n475), .A3(new_n455), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n475), .B1(new_n454), .B2(new_n455), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n468), .A3(new_n471), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n440), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT99), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n482), .A2(new_n480), .A3(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n491), .A2(KEYINPUT100), .A3(new_n437), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT100), .B1(new_n491), .B2(new_n437), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n481), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT95), .ZN(new_n496));
  INV_X1    g295(.A(new_n466), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n498));
  INV_X1    g297(.A(G43gat), .ZN(new_n499));
  INV_X1    g298(.A(G50gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G43gat), .A2(G50gat), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G29gat), .ZN(new_n505));
  INV_X1    g304(.A(G36gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT14), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT14), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(G29gat), .B2(G36gat), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n507), .B(new_n509), .C1(new_n505), .C2(new_n506), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT87), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n500), .ZN(new_n513));
  NAND2_X1  g312(.A1(KEYINPUT87), .A2(G50gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n499), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT86), .B(G43gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n500), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n513), .A2(KEYINPUT88), .A3(new_n499), .A4(new_n514), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n503), .B1(new_n521), .B2(new_n498), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n511), .B1(new_n522), .B2(new_n510), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n523), .A2(KEYINPUT17), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n526), .B(new_n511), .C1(new_n522), .C2(new_n510), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n529));
  AOI211_X1 g328(.A(new_n497), .B(new_n524), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT41), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n525), .A2(new_n527), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(new_n466), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n496), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G190gat), .B(G218gat), .Z(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n524), .B1(new_n528), .B2(new_n529), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n466), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n528), .A2(new_n497), .B1(KEYINPUT41), .B2(new_n531), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(KEYINPUT95), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n496), .B(new_n536), .C1(new_n530), .C2(new_n534), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT96), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n542), .A2(new_n546), .A3(new_n543), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n531), .A2(KEYINPUT41), .ZN(new_n548));
  XNOR2_X1  g347(.A(G134gat), .B(G162gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n544), .A2(KEYINPUT96), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT21), .B1(new_n484), .B2(new_n485), .ZN(new_n556));
  XNOR2_X1  g355(.A(G15gat), .B(G22gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT16), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(G1gat), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(G1gat), .B2(new_n557), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(G8gat), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n207), .ZN(new_n563));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT93), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n565), .B(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT21), .B1(new_n454), .B2(new_n455), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G211gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n569), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n568), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT18), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT90), .B1(new_n533), .B2(new_n561), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT90), .ZN(new_n576));
  INV_X1    g375(.A(new_n561), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n528), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n575), .A2(new_n578), .B1(new_n538), .B2(new_n561), .ZN(new_n579));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n574), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n528), .A2(new_n529), .ZN(new_n582));
  INV_X1    g381(.A(new_n524), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n561), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n576), .B1(new_n528), .B2(new_n577), .ZN(new_n585));
  AOI211_X1 g384(.A(KEYINPUT90), .B(new_n561), .C1(new_n525), .C2(new_n527), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n584), .B(new_n580), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(KEYINPUT18), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n528), .A2(new_n577), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n575), .A2(KEYINPUT91), .A3(new_n578), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT91), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n585), .B2(new_n586), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n589), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n580), .B(KEYINPUT13), .ZN(new_n594));
  OAI22_X1  g393(.A1(new_n581), .A2(new_n588), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT11), .B(G169gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G197gat), .ZN(new_n597));
  XOR2_X1   g396(.A(G113gat), .B(G141gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT12), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n589), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT91), .B1(new_n575), .B2(new_n578), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n585), .A2(new_n586), .A3(new_n591), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n594), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n587), .A2(KEYINPUT18), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n575), .A2(new_n578), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n610), .A2(new_n574), .A3(new_n580), .A4(new_n584), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n608), .A2(new_n612), .A3(new_n600), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n602), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n555), .A2(new_n573), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n433), .A2(new_n495), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n384), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g424(.A1(new_n621), .A2(new_n399), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT16), .B(G8gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(KEYINPUT42), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n627), .B(KEYINPUT103), .Z(new_n630));
  AND2_X1   g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n632));
  OAI21_X1  g431(.A(G8gat), .B1(new_n621), .B2(new_n399), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n633), .A2(KEYINPUT104), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(KEYINPUT104), .ZN(new_n635));
  OAI221_X1 g434(.A(new_n629), .B1(new_n631), .B2(new_n632), .C1(new_n634), .C2(new_n635), .ZN(G1325gat));
  INV_X1    g435(.A(new_n403), .ZN(new_n637));
  AOI21_X1  g436(.A(G15gat), .B1(new_n622), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n412), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n621), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n638), .B1(G15gat), .B2(new_n640), .ZN(G1326gat));
  NOR2_X1   g440(.A1(new_n621), .A2(new_n336), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT43), .B(G22gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT105), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n642), .B(new_n644), .ZN(G1327gat));
  NAND2_X1  g444(.A1(new_n433), .A2(new_n555), .ZN(new_n646));
  INV_X1    g445(.A(new_n573), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n647), .A2(new_n494), .A3(new_n615), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n505), .A3(new_n623), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT45), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n646), .A2(KEYINPUT44), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n432), .A2(KEYINPUT106), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n413), .A2(new_n431), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n408), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n555), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n649), .B1(new_n653), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(G29gat), .B1(new_n661), .B2(new_n384), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n652), .A2(new_n662), .ZN(G1328gat));
  INV_X1    g462(.A(new_n399), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n650), .A2(new_n506), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT46), .Z(new_n666));
  OAI21_X1  g465(.A(G36gat), .B1(new_n661), .B2(new_n399), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(G1329gat));
  NAND3_X1  g467(.A1(new_n660), .A2(new_n412), .A3(new_n518), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT47), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n646), .A2(new_n403), .A3(new_n649), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n669), .B(new_n671), .C1(new_n518), .C2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n670), .A2(KEYINPUT47), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(G1330gat));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n513), .A2(new_n514), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n660), .B2(new_n404), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n650), .A2(new_n404), .A3(new_n677), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n680), .B(new_n681), .Z(G1331gat));
  NOR2_X1   g481(.A1(new_n555), .A2(new_n573), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n657), .A2(new_n683), .A3(new_n615), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n494), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n623), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g487(.A1(new_n685), .A2(new_n399), .ZN(new_n689));
  NOR2_X1   g488(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n690));
  AND2_X1   g489(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n689), .B2(new_n690), .ZN(G1333gat));
  INV_X1    g492(.A(G71gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n685), .B2(new_n403), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n685), .A2(new_n694), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT110), .B1(new_n696), .B2(new_n412), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698));
  NOR4_X1   g497(.A1(new_n685), .A2(new_n698), .A3(new_n694), .A4(new_n639), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n695), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT50), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT50), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n702), .B(new_n695), .C1(new_n697), .C2(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(G1334gat));
  NAND2_X1  g503(.A1(new_n686), .A2(new_n404), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g505(.A1(new_n653), .A2(new_n659), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n647), .A2(new_n614), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n494), .A3(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n458), .A3(new_n384), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT111), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n413), .A2(new_n431), .A3(new_n655), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n655), .B1(new_n413), .B2(new_n431), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n402), .A2(new_n407), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(KEYINPUT35), .B2(new_n400), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n711), .B1(new_n716), .B2(new_n554), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n657), .A2(KEYINPUT111), .A3(new_n555), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n718), .A3(new_n708), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT51), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n708), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n657), .A2(new_n555), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(new_n711), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT51), .B1(new_n724), .B2(new_n718), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n623), .B(new_n494), .C1(new_n721), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n710), .B1(new_n726), .B2(new_n458), .ZN(G1336gat));
  NOR2_X1   g526(.A1(new_n399), .A2(G92gat), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n494), .B(new_n728), .C1(new_n721), .C2(new_n725), .ZN(new_n729));
  OAI21_X1  g528(.A(G92gat), .B1(new_n709), .B2(new_n399), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(new_n730), .B2(KEYINPUT112), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n729), .B(new_n730), .C1(KEYINPUT112), .C2(new_n732), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1337gat));
  NOR3_X1   g535(.A1(new_n709), .A2(new_n248), .A3(new_n639), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n637), .B(new_n494), .C1(new_n721), .C2(new_n725), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(new_n248), .ZN(G1338gat));
  NOR2_X1   g538(.A1(KEYINPUT113), .A2(G106gat), .ZN(new_n740));
  AOI211_X1 g539(.A(new_n495), .B(new_n722), .C1(new_n653), .C2(new_n659), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n404), .ZN(new_n742));
  NAND2_X1  g541(.A1(KEYINPUT113), .A2(G106gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n495), .A2(new_n336), .A3(G106gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n721), .B2(new_n725), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n719), .A2(new_n720), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n724), .A2(KEYINPUT51), .A3(new_n718), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n749), .A2(new_n750), .B1(new_n751), .B2(new_n745), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n745), .A2(new_n751), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n752), .A2(new_n753), .B1(new_n742), .B2(new_n743), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n748), .B1(new_n754), .B2(new_n747), .ZN(G1339gat));
  NAND2_X1  g554(.A1(new_n482), .A2(new_n490), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n438), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n486), .A2(new_n487), .A3(new_n440), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n478), .A2(KEYINPUT54), .A3(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n758), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n488), .A2(new_n489), .ZN(new_n762));
  AOI211_X1 g561(.A(KEYINPUT99), .B(new_n440), .C1(new_n486), .C2(new_n487), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(new_n437), .A3(new_n760), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n764), .A2(KEYINPUT55), .A3(new_n437), .A4(new_n760), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND4_X1   g569(.A1(new_n481), .A2(new_n761), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n608), .A2(new_n600), .A3(new_n612), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n600), .B1(new_n608), .B2(new_n612), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n589), .B(new_n607), .C1(new_n590), .C2(new_n592), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n579), .A2(new_n580), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n599), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n613), .A2(new_n777), .A3(new_n494), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n774), .A2(new_n778), .B1(new_n551), .B2(new_n553), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n771), .A2(new_n613), .A3(new_n777), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n554), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT116), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n761), .A2(new_n770), .A3(new_n481), .A4(new_n767), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n602), .B2(new_n613), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n613), .A2(new_n777), .A3(new_n494), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n554), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n613), .A2(new_n777), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n788), .A2(new_n551), .A3(new_n553), .A4(new_n771), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n782), .A2(new_n573), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n683), .A2(new_n495), .A3(new_n615), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n384), .A2(new_n664), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n405), .ZN(new_n797));
  OAI21_X1  g596(.A(G113gat), .B1(new_n797), .B2(new_n615), .ZN(new_n798));
  INV_X1    g597(.A(new_n341), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n615), .A2(new_n233), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(G1340gat));
  OAI21_X1  g602(.A(G120gat), .B1(new_n797), .B2(new_n495), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n800), .A2(new_n234), .A3(new_n494), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1341gat));
  AOI21_X1  g605(.A(G127gat), .B1(new_n800), .B2(new_n647), .ZN(new_n807));
  INV_X1    g606(.A(new_n797), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n647), .A2(G127gat), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(G1342gat));
  NOR3_X1   g609(.A1(new_n801), .A2(G134gat), .A3(new_n554), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT56), .ZN(new_n812));
  OAI21_X1  g611(.A(G134gat), .B1(new_n797), .B2(new_n554), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1343gat));
  NOR3_X1   g613(.A1(new_n412), .A2(new_n384), .A3(new_n664), .ZN(new_n815));
  XNOR2_X1  g614(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n793), .B2(new_n404), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n761), .A2(new_n770), .A3(new_n481), .ZN(new_n819));
  INV_X1    g618(.A(new_n765), .ZN(new_n820));
  XNOR2_X1  g619(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n614), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n555), .B1(new_n822), .B2(new_n778), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n573), .B1(new_n823), .B2(new_n781), .ZN(new_n824));
  AOI211_X1 g623(.A(new_n818), .B(new_n336), .C1(new_n824), .C2(new_n792), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n614), .B(new_n815), .C1(new_n817), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G141gat), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n336), .B1(new_n791), .B2(new_n792), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n828), .A2(new_n285), .A3(new_n614), .A4(new_n815), .ZN(new_n829));
  XOR2_X1   g628(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n826), .A2(new_n832), .A3(G141gat), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n826), .B2(G141gat), .ZN(new_n834));
  INV_X1    g633(.A(new_n829), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT121), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n840), .B(new_n831), .C1(new_n836), .C2(new_n837), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(G1344gat));
  NOR2_X1   g641(.A1(new_n412), .A2(new_n336), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n796), .A2(new_n283), .A3(new_n494), .A4(new_n843), .ZN(new_n844));
  XOR2_X1   g643(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n845));
  AOI21_X1  g644(.A(new_n336), .B1(new_n824), .B2(new_n792), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n847));
  OR3_X1    g646(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT57), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n846), .B2(KEYINPUT57), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n828), .A2(new_n816), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n851), .A2(new_n494), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n815), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n845), .B1(new_n853), .B2(G148gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n815), .B1(new_n817), .B2(new_n825), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n495), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(KEYINPUT59), .A3(new_n283), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n844), .B1(new_n854), .B2(new_n857), .ZN(G1345gat));
  NOR3_X1   g657(.A1(new_n855), .A2(new_n288), .A3(new_n573), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n828), .A2(new_n647), .A3(new_n815), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n288), .B2(new_n860), .ZN(G1346gat));
  NOR3_X1   g660(.A1(new_n855), .A2(new_n289), .A3(new_n554), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n828), .A2(new_n555), .A3(new_n815), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n289), .B2(new_n863), .ZN(G1347gat));
  AOI21_X1  g663(.A(new_n623), .B1(new_n791), .B2(new_n792), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n664), .A3(new_n341), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n221), .A3(new_n614), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n793), .A2(new_n384), .A3(new_n664), .A4(new_n405), .ZN(new_n869));
  OAI21_X1  g668(.A(G169gat), .B1(new_n869), .B2(new_n615), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1348gat));
  NOR3_X1   g670(.A1(new_n869), .A2(new_n222), .A3(new_n495), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n867), .A2(new_n494), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n222), .ZN(G1349gat));
  NAND3_X1  g673(.A1(new_n867), .A2(new_n218), .A3(new_n647), .ZN(new_n875));
  OAI21_X1  g674(.A(G183gat), .B1(new_n869), .B2(new_n573), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(KEYINPUT124), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n879));
  OAI221_X1 g678(.A(G190gat), .B1(KEYINPUT125), .B2(new_n879), .C1(new_n869), .C2(new_n554), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(KEYINPUT125), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n208), .A3(new_n555), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1351gat));
  NAND2_X1  g683(.A1(new_n843), .A2(new_n664), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT126), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n865), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(G197gat), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n888), .A3(new_n614), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n623), .A2(new_n412), .A3(new_n399), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n851), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(new_n614), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n889), .B1(new_n892), .B2(new_n888), .ZN(G1352gat));
  NAND2_X1  g692(.A1(new_n852), .A2(new_n890), .ZN(new_n894));
  XNOR2_X1  g693(.A(KEYINPUT127), .B(G204gat), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n495), .A2(new_n895), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n887), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT62), .Z(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(G1353gat));
  NAND3_X1  g699(.A1(new_n887), .A2(new_n302), .A3(new_n647), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n891), .A2(new_n647), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n902), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT63), .B1(new_n902), .B2(G211gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(G1354gat));
  AOI21_X1  g704(.A(G218gat), .B1(new_n887), .B2(new_n555), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n555), .A2(new_n304), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n891), .B2(new_n907), .ZN(G1355gat));
endmodule


