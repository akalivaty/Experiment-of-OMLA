//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n194));
  OR3_X1    g008(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G146), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT23), .B1(new_n197), .B2(G119), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G128), .ZN(new_n200));
  INV_X1    g014(.A(G110), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT68), .A2(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT68), .A2(G128), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .A4(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n201), .A3(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT24), .B(G110), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT68), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT68), .A2(G128), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n207), .A2(new_n208), .A3(new_n199), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT79), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n197), .B2(G119), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n199), .A2(KEYINPUT79), .A3(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n206), .B1(new_n209), .B2(new_n213), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n205), .A2(KEYINPUT81), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT81), .B1(new_n205), .B2(new_n214), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n193), .B(new_n196), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT80), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n209), .A2(new_n213), .A3(new_n206), .ZN(new_n219));
  AOI21_X1  g033(.A(G146), .B1(new_n194), .B2(new_n195), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(new_n221), .B2(new_n196), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n201), .B1(new_n200), .B2(new_n204), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n218), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n194), .A2(G146), .A3(new_n195), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(new_n220), .ZN(new_n227));
  NOR4_X1   g041(.A1(new_n227), .A2(new_n223), .A3(new_n219), .A4(KEYINPUT80), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n217), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT73), .A2(G953), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT73), .A2(G953), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(G221), .A3(G234), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT22), .B(G137), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n229), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n217), .B(new_n235), .C1(new_n225), .C2(new_n228), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n239), .B(KEYINPUT83), .ZN(new_n240));
  INV_X1    g054(.A(G234), .ZN(new_n241));
  OAI21_X1  g055(.A(G217), .B1(new_n241), .B2(G902), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(KEYINPUT84), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n237), .A2(new_n243), .A3(new_n238), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n248), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n237), .A2(new_n243), .A3(new_n238), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n242), .B(KEYINPUT78), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n246), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G237), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n232), .A2(G210), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT27), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n263));
  INV_X1    g077(.A(G113), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT70), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(KEYINPUT2), .B2(G113), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT2), .A2(G113), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OR2_X1    g084(.A1(KEYINPUT71), .A2(G116), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT71), .A2(G116), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(G119), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n199), .A2(G116), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n268), .A2(new_n273), .A3(new_n269), .A4(new_n274), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n279));
  INV_X1    g093(.A(G137), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n279), .B1(new_n280), .B2(G134), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(G134), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT66), .A3(G137), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G131), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n288));
  INV_X1    g102(.A(G143), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(G146), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n192), .A2(KEYINPUT65), .A3(G143), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(G146), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n290), .A2(new_n291), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n192), .A2(G143), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n202), .A2(new_n203), .B1(new_n295), .B2(KEYINPUT1), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n295), .A2(new_n293), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n280), .A2(G134), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT11), .B1(new_n283), .B2(G137), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT11), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n280), .A3(G134), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G131), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT67), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n285), .A2(new_n306), .A3(G131), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n287), .A2(new_n298), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n290), .A2(new_n293), .A3(new_n291), .ZN(new_n309));
  NAND2_X1  g123(.A1(KEYINPUT0), .A2(G128), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n310), .B(KEYINPUT64), .ZN(new_n313));
  NOR2_X1   g127(.A1(KEYINPUT0), .A2(G128), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(new_n295), .B2(new_n293), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI211_X1 g130(.A(G131), .B(new_n299), .C1(new_n300), .C2(new_n302), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n300), .A2(new_n302), .ZN(new_n318));
  INV_X1    g132(.A(new_n299), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n304), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n312), .B(new_n316), .C1(new_n317), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n308), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n278), .B1(new_n322), .B2(KEYINPUT74), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n285), .A2(new_n306), .A3(G131), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n306), .B1(new_n285), .B2(G131), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n295), .A2(new_n293), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n207), .A2(new_n208), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(G143), .B2(new_n192), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n327), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n331), .A2(new_n294), .B1(new_n303), .B2(new_n304), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n318), .A2(new_n319), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G131), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n305), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n309), .A2(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n326), .A2(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT28), .B1(new_n323), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n308), .A2(KEYINPUT72), .ZN(new_n342));
  INV_X1    g156(.A(new_n278), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT72), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n332), .A2(new_n344), .A3(new_n307), .A4(new_n287), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n342), .A2(new_n343), .A3(new_n321), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n322), .A2(new_n278), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n341), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n262), .B1(new_n340), .B2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n342), .A2(KEYINPUT30), .A3(new_n321), .A4(new_n345), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT69), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT30), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n351), .B1(new_n322), .B2(new_n352), .ZN(new_n353));
  AOI211_X1 g167(.A(KEYINPUT69), .B(KEYINPUT30), .C1(new_n308), .C2(new_n321), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n278), .B(new_n350), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n262), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n346), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n345), .A2(new_n321), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(KEYINPUT77), .A3(new_n343), .A4(new_n342), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n346), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n342), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n278), .B1(new_n366), .B2(new_n361), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT28), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n343), .B1(new_n337), .B2(new_n338), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n322), .A2(KEYINPUT74), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n341), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n369), .A2(KEYINPUT29), .A3(new_n372), .A4(new_n262), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n360), .A2(new_n243), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(G472), .A2(G902), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT31), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n346), .A2(new_n262), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n355), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n355), .B2(new_n378), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n356), .B1(new_n340), .B2(new_n348), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n376), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI22_X1  g197(.A1(G472), .A2(new_n374), .B1(new_n383), .B2(KEYINPUT32), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n346), .A2(new_n347), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT28), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n262), .B1(new_n386), .B2(new_n372), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n379), .A2(new_n387), .A3(new_n380), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT75), .B1(new_n388), .B2(new_n376), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n355), .A2(new_n378), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT31), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n355), .A2(new_n377), .A3(new_n378), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n382), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT75), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(new_n375), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT76), .B(KEYINPUT32), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n257), .B1(new_n384), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G214), .B1(G237), .B2(G902), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G110), .B(G122), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G104), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT3), .B1(new_n403), .B2(G107), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT3), .ZN(new_n405));
  INV_X1    g219(.A(G107), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(G104), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n403), .A2(G107), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n404), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT86), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT86), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n404), .A2(new_n407), .A3(new_n412), .A4(new_n408), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n410), .A2(new_n411), .A3(G101), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n278), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(G101), .A3(new_n413), .ZN(new_n416));
  INV_X1    g230(.A(G101), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n404), .A2(new_n407), .A3(new_n417), .A4(new_n408), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n418), .A2(KEYINPUT4), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT87), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n416), .A2(KEYINPUT87), .A3(new_n419), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n415), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n273), .A2(KEYINPUT5), .A3(new_n274), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G113), .B1(new_n274), .B2(KEYINPUT5), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n277), .ZN(new_n429));
  INV_X1    g243(.A(new_n408), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n403), .A2(G107), .ZN(new_n431));
  OAI21_X1  g245(.A(G101), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n418), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n428), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n402), .B1(new_n424), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n434), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n416), .A2(KEYINPUT87), .A3(new_n419), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT87), .B1(new_n416), .B2(new_n419), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n401), .B(new_n436), .C1(new_n439), .C2(new_n415), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n435), .A2(new_n440), .A3(KEYINPUT6), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n336), .A2(new_n189), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n298), .A2(G125), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G224), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G953), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n442), .A2(new_n443), .A3(new_n446), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n451), .B(new_n402), .C1(new_n424), .C2(new_n434), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n441), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n441), .A2(KEYINPUT91), .A3(new_n450), .A4(new_n452), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n446), .A2(KEYINPUT7), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n448), .B2(new_n449), .ZN(new_n459));
  INV_X1    g273(.A(new_n433), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n427), .B(KEYINPUT92), .Z(new_n461));
  OAI211_X1 g275(.A(new_n277), .B(new_n460), .C1(new_n461), .C2(new_n426), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n433), .B1(new_n428), .B2(new_n429), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n401), .B(KEYINPUT8), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n444), .A2(new_n458), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n459), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n440), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n243), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n457), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G210), .B1(G237), .B2(G902), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT94), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT93), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n457), .A2(new_n471), .A3(new_n475), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n400), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT9), .B(G234), .ZN(new_n480));
  OAI21_X1  g294(.A(G221), .B1(new_n480), .B2(G902), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT85), .ZN(new_n482));
  INV_X1    g296(.A(G469), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n414), .A2(new_n336), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n437), .B2(new_n438), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n290), .A2(new_n293), .A3(new_n291), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n289), .A2(G146), .ZN(new_n488));
  OAI21_X1  g302(.A(G128), .B1(new_n488), .B2(new_n329), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT88), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n487), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n294), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT10), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n460), .ZN(new_n496));
  INV_X1    g310(.A(new_n298), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT10), .B1(new_n497), .B2(new_n433), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n486), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n335), .ZN(new_n501));
  INV_X1    g315(.A(new_n335), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n486), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n232), .A2(G227), .ZN(new_n505));
  XOR2_X1   g319(.A(G110), .B(G140), .Z(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n507), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n511));
  AND4_X1   g325(.A1(new_n290), .A2(new_n291), .A3(new_n292), .A4(new_n293), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n490), .B2(KEYINPUT88), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n433), .B1(new_n513), .B2(new_n493), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n460), .A2(new_n298), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n335), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT12), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(KEYINPUT12), .B(new_n335), .C1(new_n514), .C2(new_n515), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n516), .A2(new_n511), .A3(new_n517), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n510), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n508), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n494), .A2(new_n460), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n497), .A2(new_n433), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n502), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT89), .B1(new_n528), .B2(KEYINPUT12), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n522), .A3(new_n519), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n422), .A2(new_n423), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n531), .A2(new_n485), .B1(new_n498), .B2(new_n496), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n507), .B1(new_n532), .B2(new_n502), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n530), .A2(new_n533), .A3(new_n524), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n483), .B(new_n243), .C1(new_n525), .C2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n509), .B1(new_n530), .B2(new_n503), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n510), .B1(new_n335), .B2(new_n500), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(G469), .B1(new_n538), .B2(G902), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n482), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT100), .B(G475), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT73), .ZN(new_n543));
  INV_X1    g357(.A(G953), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(KEYINPUT73), .A2(G953), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n545), .A2(G214), .A3(new_n258), .A4(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n547), .A2(new_n289), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n289), .ZN(new_n549));
  OAI21_X1  g363(.A(G131), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n547), .A2(new_n289), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n232), .A2(G143), .A3(G214), .A4(new_n258), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(KEYINPUT96), .A3(G131), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n555), .A3(new_n304), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n552), .A2(new_n553), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT96), .B1(new_n556), .B2(G131), .ZN(new_n560));
  AOI211_X1 g374(.A(new_n551), .B(new_n304), .C1(new_n554), .C2(new_n555), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT17), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n227), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(KEYINPUT18), .A2(G131), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n556), .B(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n191), .A2(KEYINPUT95), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n188), .A2(new_n190), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G146), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n193), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n563), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(G113), .B(G122), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT98), .B(G104), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n576), .B(new_n577), .Z(new_n578));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n578), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n563), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n542), .B1(new_n582), .B2(new_n243), .ZN(new_n583));
  NOR2_X1   g397(.A1(G475), .A2(G902), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT99), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n552), .A2(new_n557), .A3(new_n558), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT97), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n552), .A2(KEYINPUT97), .A3(new_n557), .A4(new_n558), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n567), .A2(KEYINPUT19), .A3(new_n570), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(KEYINPUT19), .B2(new_n568), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n196), .B1(new_n591), .B2(G146), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n580), .B1(new_n594), .B2(new_n574), .ZN(new_n595));
  INV_X1    g409(.A(new_n581), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n585), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT20), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT20), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n599), .B(new_n585), .C1(new_n595), .C2(new_n596), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n583), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G952), .ZN(new_n602));
  AOI211_X1 g416(.A(G953), .B(new_n602), .C1(G234), .C2(G237), .ZN(new_n603));
  AOI211_X1 g417(.A(new_n243), .B(new_n232), .C1(G234), .C2(G237), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT21), .B(G898), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G217), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n480), .A2(new_n608), .A3(G953), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n202), .A2(G143), .A3(new_n203), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n197), .A2(G143), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n283), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n271), .A2(G122), .A3(new_n272), .ZN(new_n616));
  INV_X1    g430(.A(G116), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n616), .B(new_n406), .C1(new_n617), .C2(G122), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n611), .A2(G134), .A3(new_n613), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n615), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n271), .A2(KEYINPUT14), .A3(G122), .A4(new_n272), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G107), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT14), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n617), .A2(G122), .ZN(new_n624));
  AND2_X1   g438(.A1(KEYINPUT71), .A2(G116), .ZN(new_n625));
  NOR2_X1   g439(.A1(KEYINPUT71), .A2(G116), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n624), .B1(new_n627), .B2(G122), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n622), .B1(new_n623), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT13), .B1(new_n328), .B2(G143), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n614), .B1(new_n631), .B2(new_n283), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n611), .A2(KEYINPUT13), .A3(G134), .A4(new_n613), .ZN(new_n633));
  INV_X1    g447(.A(G122), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n625), .A2(new_n626), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(G107), .B1(new_n635), .B2(new_n624), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n632), .A2(new_n633), .B1(new_n636), .B2(new_n618), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n610), .B1(new_n630), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n618), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT13), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n611), .A2(new_n640), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n641), .A2(G134), .B1(new_n613), .B2(new_n611), .ZN(new_n642));
  INV_X1    g456(.A(new_n633), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n644), .B(new_n609), .C1(new_n629), .C2(new_n620), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n638), .A2(KEYINPUT101), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n647), .B(new_n610), .C1(new_n630), .C2(new_n637), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(new_n243), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(G478), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(KEYINPUT15), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n649), .B(new_n651), .Z(new_n652));
  NAND3_X1  g466(.A1(new_n601), .A2(new_n607), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n398), .A2(new_n479), .A3(new_n540), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G101), .ZN(G3));
  NAND2_X1  g470(.A1(new_n472), .A2(new_n474), .ZN(new_n657));
  INV_X1    g471(.A(new_n474), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n457), .A2(new_n471), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n400), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n580), .B1(new_n563), .B2(new_n574), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n243), .B1(new_n596), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n541), .ZN(new_n663));
  INV_X1    g477(.A(new_n600), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n565), .B1(new_n193), .B2(new_n572), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n592), .B1(new_n586), .B2(new_n587), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n665), .B1(new_n666), .B2(new_n589), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n581), .B1(new_n667), .B2(new_n580), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n599), .B1(new_n668), .B2(new_n585), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n663), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT33), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n646), .A2(new_n671), .A3(new_n648), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n638), .A2(KEYINPUT33), .A3(new_n645), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n650), .A2(G902), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n649), .A2(new_n676), .A3(new_n650), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n676), .B1(new_n649), .B2(new_n650), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n670), .A2(new_n607), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n660), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n658), .B1(new_n457), .B2(new_n471), .ZN(new_n684));
  AOI211_X1 g498(.A(new_n474), .B(new_n470), .C1(new_n455), .C2(new_n456), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n399), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT103), .B1(new_n686), .B2(new_n680), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n388), .B2(G902), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n389), .A3(new_n395), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n257), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n540), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT34), .B(G104), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G6));
  INV_X1    g509(.A(new_n652), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n601), .A2(new_n607), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n686), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n540), .A3(new_n691), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT35), .B(G107), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G9));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n229), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n217), .B(new_n703), .C1(new_n225), .C2(new_n228), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n245), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT104), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n256), .A2(new_n702), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n252), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n247), .B2(new_n248), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n254), .B1(new_n711), .B2(new_n251), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n707), .B(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT105), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n653), .ZN(new_n717));
  INV_X1    g531(.A(new_n690), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(new_n479), .A3(new_n540), .A4(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT37), .B(G110), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G12));
  INV_X1    g535(.A(G900), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n603), .B1(new_n604), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n601), .A2(new_n696), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n716), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n384), .A2(new_n397), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n660), .A4(new_n540), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G128), .ZN(G30));
  AOI21_X1  g543(.A(new_n475), .B1(new_n457), .B2(new_n471), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n476), .B(new_n470), .C1(new_n455), .C2(new_n456), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT38), .Z(new_n733));
  NAND2_X1  g547(.A1(new_n256), .A2(new_n708), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n355), .A2(new_n346), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n262), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n736), .B(new_n243), .C1(new_n262), .C2(new_n368), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n383), .A2(KEYINPUT32), .B1(G472), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n734), .B1(new_n397), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n652), .A2(new_n400), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n670), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n733), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  XOR2_X1   g557(.A(new_n723), .B(KEYINPUT39), .Z(new_n744));
  NAND2_X1  g558(.A1(new_n540), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT40), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n289), .ZN(G45));
  NAND3_X1  g562(.A1(new_n670), .A2(new_n679), .A3(new_n724), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n716), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n727), .A3(new_n660), .A4(new_n540), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G146), .ZN(G48));
  AOI21_X1  g566(.A(new_n524), .B1(new_n530), .B2(new_n533), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n509), .B1(new_n501), .B2(new_n503), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n534), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(G469), .B1(new_n755), .B2(G902), .ZN(new_n756));
  INV_X1    g570(.A(new_n482), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n535), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT106), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n756), .A2(new_n760), .A3(new_n757), .A4(new_n535), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n398), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT107), .B1(new_n688), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n762), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n683), .A2(new_n687), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT41), .B(G113), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G15));
  NAND4_X1  g584(.A1(new_n698), .A2(new_n398), .A3(new_n759), .A4(new_n761), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G116), .ZN(G18));
  NAND3_X1  g586(.A1(new_n759), .A2(new_n660), .A3(new_n761), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n717), .A2(new_n727), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n199), .ZN(G21));
  AOI21_X1  g590(.A(new_n741), .B1(new_n659), .B2(new_n657), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n262), .B1(new_n369), .B2(new_n372), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n391), .A2(new_n392), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n375), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n689), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n606), .A3(new_n257), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n759), .A2(new_n777), .A3(new_n782), .A4(new_n761), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G122), .ZN(G24));
  NAND3_X1  g598(.A1(new_n734), .A2(new_n689), .A3(new_n780), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n749), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n759), .A2(new_n786), .A3(new_n660), .A4(new_n761), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G125), .ZN(G27));
  NOR2_X1   g602(.A1(new_n482), .A2(new_n400), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n477), .A2(new_n478), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT108), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n535), .A2(new_n791), .A3(new_n539), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n791), .B1(new_n535), .B2(new_n539), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n795));
  INV_X1    g609(.A(G472), .ZN(new_n796));
  AOI21_X1  g610(.A(G902), .B1(new_n358), .B2(new_n359), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n796), .B1(new_n797), .B2(new_n373), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n393), .A2(KEYINPUT32), .A3(new_n375), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT32), .B1(new_n393), .B2(new_n375), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n670), .A2(KEYINPUT42), .A3(new_n679), .A4(new_n724), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n801), .A2(new_n257), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n794), .A2(new_n795), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n789), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n730), .A2(new_n731), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n535), .A2(new_n539), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT108), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n535), .A2(new_n539), .A3(new_n791), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n374), .A2(G472), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n393), .A2(KEYINPUT32), .A3(new_n375), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT32), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n388), .B2(new_n376), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n679), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n601), .A2(new_n816), .A3(new_n723), .ZN(new_n817));
  INV_X1    g631(.A(new_n257), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(new_n817), .A3(KEYINPUT42), .A4(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT109), .B1(new_n810), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n792), .A2(new_n793), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n398), .A3(new_n817), .A4(new_n806), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT42), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n804), .A2(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(new_n304), .ZN(G33));
  INV_X1    g639(.A(new_n725), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n821), .A2(new_n398), .A3(new_n826), .A4(new_n806), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G134), .ZN(G36));
  OAI211_X1 g642(.A(new_n679), .B(new_n663), .C1(new_n664), .C2(new_n669), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT43), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n598), .A2(new_n600), .ZN(new_n833));
  XOR2_X1   g647(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n663), .A3(new_n679), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(KEYINPUT44), .A3(new_n690), .A4(new_n734), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n730), .A2(new_n731), .A3(new_n400), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n690), .A2(new_n734), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT44), .B1(new_n840), .B2(new_n836), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n530), .A2(new_n503), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n507), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n533), .A2(new_n501), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(KEYINPUT45), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT45), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n536), .B2(new_n537), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(G469), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(G469), .A2(G902), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(KEYINPUT46), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT110), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n850), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT46), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT110), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n849), .A2(new_n856), .A3(KEYINPUT46), .A4(new_n850), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n852), .A2(new_n855), .A3(new_n535), .A4(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n757), .A3(new_n744), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n842), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(G137), .ZN(G39));
  NAND2_X1  g676(.A1(new_n858), .A2(new_n757), .ZN(new_n863));
  XNOR2_X1  g677(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT47), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n858), .B(new_n757), .C1(KEYINPUT112), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n838), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n869), .A2(new_n727), .A3(new_n818), .A4(new_n749), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n866), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(G140), .ZN(G42));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n771), .A2(new_n783), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n775), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n768), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n822), .A2(new_n823), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n795), .B1(new_n794), .B2(new_n803), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n810), .A2(new_n819), .A3(KEYINPUT109), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n821), .A2(new_n786), .A3(new_n806), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n601), .A2(new_n652), .A3(new_n724), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n716), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n727), .A3(new_n540), .A4(new_n838), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n827), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n670), .A2(new_n679), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n601), .A2(new_n696), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n606), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n691), .A2(new_n888), .A3(new_n479), .A4(new_n540), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n655), .A2(new_n889), .A3(new_n719), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n723), .A2(new_n482), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n821), .A2(new_n739), .A3(new_n777), .A4(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n787), .A3(new_n728), .A4(new_n751), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n876), .A2(new_n880), .A3(new_n891), .A4(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n873), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n768), .A2(new_n880), .A3(new_n875), .A4(new_n891), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n894), .B(KEYINPUT52), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(KEYINPUT115), .A3(KEYINPUT53), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n902), .A2(KEYINPUT114), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n903), .B1(new_n902), .B2(KEYINPUT114), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT53), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT54), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n688), .A2(KEYINPUT107), .A3(new_n762), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n766), .B1(new_n764), .B2(new_n765), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n880), .B(new_n875), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT116), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n827), .A2(new_n881), .A3(new_n884), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n655), .A2(new_n719), .A3(new_n889), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT53), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n896), .B2(new_n897), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT116), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n768), .A2(new_n919), .A3(new_n880), .A4(new_n875), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n914), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT54), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n910), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n733), .A2(new_n399), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n759), .A2(new_n761), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n836), .A2(new_n603), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n930), .A2(new_n257), .A3(new_n781), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n927), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT50), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n929), .A2(new_n838), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(new_n930), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(new_n785), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n397), .A2(new_n818), .A3(new_n738), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n603), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n670), .A2(new_n679), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n866), .A2(new_n868), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n756), .A2(new_n535), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT113), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n482), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n838), .A3(new_n931), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n933), .A2(new_n941), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT51), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n935), .A2(new_n257), .A3(new_n801), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT48), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n934), .A2(new_n886), .A3(new_n938), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n931), .A2(new_n660), .A3(new_n929), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(G952), .A3(new_n544), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n948), .A2(new_n949), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n950), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI22_X1  g772(.A1(new_n926), .A2(new_n958), .B1(G952), .B2(G953), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n944), .B(KEYINPUT49), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n733), .A2(new_n805), .A3(new_n829), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n937), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n962), .ZN(G75));
  NOR2_X1   g777(.A1(new_n232), .A2(G952), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n243), .B1(new_n921), .B2(new_n923), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT56), .B1(new_n966), .B2(new_n474), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n441), .A2(new_n452), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(new_n450), .ZN(new_n969));
  XOR2_X1   g783(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n965), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n967), .A2(new_n971), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n973), .A2(KEYINPUT118), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(KEYINPUT118), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G51));
  AOI211_X1 g790(.A(new_n243), .B(new_n849), .C1(new_n921), .C2(new_n923), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n850), .B(KEYINPUT57), .Z(new_n978));
  AOI21_X1  g792(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n924), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n755), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT119), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n977), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n980), .A2(KEYINPUT119), .A3(new_n981), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n964), .B1(new_n984), .B2(new_n985), .ZN(G54));
  AND3_X1   g800(.A1(new_n966), .A2(KEYINPUT58), .A3(G475), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT120), .B1(new_n987), .B2(new_n668), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n964), .B1(new_n987), .B2(new_n668), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n987), .A2(KEYINPUT120), .A3(new_n668), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(G60));
  AND2_X1   g806(.A1(new_n672), .A2(new_n673), .ZN(new_n993));
  NAND2_X1  g807(.A1(G478), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT59), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n993), .B(new_n996), .C1(new_n924), .C2(new_n979), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n965), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n926), .A2(new_n996), .ZN(new_n999));
  INV_X1    g813(.A(new_n993), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(G63));
  NAND2_X1  g815(.A1(G217), .A2(G902), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT60), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(new_n921), .B2(new_n923), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n706), .A3(new_n705), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n1005), .B(new_n965), .C1(new_n240), .C2(new_n1004), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT61), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(G66));
  OAI21_X1  g822(.A(G953), .B1(new_n605), .B2(new_n445), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n876), .A2(new_n916), .ZN(new_n1010));
  INV_X1    g824(.A(new_n232), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n968), .B1(G898), .B2(new_n232), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(G69));
  INV_X1    g828(.A(KEYINPUT124), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT44), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n832), .A2(new_n835), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n690), .A2(new_n734), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1019), .A2(new_n837), .A3(new_n838), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n777), .A2(new_n818), .A3(new_n815), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n859), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n827), .A2(new_n787), .A3(new_n728), .A4(new_n751), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n1022), .A2(new_n824), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1015), .B1(new_n1024), .B2(new_n871), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n804), .A2(new_n820), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1023), .B1(new_n877), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1021), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n860), .B1(new_n842), .B2(new_n1028), .ZN(new_n1029));
  AND4_X1   g843(.A1(new_n1015), .A2(new_n1027), .A3(new_n871), .A4(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n232), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n232), .A2(G900), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1031), .A2(KEYINPUT125), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT125), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1023), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n1029), .A2(new_n880), .A3(new_n871), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(KEYINPUT124), .ZN(new_n1038));
  NAND4_X1  g852(.A1(new_n1027), .A2(new_n1015), .A3(new_n871), .A4(new_n1029), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1011), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1035), .B1(new_n1040), .B2(new_n1032), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n1042));
  INV_X1    g856(.A(new_n591), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1034), .A2(new_n1041), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n787), .A2(new_n728), .A3(new_n751), .ZN(new_n1047));
  OAI21_X1  g861(.A(KEYINPUT62), .B1(new_n747), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n886), .A2(new_n887), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n398), .A2(new_n838), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1050), .A2(new_n745), .ZN(new_n1051));
  XNOR2_X1  g865(.A(new_n1051), .B(KEYINPUT122), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n1048), .A2(new_n861), .A3(new_n871), .A4(new_n1052), .ZN(new_n1053));
  OR3_X1    g867(.A1(new_n747), .A2(new_n1047), .A3(KEYINPUT62), .ZN(new_n1054));
  OR2_X1    g868(.A1(new_n1054), .A2(KEYINPUT121), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1054), .A2(KEYINPUT121), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g871(.A(new_n1044), .B1(new_n1057), .B2(new_n1011), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1046), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g873(.A(KEYINPUT123), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1046), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n232), .B1(G227), .B2(G900), .ZN(new_n1062));
  INV_X1    g876(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n1059), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  OAI211_X1 g878(.A(new_n1046), .B(new_n1058), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1065));
  AND2_X1   g879(.A1(new_n1064), .A2(new_n1065), .ZN(G72));
  NAND2_X1  g880(.A1(new_n1057), .A2(new_n1010), .ZN(new_n1067));
  NAND2_X1  g881(.A1(G472), .A2(G902), .ZN(new_n1068));
  XOR2_X1   g882(.A(new_n1068), .B(KEYINPUT63), .Z(new_n1069));
  AOI21_X1  g883(.A(new_n736), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g884(.A1(new_n1070), .A2(new_n964), .ZN(new_n1071));
  NAND3_X1  g885(.A1(new_n736), .A2(new_n357), .A3(new_n1069), .ZN(new_n1072));
  XNOR2_X1  g886(.A(new_n1072), .B(KEYINPUT127), .ZN(new_n1073));
  OAI21_X1  g887(.A(new_n1073), .B1(new_n906), .B2(new_n909), .ZN(new_n1074));
  NAND3_X1  g888(.A1(new_n1010), .A2(new_n1039), .A3(new_n1038), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n1075), .A2(new_n1069), .ZN(new_n1076));
  XOR2_X1   g890(.A(new_n357), .B(KEYINPUT126), .Z(new_n1077));
  NAND2_X1  g891(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AND3_X1   g892(.A1(new_n1071), .A2(new_n1074), .A3(new_n1078), .ZN(G57));
endmodule


