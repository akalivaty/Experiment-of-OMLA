//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT66), .Z(G319));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(new_n463), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(KEYINPUT67), .A3(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n465), .A2(G2104), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(G2105), .B1(G101), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n470), .A2(G136), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n469), .A2(new_n465), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n482), .B(new_n484), .C1(G124), .C2(new_n485), .ZN(G162));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n466), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n470), .A2(KEYINPUT4), .A3(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n485), .B2(G126), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  OR2_X1    g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  OAI21_X1  g084(.A(G543), .B1(new_n506), .B2(new_n507), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OR3_X1    g087(.A1(new_n502), .A2(new_n503), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n503), .B1(new_n502), .B2(new_n512), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(G166));
  INV_X1    g090(.A(new_n508), .ZN(new_n516));
  INV_X1    g091(.A(new_n510), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(G89), .B1(new_n517), .B2(G51), .ZN(new_n518));
  XOR2_X1   g093(.A(KEYINPUT69), .B(KEYINPUT7), .Z(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n499), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(new_n521), .A3(new_n522), .ZN(G286));
  INV_X1    g098(.A(G286), .ZN(G168));
  AOI22_X1  g099(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(new_n501), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT6), .B(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT71), .B(G90), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n499), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(KEYINPUT70), .A2(G52), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT70), .A2(G52), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(new_n527), .A3(G543), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n529), .A2(new_n533), .A3(KEYINPUT72), .ZN(new_n534));
  AOI21_X1  g109(.A(KEYINPUT72), .B1(new_n529), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n526), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT71), .B(G90), .Z(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT70), .B(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n508), .A2(new_n539), .B1(new_n510), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n529), .A2(new_n533), .A3(KEYINPUT72), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(KEYINPUT73), .B1(new_n545), .B2(new_n526), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n538), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n501), .ZN(new_n550));
  XOR2_X1   g125(.A(KEYINPUT75), .B(G81), .Z(new_n551));
  XOR2_X1   g126(.A(KEYINPUT74), .B(G43), .Z(new_n552));
  OAI22_X1  g127(.A1(new_n508), .A2(new_n551), .B1(new_n552), .B2(new_n510), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n497), .A2(new_n561), .A3(new_n498), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT78), .B1(new_n505), .B2(new_n504), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT77), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT79), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n569), .B(G651), .C1(new_n564), .C2(new_n566), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n516), .A2(G91), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n527), .A2(KEYINPUT76), .A3(G53), .A4(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n568), .A2(new_n570), .A3(new_n571), .A4(new_n573), .ZN(G299));
  INV_X1    g149(.A(G166), .ZN(G303));
  AND2_X1   g150(.A1(new_n516), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n577));
  INV_X1    g152(.A(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n510), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G288));
  AOI22_X1  g156(.A1(new_n499), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n501), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  INV_X1    g159(.A(G48), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n508), .A2(new_n584), .B1(new_n510), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n583), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n516), .A2(G85), .B1(new_n517), .B2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n501), .B2(new_n589), .ZN(G290));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n508), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT10), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n562), .B2(new_n563), .ZN(new_n595));
  AND2_X1   g170(.A1(G79), .A2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n517), .A2(G54), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g176(.A(new_n600), .B1(G171), .B2(G868), .ZN(G321));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G299), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n603), .B2(G168), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(new_n603), .B2(G168), .ZN(G280));
  INV_X1    g181(.A(new_n599), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n464), .A2(new_n476), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(G2100), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n470), .A2(G135), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n485), .A2(G123), .ZN(new_n621));
  OR2_X1    g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n622), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n618), .A2(new_n619), .A3(new_n625), .ZN(G156));
  XOR2_X1   g201(.A(G2451), .B(G2454), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT82), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n628), .B(new_n630), .Z(new_n631));
  XOR2_X1   g206(.A(KEYINPUT80), .B(KEYINPUT14), .Z(new_n632));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT81), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2427), .B(G2430), .Z(new_n636));
  AOI21_X1  g211(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n631), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(G14), .A3(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n645), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n650), .B1(new_n653), .B2(new_n647), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT18), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n647), .A3(new_n645), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2096), .B(G2100), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT84), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n663), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n663), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(new_n673), .Z(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT85), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n674), .A2(new_n676), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n674), .A2(new_n676), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(G229));
  XNOR2_X1  g259(.A(KEYINPUT94), .B(KEYINPUT25), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G139), .B2(new_n470), .ZN(new_n688));
  AOI22_X1  g263(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n465), .B2(new_n689), .ZN(new_n690));
  MUX2_X1   g265(.A(G33), .B(new_n690), .S(G29), .Z(new_n691));
  NOR2_X1   g266(.A1(new_n691), .A2(G2072), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G21), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G168), .B2(new_n693), .ZN(new_n695));
  INV_X1    g270(.A(G1966), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G2078), .ZN(new_n698));
  NAND2_X1  g273(.A1(G164), .A2(G29), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G27), .B2(G29), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n697), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n691), .A2(G2072), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT97), .B(KEYINPUT31), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G11), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT98), .B(G28), .ZN(new_n705));
  AOI21_X1  g280(.A(G29), .B1(new_n705), .B2(KEYINPUT30), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(KEYINPUT30), .B2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n704), .B(new_n707), .C1(new_n624), .C2(new_n708), .ZN(new_n709));
  OR4_X1    g284(.A1(new_n692), .A2(new_n701), .A3(new_n702), .A4(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G5), .A2(G16), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G171), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1961), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n708), .A2(G32), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n470), .A2(G141), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT96), .Z(new_n716));
  AND2_X1   g291(.A1(new_n476), .A2(G105), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT26), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n717), .B(new_n719), .C1(G129), .C2(new_n485), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n714), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT27), .B(G1996), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n698), .B2(new_n700), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n722), .B2(new_n723), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(G34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n478), .B2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT95), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2084), .ZN(new_n733));
  NOR4_X1   g308(.A1(new_n710), .A2(new_n713), .A3(new_n726), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(KEYINPUT99), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n693), .A2(G20), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT23), .Z(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G299), .B2(G16), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1956), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n607), .A2(new_n693), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G4), .B2(new_n693), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT91), .B(G1348), .Z(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n693), .A2(G19), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n554), .B2(new_n693), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1341), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n708), .A2(G35), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G162), .B2(new_n708), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT29), .Z(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n746), .B1(new_n750), .B2(G2090), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n708), .A2(G26), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT28), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n485), .A2(G128), .ZN(new_n754));
  INV_X1    g329(.A(G140), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(new_n466), .ZN(new_n756));
  OAI21_X1  g331(.A(KEYINPUT92), .B1(G104), .B2(G2105), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g333(.A1(KEYINPUT92), .A2(G104), .A3(G2105), .ZN(new_n759));
  OAI221_X1 g334(.A(G2104), .B1(G116), .B2(new_n465), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n753), .B1(new_n763), .B2(new_n708), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT93), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G2090), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n749), .A2(new_n768), .B1(new_n741), .B2(new_n742), .ZN(new_n769));
  AND4_X1   g344(.A1(new_n743), .A2(new_n751), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n735), .A2(new_n739), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n693), .A2(G22), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G166), .B2(new_n693), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n773), .A2(G1971), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n693), .A2(G23), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n580), .B2(new_n693), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT33), .B(G1976), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n776), .B(new_n777), .Z(new_n778));
  NOR2_X1   g353(.A1(new_n773), .A2(G1971), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n693), .A2(G6), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n583), .A2(new_n586), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n693), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT32), .B(G1981), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT89), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n782), .B(new_n784), .Z(new_n785));
  NOR4_X1   g360(.A1(new_n774), .A2(new_n778), .A3(new_n779), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  MUX2_X1   g364(.A(G24), .B(G290), .S(G16), .Z(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1986), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n708), .A2(G25), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT86), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n485), .A2(G119), .ZN(new_n794));
  INV_X1    g369(.A(G131), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n466), .ZN(new_n796));
  OAI21_X1  g371(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n797));
  INV_X1    g372(.A(G107), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(G2105), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT87), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n793), .B1(new_n802), .B2(G29), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  XOR2_X1   g379(.A(new_n803), .B(new_n804), .Z(new_n805));
  NAND4_X1  g380(.A1(new_n788), .A2(new_n789), .A3(new_n791), .A4(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT90), .B(KEYINPUT36), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n734), .A2(KEYINPUT99), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n771), .A2(new_n808), .A3(new_n809), .ZN(G311));
  OR3_X1    g385(.A1(new_n771), .A2(new_n808), .A3(new_n809), .ZN(G150));
  INV_X1    g386(.A(G67), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n497), .B2(new_n498), .ZN(new_n813));
  NAND2_X1  g388(.A1(G80), .A2(G543), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(G651), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT102), .B(G93), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n516), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n517), .A2(G55), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n816), .A2(new_n817), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(G860), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n599), .A2(new_n608), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n820), .A2(new_n821), .ZN(new_n831));
  INV_X1    g406(.A(new_n823), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n554), .A2(new_n831), .A3(new_n832), .A4(new_n818), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n552), .A2(new_n510), .ZN(new_n834));
  OAI221_X1 g409(.A(new_n834), .B1(new_n508), .B2(new_n551), .C1(new_n501), .C2(new_n549), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n822), .B2(new_n823), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n830), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n825), .B1(new_n839), .B2(KEYINPUT39), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n827), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT103), .Z(G145));
  XOR2_X1   g418(.A(KEYINPUT105), .B(G37), .Z(new_n844));
  INV_X1    g419(.A(KEYINPUT104), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n495), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n489), .A2(KEYINPUT104), .A3(new_n494), .A4(new_n490), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n762), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n485), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n465), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G142), .B2(new_n470), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n849), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n721), .B(new_n690), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n801), .B(new_n615), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(G162), .B(new_n624), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n478), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n855), .A2(new_n858), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n859), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n862), .B1(new_n859), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n844), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g442(.A1(new_n833), .A2(new_n836), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n610), .B(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(G299), .A2(new_n599), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n872));
  NAND2_X1  g447(.A1(G299), .A2(new_n599), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n873), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT41), .B1(new_n875), .B2(new_n870), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT107), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n875), .A2(new_n870), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(KEYINPUT107), .A3(new_n872), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n869), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n879), .B(KEYINPUT106), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n869), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(G290), .B(new_n781), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(G166), .A2(new_n580), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(G166), .A2(new_n580), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n890), .A2(new_n886), .A3(new_n884), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n883), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n883), .A2(new_n894), .ZN(new_n897));
  OAI21_X1  g472(.A(G868), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n824), .A2(G868), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(G331));
  NAND2_X1  g476(.A1(G331), .A2(KEYINPUT108), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(G295));
  NAND2_X1  g480(.A1(new_n536), .A2(new_n537), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n545), .A2(KEYINPUT73), .A3(new_n526), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n906), .A2(G286), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(G286), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n868), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT110), .ZN(new_n911));
  OAI21_X1  g486(.A(G168), .B1(new_n538), .B2(new_n546), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(new_n907), .A3(G286), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n837), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  OAI211_X1 g490(.A(KEYINPUT110), .B(new_n868), .C1(new_n908), .C2(new_n909), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n879), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n910), .A2(KEYINPUT109), .A3(new_n914), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n920), .B(new_n868), .C1(new_n908), .C2(new_n909), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n878), .A2(new_n919), .A3(new_n880), .A4(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n892), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n918), .A2(new_n922), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT111), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n889), .B2(new_n891), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n884), .B1(new_n890), .B2(new_n886), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n887), .A2(new_n888), .A3(new_n885), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT111), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n925), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n924), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n931), .B1(new_n922), .B2(new_n918), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT112), .B1(new_n936), .B2(G37), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT43), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n882), .B1(new_n921), .B2(new_n919), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n917), .B1(new_n874), .B2(new_n876), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n932), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AND4_X1   g516(.A1(KEYINPUT43), .A2(new_n941), .A3(new_n844), .A4(new_n923), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT44), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n935), .B2(new_n937), .ZN(new_n946));
  AND4_X1   g521(.A1(new_n945), .A2(new_n941), .A3(new_n844), .A4(new_n923), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n948), .ZN(G397));
  NAND3_X1  g524(.A1(new_n513), .A2(G8), .A3(new_n514), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n472), .A2(G40), .A3(new_n477), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n953));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n495), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n952), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n846), .A2(KEYINPUT45), .A3(new_n954), .A4(new_n847), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1971), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n956), .A2(KEYINPUT113), .A3(new_n957), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n955), .A2(KEYINPUT50), .ZN(new_n964));
  INV_X1    g539(.A(new_n952), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n495), .A2(new_n966), .A3(new_n954), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n768), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n963), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n951), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n952), .A2(new_n955), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G8), .ZN(new_n976));
  NAND2_X1  g551(.A1(G305), .A2(G1981), .ZN(new_n977));
  OR3_X1    g552(.A1(new_n583), .A2(G1981), .A3(new_n586), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n977), .A2(KEYINPUT117), .A3(KEYINPUT49), .A4(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n978), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n976), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n981), .A2(KEYINPUT115), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT49), .B1(new_n981), .B2(KEYINPUT115), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT116), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT116), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1976), .ZN(new_n990));
  NOR2_X1   g565(.A1(G288), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n992));
  OAI22_X1  g567(.A1(new_n976), .A2(new_n991), .B1(KEYINPUT114), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n580), .A2(G1976), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(KEYINPUT114), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n975), .A2(G8), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(G288), .A2(new_n992), .A3(new_n990), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n989), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n972), .B1(new_n963), .B2(new_n970), .ZN(new_n1000));
  INV_X1    g575(.A(new_n951), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G2084), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n954), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n956), .A2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n969), .A2(new_n1003), .B1(new_n1005), .B2(new_n696), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1006), .A2(new_n972), .A3(G286), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n973), .A2(new_n999), .A3(new_n1002), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT63), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n989), .A2(new_n998), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n972), .B(new_n951), .C1(new_n963), .C2(new_n970), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(KEYINPUT63), .A3(new_n973), .A4(new_n1007), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT123), .ZN(new_n1016));
  AOI21_X1  g591(.A(G2078), .B1(new_n960), .B2(new_n962), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n962), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT113), .B1(new_n956), .B2(new_n957), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n698), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1018), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(KEYINPUT123), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n955), .A2(new_n953), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1026), .A2(new_n965), .A3(new_n1004), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n698), .A2(KEYINPUT53), .ZN(new_n1028));
  INV_X1    g603(.A(G1961), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1027), .A2(new_n1028), .B1(new_n968), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(G301), .B(KEYINPUT54), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n1034));
  OAI21_X1  g609(.A(G299), .B1(KEYINPUT118), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(KEYINPUT118), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1035), .B(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1956), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n968), .A2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT56), .B(G2072), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n956), .A2(new_n957), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n968), .A2(new_n742), .B1(new_n766), .B2(new_n974), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(new_n599), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1046), .A2(new_n1045), .A3(new_n599), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1048), .A2(new_n1049), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT120), .B(G1996), .Z(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT58), .B(G1341), .ZN(new_n1052));
  OAI22_X1  g627(.A1(new_n958), .A2(new_n1051), .B1(new_n974), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n554), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(KEYINPUT59), .A3(new_n554), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1046), .A2(new_n607), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1056), .B(new_n1057), .C1(KEYINPUT60), .C2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT61), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1035), .B(new_n1036), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT61), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1058), .A2(KEYINPUT60), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1046), .A2(new_n607), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1060), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1050), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT45), .B1(new_n848), .B2(new_n954), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n957), .A2(new_n965), .A3(new_n1028), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1068), .A2(new_n1069), .B1(new_n969), .B2(G1961), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(new_n1032), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G286), .A2(G8), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n1072), .B2(KEYINPUT121), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1072), .B(new_n1075), .C1(new_n1006), .C2(new_n972), .ZN(new_n1076));
  OAI22_X1  g651(.A1(new_n1027), .A2(G1966), .B1(new_n968), .B2(G2084), .ZN(new_n1077));
  OAI211_X1 g652(.A(G8), .B(new_n1074), .C1(new_n1077), .C2(G286), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(G8), .A3(G286), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1025), .A2(new_n1071), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1082), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1033), .A2(new_n1067), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(G301), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1079), .A2(KEYINPUT62), .A3(new_n1080), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT62), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1083), .B(new_n1085), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n989), .A2(new_n990), .A3(new_n580), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n976), .B1(new_n1089), .B2(new_n978), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n999), .B2(new_n1012), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1015), .A2(new_n1084), .A3(new_n1088), .A4(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1068), .A2(new_n965), .ZN(new_n1093));
  INV_X1    g668(.A(G1996), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n721), .B(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n762), .B(new_n766), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n801), .A2(new_n804), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n801), .A2(new_n804), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(G290), .B(G1986), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1093), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1092), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1097), .B(KEYINPUT124), .ZN(new_n1104));
  OAI22_X1  g679(.A1(new_n1103), .A2(new_n1104), .B1(G2067), .B2(new_n762), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n1093), .ZN(new_n1106));
  XOR2_X1   g681(.A(new_n1106), .B(KEYINPUT125), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1099), .A2(new_n1093), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT126), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G290), .A2(G1986), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1093), .A2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(new_n1111), .B(KEYINPUT48), .Z(new_n1112));
  OAI21_X1  g687(.A(new_n1107), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1114), .A2(KEYINPUT46), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(KEYINPUT46), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1096), .A2(new_n716), .A3(new_n720), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1115), .A2(new_n1116), .B1(new_n1093), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1118), .A2(KEYINPUT47), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(KEYINPUT47), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1113), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1102), .A2(new_n1121), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g697(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1124));
  NAND3_X1  g698(.A1(new_n680), .A2(new_n1124), .A3(new_n683), .ZN(new_n1125));
  NAND2_X1  g699(.A1(new_n1125), .A2(KEYINPUT127), .ZN(new_n1126));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n1127));
  NAND4_X1  g701(.A1(new_n680), .A2(new_n1124), .A3(new_n1127), .A4(new_n683), .ZN(new_n1128));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g703(.A(new_n866), .B(new_n1129), .C1(new_n946), .C2(new_n947), .ZN(G225));
  INV_X1    g704(.A(G225), .ZN(G308));
endmodule


