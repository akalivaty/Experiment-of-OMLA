

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735;

  XNOR2_X1 U372 ( .A(n535), .B(n534), .ZN(n544) );
  XNOR2_X1 U373 ( .A(n540), .B(KEYINPUT32), .ZN(n612) );
  NOR2_X1 U374 ( .A1(n602), .A2(n639), .ZN(n604) );
  OR2_X2 U375 ( .A1(n561), .A2(n566), .ZN(n681) );
  XNOR2_X2 U376 ( .A(n452), .B(n360), .ZN(n722) );
  XNOR2_X2 U377 ( .A(n414), .B(G134), .ZN(n452) );
  XNOR2_X2 U378 ( .A(n722), .B(n361), .ZN(n378) );
  INV_X1 U379 ( .A(KEYINPUT19), .ZN(n351) );
  NOR2_X1 U380 ( .A1(n624), .A2(n639), .ZN(n625) );
  NOR2_X1 U381 ( .A1(n640), .A2(n639), .ZN(n641) );
  BUF_X1 U382 ( .A(n632), .Z(n626) );
  XNOR2_X1 U383 ( .A(n352), .B(n351), .ZN(n528) );
  NOR2_X2 U384 ( .A1(n486), .A2(n485), .ZN(n352) );
  BUF_X1 U385 ( .A(n612), .Z(n353) );
  XNOR2_X1 U386 ( .A(n359), .B(n358), .ZN(n360) );
  INV_X2 U387 ( .A(G953), .ZN(n708) );
  INV_X1 U388 ( .A(KEYINPUT44), .ZN(n559) );
  AND2_X1 U389 ( .A1(n355), .A2(n354), .ZN(n507) );
  NOR2_X1 U390 ( .A1(n498), .A2(n433), .ZN(n434) );
  XNOR2_X1 U391 ( .A(n601), .B(KEYINPUT84), .ZN(n639) );
  INV_X1 U392 ( .A(KEYINPUT81), .ZN(n575) );
  XNOR2_X1 U393 ( .A(n506), .B(KEYINPUT73), .ZN(n354) );
  AND2_X1 U394 ( .A1(n497), .A2(n496), .ZN(n355) );
  NAND2_X1 U395 ( .A1(n593), .A2(n587), .ZN(n585) );
  XNOR2_X1 U396 ( .A(n584), .B(n583), .ZN(n593) );
  XNOR2_X1 U397 ( .A(n425), .B(n424), .ZN(n486) );
  BUF_X1 U398 ( .A(n549), .Z(n541) );
  XNOR2_X1 U399 ( .A(n405), .B(n442), .ZN(n408) );
  XNOR2_X1 U400 ( .A(n408), .B(n407), .ZN(n714) );
  AND2_X1 U401 ( .A1(n568), .A2(n562), .ZN(n565) );
  XOR2_X1 U402 ( .A(G140), .B(KEYINPUT98), .Z(n356) );
  XOR2_X1 U403 ( .A(n384), .B(n383), .Z(n357) );
  INV_X1 U404 ( .A(KEYINPUT12), .ZN(n436) );
  NOR2_X1 U405 ( .A1(n550), .A2(n477), .ZN(n478) );
  INV_X1 U406 ( .A(KEYINPUT48), .ZN(n509) );
  XNOR2_X1 U407 ( .A(n437), .B(n436), .ZN(n438) );
  NAND2_X1 U408 ( .A1(n605), .A2(n478), .ZN(n479) );
  XNOR2_X1 U409 ( .A(n509), .B(KEYINPUT78), .ZN(n510) );
  XNOR2_X1 U410 ( .A(n479), .B(KEYINPUT109), .ZN(n480) );
  XNOR2_X1 U411 ( .A(n511), .B(n510), .ZN(n520) );
  XNOR2_X1 U412 ( .A(n483), .B(KEYINPUT1), .ZN(n549) );
  BUF_X1 U413 ( .A(n714), .Z(n716) );
  BUF_X1 U414 ( .A(n593), .Z(n709) );
  XNOR2_X1 U415 ( .A(n493), .B(n476), .ZN(n605) );
  INV_X1 U416 ( .A(KEYINPUT63), .ZN(n603) );
  XNOR2_X2 U417 ( .A(G143), .B(G128), .ZN(n414) );
  XNOR2_X1 U418 ( .A(G131), .B(KEYINPUT68), .ZN(n359) );
  INV_X1 U419 ( .A(KEYINPUT4), .ZN(n358) );
  XNOR2_X1 U420 ( .A(KEYINPUT67), .B(G101), .ZN(n415) );
  XNOR2_X1 U421 ( .A(n415), .B(G146), .ZN(n361) );
  XOR2_X1 U422 ( .A(KEYINPUT94), .B(G116), .Z(n363) );
  XNOR2_X1 U423 ( .A(G137), .B(G113), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U425 ( .A(KEYINPUT3), .B(G119), .ZN(n406) );
  XNOR2_X1 U426 ( .A(n364), .B(n406), .ZN(n367) );
  NOR2_X1 U427 ( .A1(G953), .A2(G237), .ZN(n443) );
  NAND2_X1 U428 ( .A1(n443), .A2(G210), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n365), .B(KEYINPUT5), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n378), .B(n368), .ZN(n598) );
  INV_X1 U432 ( .A(G902), .ZN(n460) );
  NAND2_X1 U433 ( .A1(n598), .A2(n460), .ZN(n369) );
  XNOR2_X2 U434 ( .A(n369), .B(G472), .ZN(n679) );
  NOR2_X1 U435 ( .A1(G237), .A2(G902), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n370), .B(KEYINPUT70), .ZN(n421) );
  INV_X1 U437 ( .A(G214), .ZN(n371) );
  OR2_X1 U438 ( .A1(n421), .A2(n371), .ZN(n687) );
  NAND2_X1 U439 ( .A1(n679), .A2(n687), .ZN(n372) );
  XOR2_X1 U440 ( .A(n372), .B(KEYINPUT30), .Z(n400) );
  XNOR2_X1 U441 ( .A(G137), .B(G140), .ZN(n388) );
  XNOR2_X1 U442 ( .A(G107), .B(n388), .ZN(n374) );
  NAND2_X1 U443 ( .A1(G227), .A2(n708), .ZN(n373) );
  XNOR2_X1 U444 ( .A(n374), .B(n373), .ZN(n376) );
  XNOR2_X1 U445 ( .A(G104), .B(G110), .ZN(n375) );
  XNOR2_X1 U446 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U447 ( .A(n378), .B(n377), .ZN(n628) );
  NAND2_X1 U448 ( .A1(n628), .A2(n460), .ZN(n379) );
  XNOR2_X2 U449 ( .A(n379), .B(G469), .ZN(n483) );
  INV_X1 U450 ( .A(n483), .ZN(n468) );
  NAND2_X1 U451 ( .A1(G234), .A2(n708), .ZN(n380) );
  XOR2_X1 U452 ( .A(KEYINPUT8), .B(n380), .Z(n455) );
  AND2_X1 U453 ( .A1(G221), .A2(n455), .ZN(n387) );
  XOR2_X1 U454 ( .A(KEYINPUT88), .B(G110), .Z(n382) );
  XNOR2_X1 U455 ( .A(G128), .B(G119), .ZN(n381) );
  XNOR2_X1 U456 ( .A(n382), .B(n381), .ZN(n385) );
  XOR2_X1 U457 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n384) );
  XNOR2_X1 U458 ( .A(KEYINPUT23), .B(KEYINPUT90), .ZN(n383) );
  XNOR2_X1 U459 ( .A(n385), .B(n357), .ZN(n386) );
  XNOR2_X1 U460 ( .A(n387), .B(n386), .ZN(n389) );
  XNOR2_X2 U461 ( .A(G146), .B(G125), .ZN(n410) );
  XNOR2_X1 U462 ( .A(n410), .B(KEYINPUT10), .ZN(n440) );
  XNOR2_X1 U463 ( .A(n388), .B(n440), .ZN(n721) );
  XNOR2_X1 U464 ( .A(n389), .B(n721), .ZN(n615) );
  NAND2_X1 U465 ( .A1(n615), .A2(n460), .ZN(n396) );
  XOR2_X1 U466 ( .A(KEYINPUT92), .B(KEYINPUT20), .Z(n391) );
  XNOR2_X1 U467 ( .A(KEYINPUT15), .B(G902), .ZN(n419) );
  NAND2_X1 U468 ( .A1(G234), .A2(n419), .ZN(n390) );
  XNOR2_X1 U469 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U470 ( .A(KEYINPUT91), .B(n392), .ZN(n397) );
  NAND2_X1 U471 ( .A1(n397), .A2(G217), .ZN(n394) );
  XNOR2_X1 U472 ( .A(KEYINPUT25), .B(KEYINPUT93), .ZN(n393) );
  XNOR2_X1 U473 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X2 U474 ( .A(n396), .B(n395), .ZN(n542) );
  NAND2_X1 U475 ( .A1(n397), .A2(G221), .ZN(n399) );
  INV_X1 U476 ( .A(KEYINPUT21), .ZN(n398) );
  XNOR2_X1 U477 ( .A(n399), .B(n398), .ZN(n673) );
  NAND2_X1 U478 ( .A1(n542), .A2(n673), .ZN(n669) );
  NOR2_X1 U479 ( .A1(n468), .A2(n669), .ZN(n567) );
  NAND2_X1 U480 ( .A1(n400), .A2(n567), .ZN(n498) );
  XNOR2_X2 U481 ( .A(KEYINPUT69), .B(KEYINPUT16), .ZN(n401) );
  XNOR2_X1 U482 ( .A(n401), .B(G110), .ZN(n402) );
  INV_X1 U483 ( .A(n402), .ZN(n405) );
  XNOR2_X2 U484 ( .A(G122), .B(G113), .ZN(n404) );
  INV_X1 U485 ( .A(G104), .ZN(n403) );
  XNOR2_X2 U486 ( .A(n404), .B(n403), .ZN(n442) );
  XNOR2_X1 U487 ( .A(G116), .B(G107), .ZN(n450) );
  XNOR2_X1 U488 ( .A(n450), .B(n406), .ZN(n407) );
  XNOR2_X1 U489 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n409) );
  XNOR2_X1 U490 ( .A(n410), .B(n409), .ZN(n413) );
  NAND2_X1 U491 ( .A1(n708), .A2(G224), .ZN(n411) );
  XNOR2_X1 U492 ( .A(n411), .B(KEYINPUT4), .ZN(n412) );
  XNOR2_X1 U493 ( .A(n413), .B(n412), .ZN(n417) );
  XNOR2_X1 U494 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U495 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U496 ( .A(n714), .B(n418), .ZN(n633) );
  INV_X1 U497 ( .A(n419), .ZN(n587) );
  OR2_X2 U498 ( .A1(n633), .A2(n587), .ZN(n425) );
  INV_X1 U499 ( .A(G210), .ZN(n420) );
  OR2_X1 U500 ( .A1(n421), .A2(n420), .ZN(n423) );
  INV_X1 U501 ( .A(KEYINPUT85), .ZN(n422) );
  XNOR2_X1 U502 ( .A(n423), .B(n422), .ZN(n424) );
  BUF_X1 U503 ( .A(n486), .Z(n481) );
  XNOR2_X1 U504 ( .A(n481), .B(KEYINPUT38), .ZN(n688) );
  INV_X1 U505 ( .A(n688), .ZN(n432) );
  NAND2_X1 U506 ( .A1(G234), .A2(G237), .ZN(n426) );
  XNOR2_X1 U507 ( .A(n426), .B(KEYINPUT14), .ZN(n427) );
  NAND2_X1 U508 ( .A1(G952), .A2(n427), .ZN(n701) );
  NOR2_X1 U509 ( .A1(n701), .A2(G953), .ZN(n524) );
  NAND2_X1 U510 ( .A1(n427), .A2(G902), .ZN(n428) );
  XOR2_X1 U511 ( .A(KEYINPUT86), .B(n428), .Z(n521) );
  NAND2_X1 U512 ( .A1(n521), .A2(G953), .ZN(n429) );
  NOR2_X1 U513 ( .A1(G900), .A2(n429), .ZN(n430) );
  NOR2_X1 U514 ( .A1(n524), .A2(n430), .ZN(n431) );
  XNOR2_X1 U515 ( .A(KEYINPUT72), .B(n431), .ZN(n499) );
  OR2_X1 U516 ( .A1(n432), .A2(n499), .ZN(n433) );
  XNOR2_X1 U517 ( .A(n434), .B(KEYINPUT39), .ZN(n518) );
  XNOR2_X1 U518 ( .A(KEYINPUT11), .B(KEYINPUT99), .ZN(n435) );
  XNOR2_X1 U519 ( .A(n356), .B(n435), .ZN(n439) );
  XNOR2_X1 U520 ( .A(G131), .B(G143), .ZN(n437) );
  XNOR2_X1 U521 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U522 ( .A(n441), .B(n440), .ZN(n446) );
  NAND2_X1 U523 ( .A1(G214), .A2(n443), .ZN(n444) );
  XNOR2_X1 U524 ( .A(n442), .B(n444), .ZN(n445) );
  XNOR2_X1 U525 ( .A(n446), .B(n445), .ZN(n621) );
  NAND2_X1 U526 ( .A1(n621), .A2(n460), .ZN(n448) );
  XOR2_X1 U527 ( .A(KEYINPUT13), .B(G475), .Z(n447) );
  XNOR2_X1 U528 ( .A(n448), .B(n447), .ZN(n470) );
  INV_X1 U529 ( .A(KEYINPUT101), .ZN(n449) );
  XNOR2_X1 U530 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U531 ( .A(n452), .B(n451), .ZN(n459) );
  XOR2_X1 U532 ( .A(KEYINPUT100), .B(KEYINPUT7), .Z(n454) );
  XNOR2_X1 U533 ( .A(G122), .B(KEYINPUT9), .ZN(n453) );
  XNOR2_X1 U534 ( .A(n454), .B(n453), .ZN(n457) );
  NAND2_X1 U535 ( .A1(G217), .A2(n455), .ZN(n456) );
  XNOR2_X1 U536 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U537 ( .A(n459), .B(n458), .ZN(n618) );
  NAND2_X1 U538 ( .A1(n618), .A2(n460), .ZN(n462) );
  XOR2_X1 U539 ( .A(KEYINPUT102), .B(G478), .Z(n461) );
  XNOR2_X1 U540 ( .A(n462), .B(n461), .ZN(n489) );
  NAND2_X1 U541 ( .A1(n470), .A2(n489), .ZN(n493) );
  NOR2_X1 U542 ( .A1(n518), .A2(n493), .ZN(n463) );
  XOR2_X1 U543 ( .A(KEYINPUT40), .B(n463), .Z(n734) );
  INV_X1 U544 ( .A(n679), .ZN(n566) );
  INV_X1 U545 ( .A(n542), .ZN(n466) );
  INV_X1 U546 ( .A(n673), .ZN(n464) );
  NOR2_X1 U547 ( .A1(n464), .A2(n499), .ZN(n465) );
  NAND2_X1 U548 ( .A1(n466), .A2(n465), .ZN(n477) );
  NOR2_X1 U549 ( .A1(n566), .A2(n477), .ZN(n467) );
  XOR2_X1 U550 ( .A(KEYINPUT28), .B(n467), .Z(n469) );
  NOR2_X1 U551 ( .A1(n469), .A2(n468), .ZN(n487) );
  INV_X1 U552 ( .A(n489), .ZN(n500) );
  OR2_X1 U553 ( .A1(n470), .A2(n500), .ZN(n690) );
  INV_X1 U554 ( .A(n690), .ZN(n532) );
  NAND2_X1 U555 ( .A1(n688), .A2(n687), .ZN(n471) );
  XNOR2_X1 U556 ( .A(KEYINPUT113), .B(n471), .ZN(n685) );
  NAND2_X1 U557 ( .A1(n532), .A2(n685), .ZN(n472) );
  XNOR2_X1 U558 ( .A(n472), .B(KEYINPUT41), .ZN(n702) );
  NAND2_X1 U559 ( .A1(n487), .A2(n702), .ZN(n473) );
  XNOR2_X1 U560 ( .A(n473), .B(KEYINPUT42), .ZN(n735) );
  NAND2_X1 U561 ( .A1(n734), .A2(n735), .ZN(n475) );
  XNOR2_X1 U562 ( .A(KEYINPUT46), .B(KEYINPUT79), .ZN(n474) );
  XNOR2_X1 U563 ( .A(n475), .B(n474), .ZN(n508) );
  INV_X1 U564 ( .A(KEYINPUT108), .ZN(n476) );
  XNOR2_X1 U565 ( .A(n679), .B(KEYINPUT6), .ZN(n550) );
  NAND2_X1 U566 ( .A1(n480), .A2(n687), .ZN(n512) );
  NOR2_X1 U567 ( .A1(n512), .A2(n481), .ZN(n482) );
  XNOR2_X1 U568 ( .A(n482), .B(KEYINPUT36), .ZN(n484) );
  XOR2_X1 U569 ( .A(KEYINPUT83), .B(n541), .Z(n538) );
  NAND2_X1 U570 ( .A1(n484), .A2(n538), .ZN(n656) );
  XNOR2_X1 U571 ( .A(n656), .B(KEYINPUT80), .ZN(n497) );
  INV_X1 U572 ( .A(n687), .ZN(n485) );
  NAND2_X1 U573 ( .A1(n487), .A2(n528), .ZN(n488) );
  XNOR2_X1 U574 ( .A(n488), .B(KEYINPUT71), .ZN(n651) );
  XOR2_X1 U575 ( .A(n651), .B(KEYINPUT47), .Z(n495) );
  INV_X1 U576 ( .A(KEYINPUT103), .ZN(n491) );
  OR2_X1 U577 ( .A1(n470), .A2(n489), .ZN(n490) );
  XOR2_X1 U578 ( .A(n491), .B(n490), .Z(n646) );
  INV_X1 U579 ( .A(KEYINPUT104), .ZN(n492) );
  XNOR2_X1 U580 ( .A(n646), .B(n492), .ZN(n517) );
  NAND2_X1 U581 ( .A1(n517), .A2(n493), .ZN(n686) );
  INV_X1 U582 ( .A(n686), .ZN(n573) );
  NAND2_X1 U583 ( .A1(n651), .A2(n573), .ZN(n494) );
  NAND2_X1 U584 ( .A1(n495), .A2(n494), .ZN(n496) );
  NAND2_X1 U585 ( .A1(n573), .A2(KEYINPUT47), .ZN(n505) );
  NOR2_X1 U586 ( .A1(n499), .A2(n498), .ZN(n503) );
  NAND2_X1 U587 ( .A1(n470), .A2(n500), .ZN(n501) );
  XOR2_X1 U588 ( .A(KEYINPUT107), .B(n501), .Z(n555) );
  NOR2_X1 U589 ( .A1(n555), .A2(n481), .ZN(n502) );
  NAND2_X1 U590 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U591 ( .A(n504), .B(KEYINPUT112), .ZN(n733) );
  NAND2_X1 U592 ( .A1(n505), .A2(n733), .ZN(n506) );
  NAND2_X1 U593 ( .A1(n508), .A2(n507), .ZN(n511) );
  XNOR2_X1 U594 ( .A(KEYINPUT110), .B(n512), .ZN(n513) );
  NOR2_X1 U595 ( .A1(n541), .A2(n513), .ZN(n514) );
  XNOR2_X1 U596 ( .A(KEYINPUT111), .B(n514), .ZN(n515) );
  XNOR2_X1 U597 ( .A(n515), .B(KEYINPUT43), .ZN(n516) );
  AND2_X1 U598 ( .A1(n516), .A2(n481), .ZN(n610) );
  NOR2_X1 U599 ( .A1(n518), .A2(n517), .ZN(n659) );
  NOR2_X1 U600 ( .A1(n610), .A2(n659), .ZN(n519) );
  NAND2_X1 U601 ( .A1(n520), .A2(n519), .ZN(n725) );
  NOR2_X1 U602 ( .A1(G898), .A2(n708), .ZN(n718) );
  NAND2_X1 U603 ( .A1(n718), .A2(n521), .ZN(n523) );
  INV_X1 U604 ( .A(KEYINPUT87), .ZN(n522) );
  XNOR2_X1 U605 ( .A(n523), .B(n522), .ZN(n526) );
  INV_X1 U606 ( .A(n524), .ZN(n525) );
  NAND2_X1 U607 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U608 ( .A1(n528), .A2(n527), .ZN(n531) );
  INV_X1 U609 ( .A(KEYINPUT82), .ZN(n529) );
  XNOR2_X1 U610 ( .A(n529), .B(KEYINPUT0), .ZN(n530) );
  XNOR2_X2 U611 ( .A(n531), .B(n530), .ZN(n568) );
  AND2_X1 U612 ( .A1(n532), .A2(n673), .ZN(n533) );
  NAND2_X1 U613 ( .A1(n568), .A2(n533), .ZN(n535) );
  INV_X1 U614 ( .A(KEYINPUT22), .ZN(n534) );
  NAND2_X1 U615 ( .A1(n544), .A2(n550), .ZN(n576) );
  INV_X1 U616 ( .A(KEYINPUT105), .ZN(n536) );
  XNOR2_X1 U617 ( .A(n542), .B(n536), .ZN(n672) );
  INV_X1 U618 ( .A(n672), .ZN(n537) );
  NAND2_X1 U619 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X2 U620 ( .A1(n576), .A2(n539), .ZN(n540) );
  INV_X1 U621 ( .A(n541), .ZN(n670) );
  NOR2_X1 U622 ( .A1(n679), .A2(n542), .ZN(n543) );
  NAND2_X1 U623 ( .A1(n670), .A2(n543), .ZN(n547) );
  BUF_X1 U624 ( .A(n544), .Z(n545) );
  INV_X1 U625 ( .A(n545), .ZN(n546) );
  NOR2_X1 U626 ( .A1(n547), .A2(n546), .ZN(n607) );
  NOR2_X1 U627 ( .A1(n612), .A2(n607), .ZN(n558) );
  INV_X1 U628 ( .A(n669), .ZN(n548) );
  NAND2_X1 U629 ( .A1(n549), .A2(n548), .ZN(n561) );
  NOR2_X1 U630 ( .A1(n561), .A2(n550), .ZN(n552) );
  INV_X1 U631 ( .A(KEYINPUT33), .ZN(n551) );
  XNOR2_X1 U632 ( .A(n552), .B(n551), .ZN(n694) );
  AND2_X1 U633 ( .A1(n694), .A2(n568), .ZN(n554) );
  INV_X1 U634 ( .A(KEYINPUT34), .ZN(n553) );
  XNOR2_X1 U635 ( .A(n554), .B(n553), .ZN(n556) );
  NOR2_X1 U636 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U637 ( .A(n557), .B(KEYINPUT35), .ZN(n611) );
  NAND2_X1 U638 ( .A1(n558), .A2(n611), .ZN(n560) );
  XNOR2_X1 U639 ( .A(n560), .B(n559), .ZN(n582) );
  INV_X1 U640 ( .A(n681), .ZN(n562) );
  XNOR2_X1 U641 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n563) );
  XNOR2_X1 U642 ( .A(n563), .B(KEYINPUT95), .ZN(n564) );
  XNOR2_X1 U643 ( .A(n565), .B(n564), .ZN(n653) );
  NAND2_X1 U644 ( .A1(n567), .A2(n566), .ZN(n570) );
  INV_X1 U645 ( .A(n568), .ZN(n569) );
  NOR2_X1 U646 ( .A1(n570), .A2(n569), .ZN(n642) );
  NOR2_X1 U647 ( .A1(n653), .A2(n642), .ZN(n572) );
  INV_X1 U648 ( .A(KEYINPUT97), .ZN(n571) );
  XNOR2_X1 U649 ( .A(n572), .B(n571), .ZN(n574) );
  NOR2_X1 U650 ( .A1(n574), .A2(n573), .ZN(n579) );
  XNOR2_X1 U651 ( .A(n576), .B(n575), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n670), .A2(n672), .ZN(n577) );
  NOR2_X1 U653 ( .A1(n578), .A2(n577), .ZN(n609) );
  NOR2_X1 U654 ( .A1(n579), .A2(n609), .ZN(n580) );
  XNOR2_X1 U655 ( .A(n580), .B(KEYINPUT106), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U657 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n583) );
  XNOR2_X1 U658 ( .A(n585), .B(KEYINPUT76), .ZN(n586) );
  NOR2_X1 U659 ( .A1(n725), .A2(n586), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n587), .A2(KEYINPUT2), .ZN(n588) );
  XOR2_X1 U661 ( .A(KEYINPUT66), .B(n588), .Z(n589) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n591), .B(KEYINPUT65), .ZN(n597) );
  INV_X1 U664 ( .A(n725), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n592), .A2(KEYINPUT2), .ZN(n595) );
  INV_X1 U666 ( .A(n709), .ZN(n594) );
  NOR2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n661) );
  INV_X1 U668 ( .A(n661), .ZN(n596) );
  AND2_X2 U669 ( .A1(n597), .A2(n596), .ZN(n632) );
  NAND2_X1 U670 ( .A1(n632), .A2(G472), .ZN(n600) );
  XOR2_X1 U671 ( .A(KEYINPUT62), .B(n598), .Z(n599) );
  XNOR2_X1 U672 ( .A(n600), .B(n599), .ZN(n602) );
  NOR2_X1 U673 ( .A1(n708), .A2(G952), .ZN(n601) );
  XNOR2_X1 U674 ( .A(n604), .B(n603), .ZN(G57) );
  NAND2_X1 U675 ( .A1(n642), .A2(n605), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n606), .B(G104), .ZN(G6) );
  XOR2_X1 U677 ( .A(G110), .B(n607), .Z(G12) );
  NAND2_X1 U678 ( .A1(n653), .A2(n646), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n608), .B(G116), .ZN(G18) );
  XOR2_X1 U680 ( .A(G101), .B(n609), .Z(G3) );
  XOR2_X1 U681 ( .A(n610), .B(G140), .Z(G42) );
  XNOR2_X1 U682 ( .A(n611), .B(G122), .ZN(G24) );
  XOR2_X1 U683 ( .A(G119), .B(n353), .Z(G21) );
  BUF_X1 U684 ( .A(n632), .Z(n613) );
  NAND2_X1 U685 ( .A1(n613), .A2(G217), .ZN(n614) );
  XOR2_X1 U686 ( .A(n615), .B(n614), .Z(n616) );
  NOR2_X1 U687 ( .A1(n616), .A2(n639), .ZN(G66) );
  NAND2_X1 U688 ( .A1(n626), .A2(G478), .ZN(n617) );
  XOR2_X1 U689 ( .A(n618), .B(n617), .Z(n619) );
  NOR2_X1 U690 ( .A1(n619), .A2(n639), .ZN(G63) );
  NAND2_X1 U691 ( .A1(n632), .A2(G475), .ZN(n623) );
  XOR2_X1 U692 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n620) );
  XNOR2_X1 U693 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U694 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U696 ( .A1(n626), .A2(G469), .ZN(n630) );
  XNOR2_X1 U697 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X1 U700 ( .A1(n631), .A2(n639), .ZN(G54) );
  NAND2_X1 U701 ( .A1(n632), .A2(G210), .ZN(n638) );
  BUF_X1 U702 ( .A(n633), .Z(n634) );
  XNOR2_X1 U703 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n635) );
  XOR2_X1 U704 ( .A(n635), .B(KEYINPUT55), .Z(n636) );
  XNOR2_X1 U705 ( .A(n634), .B(n636), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n638), .B(n637), .ZN(n640) );
  XNOR2_X1 U707 ( .A(n641), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U708 ( .A1(n642), .A2(n646), .ZN(n644) );
  XOR2_X1 U709 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n643) );
  XNOR2_X1 U710 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U711 ( .A(G107), .B(n645), .ZN(G9) );
  XOR2_X1 U712 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n648) );
  NAND2_X1 U713 ( .A1(n651), .A2(n646), .ZN(n647) );
  XNOR2_X1 U714 ( .A(n648), .B(n647), .ZN(n650) );
  XOR2_X1 U715 ( .A(G128), .B(KEYINPUT114), .Z(n649) );
  XNOR2_X1 U716 ( .A(n650), .B(n649), .ZN(G30) );
  NAND2_X1 U717 ( .A1(n605), .A2(n651), .ZN(n652) );
  XNOR2_X1 U718 ( .A(n652), .B(G146), .ZN(G48) );
  NAND2_X1 U719 ( .A1(n653), .A2(n605), .ZN(n654) );
  XNOR2_X1 U720 ( .A(n654), .B(KEYINPUT116), .ZN(n655) );
  XNOR2_X1 U721 ( .A(G113), .B(n655), .ZN(G15) );
  XNOR2_X1 U722 ( .A(KEYINPUT37), .B(KEYINPUT117), .ZN(n657) );
  XNOR2_X1 U723 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U724 ( .A(G125), .B(n658), .ZN(G27) );
  XOR2_X1 U725 ( .A(G134), .B(n659), .Z(G36) );
  XNOR2_X1 U726 ( .A(KEYINPUT2), .B(KEYINPUT74), .ZN(n662) );
  NOR2_X1 U727 ( .A1(n709), .A2(n662), .ZN(n660) );
  NOR2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n666) );
  INV_X1 U729 ( .A(n662), .ZN(n663) );
  NAND2_X1 U730 ( .A1(n663), .A2(n725), .ZN(n664) );
  XOR2_X1 U731 ( .A(KEYINPUT75), .B(n664), .Z(n665) );
  NAND2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U733 ( .A(KEYINPUT77), .B(n667), .ZN(n668) );
  NOR2_X1 U734 ( .A1(G953), .A2(n668), .ZN(n706) );
  NAND2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U736 ( .A(KEYINPUT50), .B(n671), .ZN(n677) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n675) );
  XNOR2_X1 U738 ( .A(KEYINPUT118), .B(KEYINPUT49), .ZN(n674) );
  XNOR2_X1 U739 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U741 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U742 ( .A(n680), .B(KEYINPUT119), .ZN(n682) );
  NAND2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U744 ( .A(KEYINPUT51), .B(n683), .Z(n684) );
  NAND2_X1 U745 ( .A1(n684), .A2(n702), .ZN(n697) );
  NAND2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n693) );
  NOR2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U749 ( .A(KEYINPUT120), .B(n691), .Z(n692) );
  NAND2_X1 U750 ( .A1(n693), .A2(n692), .ZN(n695) );
  NAND2_X1 U751 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U752 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n698), .B(KEYINPUT52), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n699), .B(KEYINPUT121), .ZN(n700) );
  NOR2_X1 U755 ( .A1(n701), .A2(n700), .ZN(n704) );
  AND2_X1 U756 ( .A1(n694), .A2(n702), .ZN(n703) );
  NOR2_X1 U757 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U758 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U759 ( .A(KEYINPUT53), .B(n707), .Z(G75) );
  NAND2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U761 ( .A1(G953), .A2(G224), .ZN(n710) );
  XNOR2_X1 U762 ( .A(KEYINPUT61), .B(n710), .ZN(n711) );
  NAND2_X1 U763 ( .A1(n711), .A2(G898), .ZN(n712) );
  NAND2_X1 U764 ( .A1(n713), .A2(n712), .ZN(n720) );
  XOR2_X1 U765 ( .A(G101), .B(KEYINPUT124), .Z(n715) );
  XNOR2_X1 U766 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U767 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U768 ( .A(n720), .B(n719), .ZN(G69) );
  XNOR2_X1 U769 ( .A(n722), .B(n721), .ZN(n723) );
  XOR2_X1 U770 ( .A(n723), .B(KEYINPUT125), .Z(n728) );
  XOR2_X1 U771 ( .A(n728), .B(KEYINPUT126), .Z(n724) );
  XNOR2_X1 U772 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U773 ( .A1(G953), .A2(n726), .ZN(n727) );
  XNOR2_X1 U774 ( .A(n727), .B(KEYINPUT127), .ZN(n732) );
  XNOR2_X1 U775 ( .A(G227), .B(n728), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n729), .A2(G900), .ZN(n730) );
  NAND2_X1 U777 ( .A1(G953), .A2(n730), .ZN(n731) );
  NAND2_X1 U778 ( .A1(n732), .A2(n731), .ZN(G72) );
  XNOR2_X1 U779 ( .A(G143), .B(n733), .ZN(G45) );
  XNOR2_X1 U780 ( .A(n734), .B(G131), .ZN(G33) );
  XNOR2_X1 U781 ( .A(G137), .B(n735), .ZN(G39) );
endmodule

