//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n855, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(KEYINPUT22), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT2), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT77), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(G148gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT76), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n214), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G155gat), .B(G162gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n211), .A2(KEYINPUT77), .A3(KEYINPUT2), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n215), .A3(G148gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G141gat), .B(G148gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(KEYINPUT2), .ZN(new_n227));
  NOR2_X1   g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT75), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT75), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G155gat), .B2(G162gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n231), .A3(new_n211), .ZN(new_n232));
  OAI22_X1  g031(.A1(new_n221), .A2(new_n225), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n210), .B1(new_n234), .B2(KEYINPUT29), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n235), .A2(KEYINPUT82), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(new_n210), .B2(KEYINPUT29), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n238), .A2(new_n233), .B1(G228gat), .B2(G233gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(KEYINPUT82), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT78), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n233), .A2(new_n242), .ZN(new_n243));
  OAI221_X1 g042(.A(KEYINPUT78), .B1(new_n227), .B2(new_n232), .C1(new_n221), .C2(new_n225), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n238), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n235), .ZN(new_n246));
  OAI211_X1 g045(.A(G228gat), .B(G233gat), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n203), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G78gat), .B(G106gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G22gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n241), .A2(new_n247), .A3(new_n203), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n251), .ZN(new_n254));
  INV_X1    g053(.A(new_n252), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(new_n248), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT32), .ZN(new_n258));
  INV_X1    g057(.A(G183gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT27), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT27), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G183gat), .ZN(new_n262));
  INV_X1    g061(.A(G190gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT64), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n261), .A2(G183gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n259), .A2(KEYINPUT27), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT65), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n260), .A2(new_n262), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n265), .A2(G190gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT64), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n264), .A2(new_n275), .A3(new_n265), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n267), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n259), .A2(new_n263), .ZN(new_n278));
  AND2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT26), .ZN(new_n281));
  AOI211_X1 g080(.A(new_n278), .B(new_n281), .C1(KEYINPUT26), .C2(new_n280), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(KEYINPUT24), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(new_n279), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n259), .A2(new_n263), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT24), .A3(new_n284), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n286), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT25), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n286), .A2(new_n290), .A3(KEYINPUT25), .A4(new_n292), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n283), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G134gat), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G127gat), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT66), .ZN(new_n303));
  INV_X1    g102(.A(G120gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G113gat), .ZN(new_n305));
  INV_X1    g104(.A(G113gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G120gat), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT1), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n300), .A2(KEYINPUT66), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n303), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n301), .A2(G127gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n299), .A2(G134gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT67), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n300), .A2(new_n302), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n308), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT68), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n313), .A2(KEYINPUT68), .A3(new_n308), .A4(new_n315), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n310), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT69), .B1(new_n298), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n277), .A2(new_n282), .B1(new_n295), .B2(new_n296), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n320), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n298), .A2(new_n321), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n258), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT33), .B1(new_n327), .B2(new_n329), .ZN(new_n331));
  XOR2_X1   g130(.A(G15gat), .B(G43gat), .Z(new_n332));
  XNOR2_X1  g131(.A(G71gat), .B(G99gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OR3_X1    g134(.A1(new_n330), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n322), .A2(new_n328), .A3(new_n325), .A4(new_n326), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT70), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT34), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n339), .A2(KEYINPUT34), .ZN(new_n341));
  AOI221_X4 g140(.A(new_n258), .B1(KEYINPUT33), .B2(new_n334), .C1(new_n327), .C2(new_n329), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n336), .A2(new_n340), .A3(new_n341), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n340), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n330), .A2(new_n331), .A3(new_n335), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(new_n342), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n257), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n320), .A2(new_n234), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT3), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(KEYINPUT5), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT4), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n318), .A2(new_n319), .ZN(new_n358));
  INV_X1    g157(.A(new_n225), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n226), .A2(KEYINPUT76), .B1(new_n213), .B2(new_n212), .ZN(new_n360));
  OR2_X1    g159(.A1(new_n226), .A2(KEYINPUT2), .ZN(new_n361));
  INV_X1    g160(.A(new_n232), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n359), .A2(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n310), .ZN(new_n364));
  AND4_X1   g163(.A1(new_n357), .A2(new_n358), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n357), .B1(new_n320), .B2(new_n363), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT80), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n358), .A2(new_n363), .A3(new_n364), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT4), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n358), .A2(new_n357), .A3(new_n363), .A4(new_n364), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n353), .B(new_n356), .C1(new_n367), .C2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n320), .A2(KEYINPUT79), .A3(new_n357), .A4(new_n363), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n370), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n355), .B1(new_n350), .B2(new_n351), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT5), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n243), .A2(new_n244), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n369), .B1(new_n381), .B2(new_n320), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n382), .B2(new_n355), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n373), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G1gat), .B(G29gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT0), .ZN(new_n387));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(KEYINPUT6), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT80), .B1(new_n365), .B2(new_n366), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n370), .A2(new_n368), .A3(new_n371), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n352), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n394), .A2(new_n356), .B1(new_n379), .B2(new_n383), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n396), .A3(new_n389), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n385), .A2(new_n390), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n396), .B1(new_n395), .B2(new_n389), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n391), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G226gat), .ZN(new_n403));
  INV_X1    g202(.A(G233gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n323), .B2(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n298), .A2(new_n405), .ZN(new_n408));
  INV_X1    g207(.A(new_n210), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT72), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT72), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n407), .A2(new_n408), .A3(new_n412), .A4(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT71), .B1(new_n407), .B2(new_n408), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT71), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT29), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n298), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(new_n406), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n210), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT73), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND2_X1  g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n425), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n414), .A2(new_n420), .A3(KEYINPUT30), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n420), .A3(new_n427), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n430), .A2(KEYINPUT74), .A3(new_n431), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n429), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n402), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT35), .B1(new_n349), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n391), .A2(KEYINPUT84), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n395), .A2(new_n389), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT6), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n439), .B(new_n442), .C1(new_n400), .C2(new_n401), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT35), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n348), .A2(new_n443), .A3(new_n444), .A4(new_n436), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n438), .A2(new_n445), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n344), .A2(KEYINPUT36), .A3(new_n347), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT36), .B1(new_n344), .B2(new_n347), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n391), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n398), .B1(new_n395), .B2(new_n389), .ZN(new_n451));
  AND4_X1   g250(.A1(new_n396), .A2(new_n373), .A3(new_n384), .A4(new_n389), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n401), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n430), .A2(KEYINPUT74), .A3(new_n431), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT74), .B1(new_n430), .B2(new_n431), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n426), .B(new_n428), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n257), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n414), .A2(new_n420), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n425), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n414), .B2(new_n420), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT38), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n407), .A2(new_n408), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n460), .B1(new_n465), .B2(new_n210), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n409), .B1(new_n415), .B2(new_n419), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT38), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(new_n461), .A3(new_n425), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT83), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n468), .A2(new_n461), .A3(new_n471), .A4(new_n425), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n464), .A2(new_n470), .A3(new_n430), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(new_n443), .ZN(new_n474));
  INV_X1    g273(.A(new_n257), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n353), .B1(new_n367), .B2(new_n372), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT39), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n355), .ZN(new_n478));
  INV_X1    g277(.A(new_n382), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n479), .B2(new_n354), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(new_n394), .B2(new_n354), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n481), .A3(new_n389), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT40), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n440), .B1(new_n483), .B2(new_n482), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n475), .B1(new_n486), .B2(new_n436), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n449), .B(new_n459), .C1(new_n474), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n446), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G113gat), .B(G141gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  XOR2_X1   g291(.A(G169gat), .B(G197gat), .Z(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(KEYINPUT12), .ZN(new_n495));
  INV_X1    g294(.A(G8gat), .ZN(new_n496));
  XOR2_X1   g295(.A(G15gat), .B(G22gat), .Z(new_n497));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G1gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT89), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n496), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n501), .B(new_n498), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n500), .A2(KEYINPUT16), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  OAI221_X1 g308(.A(new_n503), .B1(new_n504), .B2(new_n496), .C1(new_n506), .C2(new_n507), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT87), .B(G29gat), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT86), .B1(G29gat), .B2(G36gat), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n512), .A2(G36gat), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR3_X1    g315(.A1(KEYINPUT86), .A2(G29gat), .A3(G36gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT14), .A3(new_n513), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G43gat), .B(G50gat), .Z(new_n524));
  INV_X1    g323(.A(KEYINPUT15), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n516), .A2(new_n526), .A3(new_n521), .A4(new_n518), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n511), .A2(new_n528), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT13), .Z(new_n534));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT17), .B1(new_n528), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n537));
  AOI211_X1 g336(.A(KEYINPUT88), .B(new_n537), .C1(new_n523), .C2(new_n527), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n533), .B(new_n529), .C1(new_n539), .C2(new_n511), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n532), .A2(new_n534), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n527), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n521), .B1(new_n516), .B2(new_n518), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n535), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n537), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n535), .A3(KEYINPUT17), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n509), .A2(new_n510), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n533), .A4(new_n529), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n495), .B1(new_n542), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n540), .A2(new_n541), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n534), .B1(new_n530), .B2(new_n531), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n553), .A2(new_n551), .A3(new_n554), .A4(new_n495), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT91), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(new_n551), .A3(new_n554), .ZN(new_n558));
  INV_X1    g357(.A(new_n495), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(KEYINPUT91), .A3(new_n555), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n489), .A2(KEYINPUT92), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT92), .B1(new_n489), .B2(new_n563), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n567), .A2(KEYINPUT41), .ZN(new_n568));
  XNOR2_X1  g367(.A(G134gat), .B(G162gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G190gat), .B(G218gat), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n574));
  NAND2_X1  g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT7), .ZN(new_n576));
  XOR2_X1   g375(.A(G99gat), .B(G106gat), .Z(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n576), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n577), .B1(new_n576), .B2(new_n581), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n574), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n576), .A2(new_n581), .ZN(new_n586));
  INV_X1    g385(.A(new_n577), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(KEYINPUT97), .A3(new_n582), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT98), .B1(new_n539), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT98), .ZN(new_n592));
  INV_X1    g391(.A(new_n590), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n548), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n588), .A2(new_n582), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n528), .A2(new_n596), .B1(KEYINPUT41), .B2(new_n567), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n573), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  AOI211_X1 g398(.A(new_n572), .B(new_n599), .C1(new_n591), .C2(new_n594), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n571), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n592), .B1(new_n548), .B2(new_n593), .ZN(new_n602));
  AOI211_X1 g401(.A(KEYINPUT98), .B(new_n590), .C1(new_n546), .C2(new_n547), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n572), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n595), .A2(new_n573), .A3(new_n597), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n570), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT21), .ZN(new_n609));
  INV_X1    g408(.A(G64gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(G57gat), .ZN(new_n611));
  XOR2_X1   g410(.A(KEYINPUT94), .B(G57gat), .Z(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(new_n610), .ZN(new_n613));
  NAND2_X1  g412(.A1(G71gat), .A2(G78gat), .ZN(new_n614));
  OR2_X1    g413(.A1(G71gat), .A2(G78gat), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT9), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n615), .A2(new_n614), .ZN(new_n619));
  XNOR2_X1  g418(.A(G57gat), .B(G64gat), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n619), .B(KEYINPUT93), .C1(new_n616), .C2(new_n620), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n614), .B(new_n615), .C1(new_n620), .C2(new_n616), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT93), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n549), .B1(new_n609), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n609), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n626), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G127gat), .B(G155gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT96), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT95), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n632), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G183gat), .B(G211gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n630), .B(new_n637), .Z(new_n638));
  NAND2_X1  g437(.A1(new_n608), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n586), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n577), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n613), .A2(new_n617), .B1(new_n622), .B2(new_n623), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n586), .A2(new_n640), .A3(new_n587), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n621), .A4(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n625), .A2(new_n596), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT10), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n596), .A2(new_n643), .A3(KEYINPUT10), .A4(new_n621), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(G230gat), .ZN(new_n650));
  OAI22_X1  g449(.A1(new_n647), .A2(new_n649), .B1(new_n650), .B2(new_n404), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n404), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n645), .A2(new_n646), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n651), .A2(new_n653), .A3(new_n657), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n639), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n455), .B(KEYINPUT100), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n566), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(new_n500), .ZN(G1324gat));
  OAI211_X1 g465(.A(new_n458), .B(new_n662), .C1(new_n564), .C2(new_n565), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT102), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT102), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(G8gat), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT42), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(KEYINPUT103), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n668), .B2(new_n669), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n675));
  OAI221_X1 g474(.A(new_n670), .B1(new_n667), .B2(new_n672), .C1(new_n674), .C2(new_n675), .ZN(G1325gat));
  NOR2_X1   g475(.A1(new_n566), .A2(new_n663), .ZN(new_n677));
  INV_X1    g476(.A(new_n344), .ZN(new_n678));
  INV_X1    g477(.A(new_n347), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(G15gat), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n449), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G15gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT104), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n682), .B1(new_n677), .B2(new_n685), .ZN(G1326gat));
  NAND2_X1  g485(.A1(new_n677), .A2(new_n257), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT43), .B(G22gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  INV_X1    g488(.A(new_n566), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n608), .A2(new_n638), .A3(new_n661), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n664), .A2(new_n512), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  INV_X1    g493(.A(new_n608), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n489), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT44), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n552), .A2(new_n556), .ZN(new_n700));
  AOI211_X1 g499(.A(KEYINPUT91), .B(new_n495), .C1(new_n542), .C2(new_n551), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n557), .A2(new_n561), .A3(KEYINPUT105), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n661), .B(KEYINPUT106), .Z(new_n705));
  NOR3_X1   g504(.A1(new_n704), .A2(new_n638), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n608), .B1(new_n446), .B2(new_n488), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT107), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI221_X1 g508(.A(new_n475), .B1(new_n486), .B2(new_n436), .C1(new_n473), .C2(new_n443), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n459), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n437), .A2(KEYINPUT108), .A3(new_n257), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n710), .A2(new_n712), .A3(new_n449), .A4(new_n713), .ZN(new_n714));
  AOI211_X1 g513(.A(KEYINPUT44), .B(new_n608), .C1(new_n714), .C2(new_n446), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n698), .B(new_n706), .C1(new_n709), .C2(new_n715), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n716), .A2(KEYINPUT109), .A3(new_n664), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT109), .B1(new_n716), .B2(new_n664), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n512), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n694), .A2(new_n719), .ZN(G1328gat));
  AND2_X1   g519(.A1(new_n690), .A2(new_n691), .ZN(new_n721));
  INV_X1    g520(.A(G36gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n722), .A3(new_n458), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT46), .ZN(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n716), .B2(new_n436), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n721), .A2(new_n726), .A3(new_n722), .A4(new_n458), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(G1329gat));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n732));
  OAI21_X1  g531(.A(G43gat), .B1(new_n716), .B2(new_n449), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n680), .A2(G43gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n690), .A2(new_n691), .A3(new_n734), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n731), .B(new_n732), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  AND4_X1   g535(.A1(new_n729), .A2(new_n733), .A3(new_n730), .A4(new_n735), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1330gat));
  OAI21_X1  g537(.A(KEYINPUT112), .B1(new_n716), .B2(new_n475), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G50gat), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n716), .A2(KEYINPUT112), .A3(new_n475), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n475), .A2(G50gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT111), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n690), .A2(new_n691), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT48), .ZN(new_n746));
  OAI21_X1  g545(.A(G50gat), .B1(new_n716), .B2(new_n475), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(new_n745), .ZN(new_n748));
  OAI22_X1  g547(.A1(new_n742), .A2(new_n746), .B1(KEYINPUT48), .B2(new_n748), .ZN(G1331gat));
  NAND2_X1  g548(.A1(new_n712), .A2(new_n713), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n449), .B1(new_n474), .B2(new_n487), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n446), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n704), .ZN(new_n753));
  INV_X1    g552(.A(new_n705), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n753), .A2(new_n639), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n664), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(new_n612), .ZN(G1332gat));
  NOR2_X1   g559(.A1(new_n756), .A2(new_n436), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  AND2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n761), .B2(new_n762), .ZN(G1333gat));
  NOR3_X1   g564(.A1(new_n756), .A2(G71gat), .A3(new_n680), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n757), .A2(new_n683), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(G71gat), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n757), .A2(new_n257), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT114), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT113), .B(G78gat), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1335gat));
  NOR2_X1   g572(.A1(new_n753), .A2(new_n638), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n752), .A2(KEYINPUT51), .A3(new_n695), .A4(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n752), .A2(new_n695), .A3(new_n774), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n608), .B1(new_n714), .B2(new_n446), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n781), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n774), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n777), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n777), .A2(new_n780), .A3(new_n782), .A4(KEYINPUT116), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n661), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n664), .A2(G85gat), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n753), .A2(new_n638), .A3(new_n788), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n698), .B(new_n792), .C1(new_n709), .C2(new_n715), .ZN(new_n793));
  OAI21_X1  g592(.A(G85gat), .B1(new_n793), .B2(new_n664), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n790), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n789), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n785), .B2(new_n786), .ZN(new_n797));
  INV_X1    g596(.A(new_n794), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT117), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(G1336gat));
  OR2_X1    g599(.A1(new_n793), .A2(new_n436), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G92gat), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n754), .A2(G92gat), .A3(new_n436), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(new_n783), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n780), .A2(new_n775), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n801), .A2(G92gat), .B1(new_n806), .B2(new_n803), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(G1337gat));
  NOR3_X1   g608(.A1(new_n680), .A2(G99gat), .A3(new_n788), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n787), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G99gat), .B1(new_n793), .B2(new_n449), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1338gat));
  NOR3_X1   g612(.A1(new_n754), .A2(G106gat), .A3(new_n475), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT53), .B1(new_n783), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT118), .B1(new_n793), .B2(new_n475), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G106gat), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n793), .A2(KEYINPUT118), .A3(new_n475), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G106gat), .B1(new_n793), .B2(new_n475), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n806), .A2(new_n814), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1339gat));
  NAND4_X1  g623(.A1(new_n704), .A2(new_n638), .A3(new_n608), .A4(new_n788), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n645), .A2(new_n646), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n652), .B(new_n648), .C1(new_n827), .C2(KEYINPUT10), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n828), .A2(new_n651), .A3(KEYINPUT54), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  OAI221_X1 g629(.A(new_n830), .B1(new_n650), .B2(new_n404), .C1(new_n647), .C2(new_n649), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n658), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n826), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n651), .A3(KEYINPUT54), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n834), .A2(KEYINPUT55), .A3(new_n658), .A4(new_n831), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n833), .A2(new_n660), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n532), .A2(new_n534), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n533), .B1(new_n550), .B2(new_n529), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n494), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(new_n555), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n695), .A2(new_n836), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n702), .A2(new_n703), .A3(new_n836), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n661), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n841), .B1(new_n844), .B2(new_n608), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n825), .B1(new_n845), .B2(new_n638), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NOR4_X1   g646(.A1(new_n847), .A2(new_n458), .A3(new_n349), .A4(new_n664), .ZN(new_n848));
  AOI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n753), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n562), .A2(new_n306), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n848), .B2(new_n850), .ZN(G1340gat));
  AOI21_X1  g650(.A(G120gat), .B1(new_n848), .B2(new_n661), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n754), .A2(new_n304), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n848), .B2(new_n853), .ZN(G1341gat));
  NAND2_X1  g653(.A1(new_n848), .A2(new_n638), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(G127gat), .ZN(G1342gat));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n848), .B(new_n695), .C1(new_n857), .C2(new_n301), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n301), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n858), .B(new_n859), .ZN(G1343gat));
  NOR3_X1   g659(.A1(new_n664), .A2(new_n683), .A3(new_n458), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n846), .B2(new_n257), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  INV_X1    g662(.A(new_n638), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n836), .A2(new_n557), .A3(new_n561), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n695), .B1(new_n865), .B2(new_n843), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n864), .B1(new_n866), .B2(new_n841), .ZN(new_n867));
  AOI211_X1 g666(.A(new_n863), .B(new_n475), .C1(new_n867), .C2(new_n825), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n861), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G141gat), .B1(new_n869), .B2(new_n562), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n846), .A2(new_n257), .A3(new_n861), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n562), .A2(G141gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n753), .B(new_n861), .C1(new_n862), .C2(new_n868), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(G141gat), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n874), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n876), .B1(new_n879), .B2(KEYINPUT58), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n877), .A2(G141gat), .B1(new_n872), .B2(new_n873), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(KEYINPUT119), .A3(new_n871), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n875), .B1(new_n880), .B2(new_n882), .ZN(G1344gat));
  NAND2_X1  g682(.A1(new_n861), .A2(new_n661), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n847), .A2(new_n475), .A3(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n217), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n661), .A2(new_n886), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n662), .A2(KEYINPUT120), .A3(new_n562), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT120), .B1(new_n662), .B2(new_n562), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n865), .A2(new_n843), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n608), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n833), .A2(new_n660), .A3(new_n835), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT121), .B1(new_n608), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n836), .A2(new_n896), .A3(new_n607), .A4(new_n601), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n897), .A3(new_n840), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n638), .B1(new_n899), .B2(KEYINPUT122), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n893), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n891), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n257), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n895), .A2(new_n840), .A3(new_n897), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT122), .B1(new_n906), .B2(new_n866), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n864), .A3(new_n902), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n889), .A2(new_n890), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(KEYINPUT123), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n863), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n475), .A2(new_n863), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n846), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n884), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n916));
  OAI221_X1 g715(.A(new_n887), .B1(new_n869), .B2(new_n888), .C1(new_n915), .C2(new_n916), .ZN(G1345gat));
  OAI21_X1  g716(.A(G155gat), .B1(new_n869), .B2(new_n864), .ZN(new_n918));
  INV_X1    g717(.A(new_n872), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n864), .A2(G155gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G1346gat));
  OAI21_X1  g720(.A(G162gat), .B1(new_n869), .B2(new_n608), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n608), .A2(G162gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n919), .B2(new_n923), .ZN(G1347gat));
  NAND2_X1  g723(.A1(new_n846), .A2(new_n664), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(new_n436), .A3(new_n349), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(G169gat), .A3(new_n563), .ZN(new_n927));
  AOI21_X1  g726(.A(G169gat), .B1(new_n926), .B2(new_n753), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(G1348gat));
  AND3_X1   g728(.A1(new_n846), .A2(new_n348), .A3(new_n664), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n930), .A2(G176gat), .A3(new_n458), .A4(new_n705), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT124), .ZN(new_n932));
  AOI21_X1  g731(.A(G176gat), .B1(new_n926), .B2(new_n661), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(G1349gat));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n458), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n259), .B1(new_n935), .B2(new_n864), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n270), .A2(new_n272), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n926), .A2(new_n937), .A3(new_n638), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(G1350gat));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n930), .A2(new_n458), .A3(new_n695), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n944), .A3(G190gat), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n943), .B2(G190gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n942), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n947), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(KEYINPUT61), .A3(new_n945), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n948), .B(new_n950), .C1(G190gat), .C2(new_n943), .ZN(G1351gat));
  NOR4_X1   g750(.A1(new_n925), .A2(new_n436), .A3(new_n475), .A4(new_n683), .ZN(new_n952));
  INV_X1    g751(.A(G197gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n953), .A3(new_n753), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT126), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n912), .A2(new_n914), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n758), .A2(new_n436), .A3(new_n683), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n563), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G197gat), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n955), .A2(new_n959), .ZN(G1352gat));
  AOI21_X1  g759(.A(new_n475), .B1(new_n910), .B2(KEYINPUT123), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n903), .A2(new_n904), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT57), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n914), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n705), .B(new_n957), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n956), .A2(KEYINPUT127), .A3(new_n705), .A4(new_n957), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n968), .A3(G204gat), .ZN(new_n969));
  INV_X1    g768(.A(G204gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n952), .A2(new_n970), .A3(new_n661), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n969), .A2(new_n973), .ZN(G1353gat));
  NAND3_X1  g773(.A1(new_n952), .A2(new_n205), .A3(new_n638), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n638), .B(new_n957), .C1(new_n963), .C2(new_n964), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  NAND3_X1  g778(.A1(new_n952), .A2(new_n206), .A3(new_n695), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n956), .A2(new_n695), .A3(new_n957), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n981), .B2(new_n206), .ZN(G1355gat));
endmodule


