//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n607, new_n608, new_n610, new_n611, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n457), .A2(KEYINPUT68), .B1(G567), .B2(new_n453), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n458), .B1(KEYINPUT68), .B2(new_n457), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(KEYINPUT70), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n464), .A2(new_n469), .A3(G125), .ZN(new_n470));
  INV_X1    g045(.A(G113), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(new_n466), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n466), .A2(G2105), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n474), .A2(G137), .B1(G101), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n474), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(new_n467), .B2(new_n468), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n479), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT71), .Z(G162));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(new_n474), .B2(G138), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n487), .A2(new_n480), .A3(G138), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n464), .A2(new_n469), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT73), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT73), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n464), .A2(new_n469), .A3(new_n492), .A4(new_n489), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n488), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n480), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT72), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT72), .B1(new_n496), .B2(new_n497), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT74), .B(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n510), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  AND3_X1   g093(.A1(new_n505), .A2(KEYINPUT75), .A3(new_n506), .ZN(new_n519));
  AOI21_X1  g094(.A(KEYINPUT75), .B1(new_n505), .B2(new_n506), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI221_X1 g101(.A(new_n524), .B1(new_n514), .B2(new_n525), .C1(new_n526), .C2(new_n512), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n522), .A2(new_n527), .ZN(G168));
  INV_X1    g103(.A(new_n519), .ZN(new_n529));
  INV_X1    g104(.A(new_n520), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n529), .A2(G64), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n509), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n507), .A2(new_n511), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n511), .A2(G543), .ZN(new_n535));
  AOI22_X1  g110(.A1(G90), .A2(new_n534), .B1(new_n535), .B2(G52), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G171));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n512), .A2(new_n539), .B1(new_n514), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n529), .A2(new_n530), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n541), .B1(new_n545), .B2(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT76), .ZN(G188));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OR3_X1    g128(.A1(new_n514), .A2(KEYINPUT9), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT9), .B1(new_n514), .B2(new_n553), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT77), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n505), .A2(new_n506), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n561), .A2(G651), .B1(G91), .B2(new_n534), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n556), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n564));
  INV_X1    g139(.A(new_n533), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n564), .B1(new_n565), .B2(new_n536), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n533), .A2(new_n537), .A3(KEYINPUT78), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G74), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n570), .B1(new_n519), .B2(new_n520), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(G87), .B2(new_n534), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n511), .A2(G49), .A3(G543), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT79), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n559), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(G48), .B2(new_n535), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n512), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n512), .A2(new_n581), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT80), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n579), .A2(new_n582), .A3(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(new_n509), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n512), .A2(new_n588), .B1(new_n514), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n587), .A2(new_n592), .ZN(G290));
  AND3_X1   g168(.A1(new_n507), .A2(new_n511), .A3(G92), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n559), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G54), .B2(new_n535), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(G301), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G284));
  AOI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G321));
  MUX2_X1   g179(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g180(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g181(.A(new_n600), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g187(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n613));
  XNOR2_X1  g188(.A(G323), .B(new_n613), .ZN(G282));
  AND2_X1   g189(.A1(new_n464), .A2(new_n469), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n475), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n474), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n481), .A2(G123), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n480), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT83), .B(G2096), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n620), .A2(new_n621), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT84), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n644), .A2(G14), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(KEYINPUT85), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(KEYINPUT85), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(G401));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT86), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  NOR3_X1   g229(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT88), .B(KEYINPUT17), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(new_n652), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n652), .B1(new_n651), .B2(new_n654), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n651), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(new_n658), .ZN(new_n664));
  INV_X1    g239(.A(new_n660), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n664), .B1(new_n665), .B2(KEYINPUT87), .ZN(new_n666));
  OAI221_X1 g241(.A(new_n656), .B1(new_n658), .B2(new_n659), .C1(new_n662), .C2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n673), .B(new_n674), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n677), .B(new_n678), .C1(new_n672), .C2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT90), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G24), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n587), .A2(new_n592), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  INV_X1    g268(.A(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT92), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(KEYINPUT92), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n474), .A2(G131), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n481), .A2(G119), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n480), .A2(G107), .ZN(new_n700));
  OAI21_X1  g275(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n698), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT91), .B(G29), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G25), .B(new_n702), .S(new_n704), .Z(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT35), .B(G1991), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  NAND3_X1  g282(.A1(new_n696), .A2(new_n697), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n690), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n690), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n690), .A2(G6), .ZN(new_n714));
  INV_X1    g289(.A(G305), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n690), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT32), .B(G1981), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n690), .A2(G22), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT93), .Z(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G303), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1971), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n713), .A2(new_n718), .A3(new_n719), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT34), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n708), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT36), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n704), .A2(G35), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n704), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT29), .Z(new_n730));
  INV_X1    g305(.A(G2090), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT100), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n731), .ZN(new_n734));
  NAND2_X1  g309(.A1(G160), .A2(G29), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT24), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G34), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(G34), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n703), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(G2084), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT98), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n703), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n474), .A2(G140), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT94), .Z(new_n746));
  OAI21_X1  g321(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n747));
  INV_X1    g322(.A(G116), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G2105), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n481), .B2(G128), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G29), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n744), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G2067), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n690), .A2(G5), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G171), .B2(new_n690), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(G1961), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n735), .A2(G2084), .A3(new_n739), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(G1961), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n756), .A2(new_n759), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT31), .B(G11), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT30), .B(G28), .Z(new_n764));
  OAI221_X1 g339(.A(new_n763), .B1(G29), .B2(new_n764), .C1(new_n626), .C2(new_n703), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n690), .A2(G4), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n607), .B2(new_n690), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G1348), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G168), .A2(new_n690), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n690), .B2(G21), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n772), .A2(new_n773), .B1(new_n767), .B2(G1348), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n690), .A2(G20), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT23), .Z(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G299), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1956), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n770), .A2(new_n774), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n742), .A2(new_n762), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n615), .A2(G127), .ZN(new_n782));
  NAND2_X1  g357(.A1(G115), .A2(G2104), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n480), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT25), .ZN(new_n787));
  NAND2_X1  g362(.A1(G103), .A2(G2104), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(G2105), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n480), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n474), .A2(G139), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n784), .B2(new_n785), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n786), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(KEYINPUT96), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n786), .B2(new_n792), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G33), .B(new_n797), .S(G29), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2072), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n753), .A2(G32), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT97), .B(KEYINPUT26), .Z(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n475), .A2(G105), .ZN(new_n805));
  AOI22_X1  g380(.A1(G129), .A2(new_n481), .B1(new_n474), .B2(G141), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n801), .B1(new_n807), .B2(new_n753), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT27), .ZN(new_n809));
  INV_X1    g384(.A(G1996), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n690), .A2(G19), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n546), .B2(new_n690), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G1341), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n703), .A2(G27), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT99), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G164), .B2(new_n703), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n814), .B1(G2078), .B2(new_n817), .ZN(new_n818));
  AOI211_X1 g393(.A(new_n811), .B(new_n818), .C1(G2078), .C2(new_n817), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n733), .A2(new_n781), .A3(new_n800), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n727), .A2(new_n820), .ZN(G311));
  INV_X1    g396(.A(G311), .ZN(G150));
  NAND2_X1  g397(.A1(new_n521), .A2(G67), .ZN(new_n823));
  NAND2_X1  g398(.A1(G80), .A2(G543), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n509), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT101), .B(G93), .Z(new_n826));
  INV_X1    g401(.A(G55), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n512), .A2(new_n826), .B1(new_n514), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT102), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n825), .A2(KEYINPUT102), .A3(new_n828), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G860), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT104), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n600), .A2(new_n608), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n838));
  XOR2_X1   g413(.A(new_n837), .B(new_n838), .Z(new_n839));
  INV_X1    g414(.A(new_n546), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n830), .B2(new_n831), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n823), .A2(new_n824), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n828), .B1(new_n842), .B2(G651), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n546), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n839), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n833), .B1(new_n847), .B2(KEYINPUT39), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n836), .B1(new_n848), .B2(new_n849), .ZN(G145));
  XNOR2_X1  g425(.A(new_n477), .B(new_n626), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(G162), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n797), .A2(KEYINPUT105), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n794), .A2(new_n854), .A3(new_n796), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n491), .A2(new_n493), .ZN(new_n856));
  INV_X1    g431(.A(new_n488), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n496), .A2(new_n497), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(new_n807), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n807), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n752), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n861), .B(new_n807), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n751), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n853), .A2(new_n855), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n474), .A2(G142), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n481), .A2(G130), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n480), .A2(G118), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT106), .Z(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(new_n617), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n617), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n874), .A2(new_n875), .A3(new_n702), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n702), .B1(new_n874), .B2(new_n875), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n866), .A2(new_n864), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(KEYINPUT105), .A3(new_n797), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n867), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n878), .B1(new_n867), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n852), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n867), .A2(new_n880), .ZN(new_n884));
  INV_X1    g459(.A(new_n878), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n852), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n867), .A2(new_n880), .A3(new_n878), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT107), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n883), .A2(new_n889), .A3(new_n893), .A4(new_n890), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n892), .A2(KEYINPUT40), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT40), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(G395));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n898));
  XNOR2_X1  g473(.A(G303), .B(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(new_n715), .ZN(new_n900));
  XNOR2_X1  g475(.A(G303), .B(KEYINPUT108), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(G305), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n692), .A2(G288), .ZN(new_n903));
  NOR2_X1   g478(.A1(G290), .A2(new_n710), .ZN(new_n904));
  OAI22_X1  g479(.A1(new_n900), .A2(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(G290), .B(G288), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(G305), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n899), .A2(new_n715), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT42), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n845), .B(new_n610), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n600), .A2(G299), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n595), .A2(new_n562), .A3(new_n556), .A4(new_n599), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n913), .A2(new_n918), .A3(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n916), .B1(new_n920), .B2(new_n912), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n911), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(G868), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(G868), .B2(new_n832), .ZN(G295));
  OAI21_X1  g499(.A(new_n923), .B1(G868), .B2(new_n832), .ZN(G331));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT113), .ZN(new_n927));
  NAND2_X1  g502(.A1(G171), .A2(new_n564), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT78), .B1(new_n533), .B2(new_n537), .ZN(new_n929));
  AOI21_X1  g504(.A(G286), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(G171), .A2(G168), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n841), .B(new_n844), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(G168), .B1(new_n566), .B2(new_n567), .ZN(new_n933));
  INV_X1    g508(.A(new_n931), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n843), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n546), .B1(new_n936), .B2(new_n829), .ZN(new_n937));
  INV_X1    g512(.A(new_n844), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n933), .B(new_n934), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n932), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n915), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n932), .A2(new_n939), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n919), .A2(KEYINPUT110), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n917), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n919), .A2(KEYINPUT110), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n915), .A2(KEYINPUT111), .A3(KEYINPUT41), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n944), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n942), .A2(KEYINPUT112), .B1(new_n943), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n915), .B1(new_n932), .B2(new_n939), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n910), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n920), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n910), .B(new_n942), .C1(new_n955), .C2(new_n940), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n890), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n927), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n905), .A2(new_n909), .ZN(new_n959));
  INV_X1    g534(.A(new_n949), .ZN(new_n960));
  OAI22_X1  g535(.A1(new_n960), .A2(new_n940), .B1(new_n951), .B2(new_n952), .ZN(new_n961));
  INV_X1    g536(.A(new_n953), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n940), .A2(new_n955), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(new_n951), .ZN(new_n965));
  AOI21_X1  g540(.A(G37), .B1(new_n965), .B2(new_n910), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n966), .A3(KEYINPUT113), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n926), .B1(new_n958), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n959), .B1(new_n964), .B2(new_n951), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT43), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT44), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n956), .A3(new_n890), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT109), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n972), .A2(new_n975), .A3(KEYINPUT43), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n963), .A2(new_n966), .A3(new_n926), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n971), .A2(new_n980), .ZN(G397));
  XNOR2_X1  g556(.A(KEYINPUT114), .B(G1384), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT45), .B1(new_n861), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n473), .A2(G40), .A3(new_n476), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(new_n810), .A3(new_n807), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT115), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n751), .B(new_n755), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n810), .B2(new_n807), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n986), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n702), .B(new_n706), .Z(new_n992));
  OAI211_X1 g567(.A(new_n988), .B(new_n991), .C1(new_n985), .C2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n692), .A2(new_n694), .ZN(new_n994));
  NAND2_X1  g569(.A1(G290), .A2(G1986), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n985), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n858), .B2(new_n860), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n984), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n999), .B(new_n1003), .C1(new_n494), .C2(new_n500), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n473), .A2(G40), .A3(new_n476), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1003), .B1(new_n494), .B2(new_n859), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1005), .B1(new_n1008), .B2(KEYINPUT117), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1002), .A2(new_n1009), .A3(new_n731), .ZN(new_n1010));
  OAI211_X1 g585(.A(KEYINPUT45), .B(new_n982), .C1(new_n494), .C2(new_n859), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1011), .A2(new_n984), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1003), .B1(new_n494), .B2(new_n500), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1971), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1010), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(G8), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G303), .A2(G8), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT55), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1022), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT118), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1976), .B1(new_n572), .B2(new_n574), .ZN(new_n1028));
  OR3_X1    g603(.A1(new_n1028), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT116), .B1(new_n1028), .B2(KEYINPUT52), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  OAI221_X1 g607(.A(G8), .B1(G288), .B2(new_n1032), .C1(new_n1007), .C2(new_n1006), .ZN(new_n1033));
  INV_X1    g608(.A(G1981), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n579), .A2(new_n1034), .A3(new_n582), .A4(new_n584), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1036));
  INV_X1    g611(.A(G48), .ZN(new_n1037));
  OAI22_X1  g612(.A1(new_n1036), .A2(new_n509), .B1(new_n1037), .B2(new_n514), .ZN(new_n1038));
  OAI21_X1  g613(.A(G1981), .B1(new_n1038), .B2(new_n583), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1035), .A2(KEYINPUT49), .A3(new_n1039), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n1007), .B2(new_n1006), .ZN(new_n1045));
  OAI22_X1  g620(.A1(new_n1031), .A2(new_n1033), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1033), .A2(KEYINPUT52), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n999), .B(new_n1003), .C1(new_n494), .C2(new_n859), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n984), .A3(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(G2090), .ZN(new_n1053));
  OAI211_X1 g628(.A(G8), .B(new_n1026), .C1(new_n1053), .C2(new_n1016), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT45), .B(new_n1003), .C1(new_n494), .C2(new_n500), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n984), .B(new_n1056), .C1(new_n998), .C2(KEYINPUT45), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n773), .ZN(new_n1058));
  INV_X1    g633(.A(G2084), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1050), .A2(new_n1059), .A3(new_n984), .A4(new_n1051), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1024), .B(G286), .C1(new_n1058), .C2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1023), .A2(new_n1027), .A3(new_n1055), .A4(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1061), .A2(KEYINPUT63), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1053), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1024), .B1(new_n1066), .B2(new_n1017), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1022), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1055), .B(new_n1065), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1064), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1058), .A2(G168), .A3(new_n1060), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1024), .B1(KEYINPUT125), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(KEYINPUT125), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(G8), .A3(G286), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1077), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1081), .A2(KEYINPUT62), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G2078), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1015), .A2(new_n1084), .A3(new_n984), .A4(new_n1011), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1052), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1006), .B1(new_n1007), .B2(new_n1014), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1086), .A2(G2078), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1091), .A3(new_n1056), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1087), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n602), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1083), .A2(new_n1094), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1023), .A2(new_n1027), .A3(new_n1055), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT62), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1032), .B(new_n710), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1045), .B1(new_n1099), .B2(new_n1035), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1054), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n1101), .B2(new_n1049), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1072), .A2(new_n1098), .A3(new_n1102), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1082), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n861), .A2(new_n982), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1012), .B(new_n1091), .C1(new_n1107), .C2(KEYINPUT45), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1108), .A2(new_n1087), .A3(G301), .A4(new_n1089), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1094), .A2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1104), .A2(new_n1105), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(new_n1020), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1108), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G171), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1116), .B(KEYINPUT54), .C1(new_n602), .C2(new_n1093), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1111), .A2(new_n1027), .A3(new_n1114), .A4(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(G1956), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1012), .A2(new_n1015), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT122), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G1956), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT117), .B(new_n984), .C1(new_n998), .C2(new_n999), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1004), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1008), .A2(KEYINPUT117), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n1121), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n562), .B2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(G299), .Z(new_n1133));
  NAND3_X1  g708(.A1(new_n1123), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1123), .A2(new_n1130), .A3(KEYINPUT123), .A4(new_n1133), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1052), .A2(new_n769), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1007), .A2(new_n1006), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n755), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n607), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1136), .A2(new_n1137), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1133), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1138), .A2(KEYINPUT60), .A3(new_n1140), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1148), .A2(KEYINPUT124), .A3(new_n600), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n600), .B1(new_n1148), .B2(KEYINPUT124), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1149), .A2(new_n1150), .B1(KEYINPUT124), .B2(new_n1148), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1141), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1144), .A2(new_n1155), .A3(new_n1145), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1155), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1146), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT58), .B(G1341), .ZN(new_n1160));
  OAI22_X1  g735(.A1(new_n1159), .A2(G1996), .B1(new_n1139), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n546), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT59), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1154), .A2(new_n1156), .A3(new_n1158), .A4(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1118), .B1(new_n1147), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n997), .B1(new_n1103), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n985), .B1(new_n807), .B2(new_n989), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT126), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n986), .A2(new_n810), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT46), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1171), .A2(KEYINPUT47), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(KEYINPUT47), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n985), .A2(new_n994), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT127), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT48), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1172), .A2(new_n1173), .B1(new_n1176), .B2(new_n993), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n702), .A2(new_n706), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n988), .A2(new_n1178), .A3(new_n991), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n752), .A2(new_n755), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n985), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1166), .A2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g758(.A1(G227), .A2(new_n459), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n688), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g760(.A(new_n1186), .B1(new_n647), .B2(new_n648), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n892), .A2(new_n894), .ZN(new_n1188));
  AND3_X1   g762(.A1(new_n1187), .A2(new_n1188), .A3(new_n978), .ZN(G308));
  NAND3_X1  g763(.A1(new_n1187), .A2(new_n1188), .A3(new_n978), .ZN(G225));
endmodule


