//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n192), .B1(new_n187), .B2(KEYINPUT16), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(KEYINPUT69), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n196), .B1(new_n200), .B2(G128), .ZN(new_n201));
  XOR2_X1   g015(.A(KEYINPUT24), .B(G110), .Z(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(KEYINPUT23), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT69), .B(G119), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(G110), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n189), .B(new_n194), .C1(new_n205), .C2(new_n211), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n193), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n194), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n201), .A2(new_n202), .ZN(new_n215));
  INV_X1    g029(.A(G110), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n206), .A2(new_n210), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G137), .ZN(new_n220));
  INV_X1    g034(.A(G221), .ZN(new_n221));
  INV_X1    g035(.A(G234), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n221), .A2(new_n222), .A3(G953), .ZN(new_n223));
  XOR2_X1   g037(.A(new_n220), .B(new_n223), .Z(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n212), .A2(new_n218), .A3(new_n224), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n229), .A2(new_n230), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G217), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(G234), .B2(new_n227), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n226), .A2(new_n228), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n235), .A2(G902), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(G472), .A2(G902), .ZN(new_n242));
  INV_X1    g056(.A(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT2), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G113), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G119), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n247), .B(new_n249), .C1(new_n207), .C2(new_n248), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT70), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n200), .A2(G116), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n252), .A2(new_n253), .A3(new_n247), .A4(new_n249), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n249), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n244), .A3(new_n246), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n188), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(G143), .B2(new_n188), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n262), .B1(new_n264), .B2(new_n209), .ZN(new_n265));
  XNOR2_X1  g079(.A(G143), .B(G146), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n263), .A3(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT71), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT11), .B1(new_n273), .B2(G137), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  INV_X1    g089(.A(G137), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(G134), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n274), .A2(new_n277), .B1(new_n273), .B2(G137), .ZN(new_n278));
  INV_X1    g092(.A(G131), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n281), .B1(new_n276), .B2(G134), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n276), .A2(G134), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n273), .A2(KEYINPUT66), .A3(G137), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G131), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT67), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n288), .A3(G131), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n272), .A2(new_n280), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n274), .A2(new_n277), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n273), .A2(G137), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G131), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n280), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT0), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n209), .ZN(new_n299));
  NAND2_X1  g113(.A1(KEYINPUT0), .A2(G128), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n262), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n266), .A2(new_n300), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n293), .A2(KEYINPUT65), .A3(G131), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n296), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n290), .A2(KEYINPUT30), .A3(new_n307), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n296), .A2(new_n305), .A3(new_n306), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n287), .A2(new_n310), .A3(new_n280), .A4(new_n289), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n311), .A2(new_n268), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n287), .A2(new_n280), .A3(new_n289), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT68), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n309), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n258), .B(new_n308), .C1(new_n315), .C2(KEYINPUT30), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT31), .ZN(new_n317));
  INV_X1    g131(.A(new_n258), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n290), .A2(new_n318), .A3(new_n307), .ZN(new_n319));
  NOR2_X1   g133(.A1(G237), .A2(G953), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G210), .ZN(new_n321));
  INV_X1    g135(.A(G101), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n323), .B(new_n324), .Z(new_n325));
  NAND4_X1  g139(.A1(new_n316), .A2(new_n317), .A3(new_n319), .A4(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n326), .A2(new_n327), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n316), .A2(new_n319), .A3(new_n325), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT31), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n319), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n315), .B2(new_n318), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n314), .A2(new_n268), .A3(new_n311), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n307), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT74), .A3(new_n258), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n319), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n334), .B1(new_n340), .B2(KEYINPUT28), .ZN(new_n341));
  XOR2_X1   g155(.A(new_n325), .B(KEYINPUT73), .Z(new_n342));
  OAI21_X1  g156(.A(new_n332), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n242), .B1(new_n330), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT32), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI221_X1 g160(.A(new_n332), .B1(new_n341), .B2(new_n342), .C1(new_n328), .C2(new_n329), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT32), .A3(new_n242), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n341), .A2(new_n342), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n341), .A2(KEYINPUT75), .A3(new_n342), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n316), .A2(new_n319), .ZN(new_n355));
  INV_X1    g169(.A(new_n325), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n352), .A2(new_n353), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n334), .A2(KEYINPUT77), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n313), .B1(new_n269), .B2(new_n271), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n258), .B1(new_n360), .B2(new_n309), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n319), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n290), .A2(new_n307), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(KEYINPUT76), .A3(new_n258), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(KEYINPUT28), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n363), .A2(KEYINPUT77), .A3(KEYINPUT28), .A4(new_n365), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT29), .A3(new_n325), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n227), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n358), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G472), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n241), .B1(new_n349), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G140), .ZN(new_n377));
  INV_X1    g191(.A(G227), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(G953), .ZN(new_n379));
  XOR2_X1   g193(.A(new_n377), .B(new_n379), .Z(new_n380));
  INV_X1    g194(.A(KEYINPUT12), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n296), .A2(new_n306), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT79), .B1(new_n384), .B2(G104), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(G107), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT3), .B1(new_n387), .B2(G107), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n384), .A3(G104), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n389), .A2(new_n322), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n390), .A2(new_n392), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n396), .A2(KEYINPUT80), .A3(new_n322), .A4(new_n389), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n384), .A2(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n387), .A2(G107), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n322), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n403));
  OAI21_X1  g217(.A(G128), .B1(new_n264), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n259), .A2(new_n403), .A3(KEYINPUT1), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n262), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n267), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n398), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n401), .B1(new_n395), .B2(new_n397), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(new_n268), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n381), .B(new_n383), .C1(new_n409), .C2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n398), .A2(new_n402), .A3(new_n408), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n410), .B2(new_n268), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n381), .B1(new_n415), .B2(new_n383), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n396), .A2(new_n389), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(G101), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n398), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT81), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n418), .A3(G101), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n398), .A2(new_n424), .A3(new_n420), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n422), .A2(new_n305), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT10), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(new_n269), .B2(new_n271), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n414), .A2(new_n427), .B1(new_n429), .B2(new_n410), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n430), .A3(new_n382), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n380), .B1(new_n417), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n426), .A2(new_n430), .A3(new_n382), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n382), .B1(new_n426), .B2(new_n430), .ZN(new_n434));
  INV_X1    g248(.A(new_n380), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n376), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n416), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n431), .A3(new_n412), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n435), .ZN(new_n440));
  INV_X1    g254(.A(new_n434), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n431), .A3(new_n380), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n442), .A3(KEYINPUT84), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(G469), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n417), .A2(new_n431), .A3(new_n380), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n435), .B1(new_n433), .B2(new_n434), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G469), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n227), .ZN(new_n449));
  NAND2_X1  g263(.A1(G469), .A2(G902), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT9), .B(G234), .Z(new_n452));
  AOI21_X1  g266(.A(new_n221), .B1(new_n452), .B2(new_n227), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G214), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(G952), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G953), .ZN(new_n459));
  INV_X1    g273(.A(G237), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n222), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G953), .ZN(new_n463));
  AOI211_X1 g277(.A(new_n227), .B(new_n463), .C1(G234), .C2(G237), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT21), .B(G898), .Z(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n470));
  XNOR2_X1  g284(.A(G110), .B(G122), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n471), .B(KEYINPUT8), .Z(new_n472));
  NAND2_X1  g286(.A1(new_n398), .A2(new_n402), .ZN(new_n473));
  OAI211_X1 g287(.A(KEYINPUT5), .B(new_n249), .C1(new_n207), .C2(new_n248), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(G113), .C1(KEYINPUT5), .C2(new_n252), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n255), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n410), .A2(new_n255), .A3(new_n475), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G125), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n303), .B2(new_n304), .ZN(new_n481));
  AOI21_X1  g295(.A(G125), .B1(new_n265), .B2(new_n267), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n463), .A2(G224), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n484), .A2(KEYINPUT7), .ZN(new_n485));
  OAI22_X1  g299(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n483), .B(new_n485), .C1(new_n481), .C2(new_n482), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n470), .B1(new_n479), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n472), .ZN(new_n492));
  AND4_X1   g306(.A1(new_n398), .A2(new_n255), .A3(new_n402), .A4(new_n475), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n398), .A2(new_n402), .B1(new_n255), .B2(new_n475), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n488), .A2(new_n489), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT88), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n422), .A2(new_n423), .A3(new_n425), .A4(new_n258), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n478), .A4(new_n471), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n478), .A3(new_n471), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT85), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n498), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n469), .B1(new_n504), .B2(G902), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n501), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n479), .A2(new_n470), .A3(new_n490), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT88), .B1(new_n495), .B2(new_n496), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT89), .A3(new_n227), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G210), .B1(G237), .B2(G902), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n471), .B1(new_n499), .B2(new_n478), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n514), .B1(new_n503), .B2(new_n501), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT6), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n481), .A2(new_n482), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n484), .B(KEYINPUT86), .Z(new_n520));
  XOR2_X1   g334(.A(new_n519), .B(new_n520), .Z(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n512), .A2(new_n513), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n513), .B1(new_n512), .B2(new_n522), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n457), .B(new_n468), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n320), .A2(G214), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n260), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n320), .A2(G143), .A3(G214), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G131), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n279), .A3(new_n529), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n531), .A2(new_n532), .B1(new_n193), .B2(G146), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n480), .A2(G140), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT19), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n191), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT90), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n187), .B2(new_n535), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n191), .A2(new_n534), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n538), .A2(new_n188), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n533), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n530), .ZN(new_n546));
  NAND2_X1  g360(.A1(KEYINPUT18), .A2(G131), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n541), .A2(G146), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n546), .A2(new_n547), .B1(new_n189), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n530), .A2(KEYINPUT18), .A3(G131), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G113), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n387), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(KEYINPUT92), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n533), .A2(new_n544), .B1(new_n549), .B2(new_n550), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(new_n554), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n531), .A2(new_n560), .A3(new_n532), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n530), .A2(KEYINPUT17), .A3(G131), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n561), .A2(new_n213), .A3(new_n194), .A4(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n554), .A3(new_n551), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n556), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT93), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT20), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G475), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n568), .A3(new_n227), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n567), .B(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n564), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n554), .B1(new_n563), .B2(new_n551), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n227), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(G475), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT95), .B1(new_n570), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT95), .ZN(new_n580));
  AND4_X1   g394(.A1(new_n568), .A2(new_n567), .A3(new_n227), .A4(new_n565), .ZN(new_n581));
  INV_X1    g395(.A(new_n565), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(G475), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n567), .B1(new_n583), .B2(new_n227), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n580), .B(new_n577), .C1(new_n581), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT99), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n587), .A2(KEYINPUT15), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(KEYINPUT15), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(G478), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n209), .A2(G143), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n260), .A2(G128), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n273), .ZN(new_n595));
  XNOR2_X1  g409(.A(G116), .B(G122), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n384), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n384), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n600), .A2(KEYINPUT97), .A3(new_n592), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT97), .B1(new_n600), .B2(new_n592), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n600), .A2(new_n592), .ZN(new_n603));
  NOR4_X1   g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n593), .ZN(new_n604));
  OAI221_X1 g418(.A(new_n595), .B1(new_n597), .B2(new_n599), .C1(new_n604), .C2(new_n273), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n599), .A2(KEYINPUT98), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n594), .B(new_n273), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n248), .A2(KEYINPUT14), .A3(G122), .ZN(new_n608));
  INV_X1    g422(.A(new_n596), .ZN(new_n609));
  OAI211_X1 g423(.A(G107), .B(new_n608), .C1(new_n609), .C2(KEYINPUT14), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n599), .A2(KEYINPUT98), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n606), .A2(new_n607), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n452), .A2(G217), .A3(new_n463), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n614), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n605), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n227), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n591), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n619), .B(new_n620), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n622), .B2(new_n591), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n586), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n375), .A2(new_n456), .A3(new_n526), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  AND3_X1   g441(.A1(new_n615), .A2(KEYINPUT33), .A3(new_n617), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT33), .B1(new_n615), .B2(new_n617), .ZN(new_n629));
  OAI21_X1  g443(.A(G478), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(G478), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n227), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n630), .B(new_n633), .C1(G478), .C2(new_n619), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n586), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT101), .B1(new_n525), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n347), .A2(new_n227), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(G472), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n344), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n640), .A2(new_n455), .A3(new_n241), .ZN(new_n641));
  INV_X1    g455(.A(new_n457), .ZN(new_n642));
  INV_X1    g456(.A(new_n513), .ZN(new_n643));
  AOI21_X1  g457(.A(KEYINPUT89), .B1(new_n510), .B2(new_n227), .ZN(new_n644));
  AOI211_X1 g458(.A(new_n469), .B(G902), .C1(new_n506), .C2(new_n509), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n518), .A2(new_n521), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n512), .A2(new_n513), .A3(new_n522), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n642), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n636), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n650), .A2(new_n651), .A3(new_n652), .A4(new_n468), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n637), .A2(new_n641), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  INV_X1    g470(.A(KEYINPUT20), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(KEYINPUT102), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n657), .A2(KEYINPUT102), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n569), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n569), .A2(new_n659), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n578), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n650), .A2(new_n468), .A3(new_n624), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n641), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NOR2_X1   g480(.A1(new_n640), .A2(new_n455), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n219), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n239), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT103), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n669), .A2(new_n672), .A3(new_n239), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n671), .B(new_n673), .C1(new_n233), .C2(new_n236), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n667), .A2(new_n526), .A3(new_n625), .A4(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n462), .B1(new_n464), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n662), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n623), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n650), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n451), .A2(new_n454), .A3(new_n674), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n346), .A2(new_n348), .ZN(new_n685));
  INV_X1    g499(.A(G472), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n358), .B2(new_n372), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n209), .ZN(G30));
  XOR2_X1   g504(.A(new_n679), .B(KEYINPUT39), .Z(new_n691));
  NAND2_X1  g505(.A1(new_n456), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n692), .A2(KEYINPUT40), .ZN(new_n693));
  INV_X1    g507(.A(new_n674), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(KEYINPUT40), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n693), .A2(new_n457), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n648), .A2(new_n649), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT38), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n623), .B1(new_n585), .B2(new_n579), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n331), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n363), .A2(new_n365), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n342), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n227), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G472), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n346), .A2(new_n348), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n696), .A2(new_n700), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n260), .ZN(G45));
  AOI211_X1 g523(.A(new_n679), .B(new_n634), .C1(new_n579), .C2(new_n585), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n697), .A3(new_n457), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n688), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n188), .ZN(G48));
  AND2_X1   g527(.A1(new_n354), .A2(new_n353), .ZN(new_n714));
  INV_X1    g528(.A(new_n357), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n350), .B2(new_n351), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n371), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n346), .B(new_n348), .C1(new_n717), .C2(new_n686), .ZN(new_n718));
  INV_X1    g532(.A(new_n449), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n448), .B1(new_n447), .B2(new_n227), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n719), .A2(new_n453), .A3(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n718), .A2(new_n240), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n637), .A3(new_n653), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NAND2_X1  g539(.A1(new_n663), .A2(new_n722), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  OAI211_X1 g541(.A(new_n721), .B(new_n457), .C1(new_n523), .C2(new_n524), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n697), .A2(KEYINPUT104), .A3(new_n457), .A4(new_n721), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n718), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n467), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n586), .A2(new_n624), .A3(new_n694), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT105), .B(G119), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G21));
  OAI221_X1 g552(.A(new_n332), .B1(new_n369), .B2(new_n342), .C1(new_n328), .C2(new_n329), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n638), .A2(G472), .B1(new_n242), .B2(new_n739), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(new_n240), .A3(new_n721), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n526), .A3(new_n699), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NAND3_X1  g557(.A1(new_n740), .A2(new_n710), .A3(new_n674), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n730), .B2(new_n731), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n480), .ZN(G27));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n432), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n440), .A2(KEYINPUT107), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n749), .A3(G469), .A4(new_n442), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n450), .B(KEYINPUT106), .Z(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n449), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n453), .A2(new_n642), .ZN(new_n753));
  AND4_X1   g567(.A1(new_n648), .A2(new_n649), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n718), .A3(new_n240), .A4(new_n710), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n375), .A2(KEYINPUT42), .A3(new_n710), .A4(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  NAND3_X1  g574(.A1(new_n375), .A2(new_n682), .A3(new_n754), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NAND3_X1  g576(.A1(new_n579), .A2(new_n585), .A3(new_n635), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT43), .Z(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n640), .A3(new_n674), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n697), .A2(new_n642), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n764), .A2(KEYINPUT44), .A3(new_n640), .A4(new_n674), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n448), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n444), .A2(KEYINPUT108), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT108), .B1(new_n444), .B2(new_n774), .ZN(new_n776));
  AND4_X1   g590(.A1(KEYINPUT45), .A2(new_n749), .A3(new_n442), .A4(new_n748), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT46), .ZN(new_n779));
  INV_X1    g593(.A(new_n751), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n449), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n454), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT109), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n767), .A2(new_n786), .A3(new_n768), .A4(new_n769), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n771), .A2(new_n691), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  NAND2_X1  g603(.A1(new_n784), .A2(KEYINPUT47), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n783), .A2(new_n791), .A3(new_n454), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n790), .A2(new_n710), .A3(new_n768), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n733), .A2(new_n241), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  INV_X1    g610(.A(new_n698), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n706), .A2(new_n241), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n719), .A2(new_n720), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n753), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI211_X1 g615(.A(new_n763), .B(new_n801), .C1(new_n800), .C2(new_n799), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n797), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  INV_X1    g618(.A(new_n768), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n790), .A2(new_n792), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n799), .A2(new_n453), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n764), .A2(new_n462), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT114), .Z(new_n810));
  AND3_X1   g624(.A1(new_n810), .A2(new_n240), .A3(new_n740), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n804), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n810), .A2(new_n642), .A3(new_n797), .A4(new_n741), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n740), .A2(new_n674), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n523), .A2(new_n524), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n799), .A3(new_n753), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT115), .Z(new_n823));
  AND2_X1   g637(.A1(new_n810), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n808), .A2(new_n811), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n462), .A3(new_n798), .ZN(new_n826));
  OR3_X1    g640(.A1(new_n826), .A2(new_n586), .A3(new_n635), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n818), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n815), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n814), .A2(new_n827), .A3(new_n818), .A4(new_n825), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n826), .A2(new_n636), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n829), .A2(new_n830), .A3(new_n459), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n744), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n754), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n624), .A2(new_n681), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n821), .A2(new_n457), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT110), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT110), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n768), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n451), .A2(new_n454), .A3(new_n674), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n349), .B2(new_n374), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n837), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n759), .A2(new_n761), .A3(new_n834), .A4(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n736), .A2(new_n723), .A3(new_n726), .A4(new_n742), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n625), .B1(new_n586), .B2(new_n634), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n641), .A2(new_n526), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n626), .A2(new_n846), .A3(new_n675), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n688), .B1(new_n683), .B2(new_n711), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n745), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n679), .A2(new_n453), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n706), .A2(new_n694), .A3(new_n752), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n697), .A2(new_n457), .A3(new_n699), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n849), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n745), .A2(new_n850), .A3(new_n855), .A4(KEYINPUT52), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT112), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n732), .A2(new_n833), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n841), .B(new_n650), .C1(new_n682), .C2(new_n710), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n856), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT52), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n851), .A2(new_n849), .A3(new_n856), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT112), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n848), .A2(new_n859), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n863), .A2(new_n864), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n868), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n848), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT113), .B1(new_n873), .B2(KEYINPUT54), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n870), .B1(new_n848), .B2(KEYINPUT111), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT111), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n844), .A2(new_n847), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n878), .B2(new_n843), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT53), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n867), .A2(new_n868), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT54), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n811), .A2(new_n732), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n867), .A2(new_n868), .B1(new_n848), .B2(new_n871), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT113), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n874), .A2(new_n882), .A3(new_n883), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n824), .A2(new_n375), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT48), .Z(new_n890));
  NOR3_X1   g704(.A1(new_n832), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(G952), .A2(G953), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n803), .B1(new_n891), .B2(new_n892), .ZN(G75));
  NOR2_X1   g707(.A1(new_n884), .A2(new_n227), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT56), .B1(new_n894), .B2(G210), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n518), .B(new_n521), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT55), .Z(new_n897));
  AND2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n895), .A2(new_n897), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n458), .A2(G953), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT117), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(G51));
  XNOR2_X1  g717(.A(new_n884), .B(new_n886), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n751), .B(KEYINPUT57), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n447), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n894), .A2(new_n778), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n902), .B1(new_n907), .B2(new_n908), .ZN(G54));
  INV_X1    g723(.A(KEYINPUT58), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT118), .B1(new_n910), .B2(new_n568), .ZN(new_n911));
  OR3_X1    g725(.A1(new_n910), .A2(new_n568), .A3(KEYINPUT118), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n894), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n582), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n902), .ZN(G60));
  OR2_X1    g729(.A1(new_n628), .A2(new_n629), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n632), .B(KEYINPUT59), .Z(new_n918));
  AND2_X1   g732(.A1(new_n884), .A2(new_n886), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n884), .A2(new_n886), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n917), .B(new_n918), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n904), .A2(KEYINPUT119), .A3(new_n917), .A4(new_n918), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n874), .A2(new_n882), .A3(new_n887), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n918), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n916), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n925), .A2(new_n928), .A3(new_n901), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT60), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n873), .A2(new_n669), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT121), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n873), .A2(new_n935), .A3(new_n669), .A4(new_n932), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n238), .B(KEYINPUT122), .Z(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n884), .B2(new_n931), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n934), .A2(new_n901), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT61), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT61), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(G66));
  INV_X1    g757(.A(G224), .ZN(new_n944));
  OAI21_X1  g758(.A(G953), .B1(new_n466), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n877), .B2(G953), .ZN(new_n946));
  INV_X1    g760(.A(new_n518), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(G898), .B2(new_n463), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(G69));
  OAI21_X1  g763(.A(G953), .B1(new_n378), .B2(new_n678), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n678), .A2(G953), .ZN(new_n952));
  MUX2_X1   g766(.A(new_n315), .B(new_n364), .S(KEYINPUT30), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n538), .A2(new_n543), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT123), .Z(new_n955));
  XOR2_X1   g769(.A(new_n953), .B(new_n955), .Z(new_n956));
  OAI21_X1  g770(.A(new_n788), .B1(new_n793), .B2(new_n794), .ZN(new_n957));
  INV_X1    g771(.A(new_n375), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(new_n854), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n785), .A2(new_n691), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n851), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n759), .A2(new_n761), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT125), .Z(new_n963));
  NOR3_X1   g777(.A1(new_n957), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n952), .B(new_n956), .C1(new_n964), .C2(G953), .ZN(new_n965));
  INV_X1    g779(.A(new_n956), .ZN(new_n966));
  INV_X1    g780(.A(new_n845), .ZN(new_n967));
  NOR4_X1   g781(.A1(new_n958), .A2(new_n967), .A3(new_n805), .A4(new_n692), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n708), .ZN(new_n970));
  XOR2_X1   g784(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n851), .A3(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n795), .A2(new_n788), .A3(new_n969), .A4(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT62), .ZN(new_n974));
  AOI22_X1  g788(.A1(new_n970), .A2(new_n851), .B1(KEYINPUT124), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n463), .B(new_n966), .C1(new_n973), .C2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n965), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n977), .B1(new_n965), .B2(new_n976), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n951), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n980), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n982), .A2(new_n950), .A3(new_n978), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n983), .ZN(G72));
  OAI211_X1 g798(.A(new_n788), .B(new_n972), .C1(new_n793), .C2(new_n794), .ZN(new_n985));
  NOR4_X1   g799(.A1(new_n985), .A2(new_n975), .A3(new_n878), .A4(new_n968), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OR3_X1    g804(.A1(new_n986), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n987), .B1(new_n986), .B2(new_n990), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n991), .A2(new_n325), .A3(new_n355), .A4(new_n992), .ZN(new_n993));
  OAI221_X1 g807(.A(new_n989), .B1(new_n715), .B2(new_n701), .C1(new_n880), .C2(new_n881), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n964), .A2(new_n877), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n355), .B1(new_n995), .B2(new_n989), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n902), .B1(new_n996), .B2(new_n356), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n993), .A2(new_n994), .A3(new_n997), .ZN(G57));
endmodule


