

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(n670), .A2(n845), .ZN(n618) );
  INV_X1 U558 ( .A(KEYINPUT29), .ZN(n650) );
  XNOR2_X1 U559 ( .A(n651), .B(n650), .ZN(n652) );
  OR2_X2 U560 ( .A1(n710), .A2(n602), .ZN(n670) );
  AND2_X1 U561 ( .A1(G2104), .A2(n545), .ZN(n540) );
  XNOR2_X1 U562 ( .A(n540), .B(KEYINPUT64), .ZN(n690) );
  NOR2_X1 U563 ( .A1(G651), .A2(n557), .ZN(n792) );
  XNOR2_X1 U564 ( .A(n758), .B(KEYINPUT40), .ZN(n759) );
  XNOR2_X1 U565 ( .A(n760), .B(n759), .ZN(G329) );
  XOR2_X1 U566 ( .A(KEYINPUT4), .B(KEYINPUT70), .Z(n526) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n795) );
  NAND2_X1 U568 ( .A1(G89), .A2(n795), .ZN(n525) );
  XNOR2_X1 U569 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U570 ( .A(KEYINPUT69), .B(n527), .ZN(n529) );
  XOR2_X1 U571 ( .A(G543), .B(KEYINPUT0), .Z(n557) );
  INV_X1 U572 ( .A(G651), .ZN(n531) );
  NOR2_X1 U573 ( .A1(n557), .A2(n531), .ZN(n791) );
  NAND2_X1 U574 ( .A1(n791), .A2(G76), .ZN(n528) );
  NAND2_X1 U575 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U576 ( .A(n530), .B(KEYINPUT5), .ZN(n538) );
  NOR2_X1 U577 ( .A1(G543), .A2(n531), .ZN(n532) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n532), .Z(n533) );
  BUF_X1 U579 ( .A(n533), .Z(n796) );
  NAND2_X1 U580 ( .A1(G63), .A2(n796), .ZN(n535) );
  NAND2_X1 U581 ( .A1(G51), .A2(n792), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U583 ( .A(KEYINPUT6), .B(n536), .Z(n537) );
  NAND2_X1 U584 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U585 ( .A(n539), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U586 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U588 ( .A1(n885), .A2(G113), .ZN(n543) );
  INV_X1 U589 ( .A(G2105), .ZN(n545) );
  NAND2_X1 U590 ( .A1(n690), .A2(G101), .ZN(n541) );
  XOR2_X1 U591 ( .A(KEYINPUT23), .B(n541), .Z(n542) );
  NAND2_X1 U592 ( .A1(n543), .A2(n542), .ZN(n549) );
  NOR2_X1 U593 ( .A1(G2105), .A2(G2104), .ZN(n544) );
  XOR2_X1 U594 ( .A(KEYINPUT17), .B(n544), .Z(n695) );
  NAND2_X1 U595 ( .A1(G137), .A2(n695), .ZN(n547) );
  NOR2_X1 U596 ( .A1(G2104), .A2(n545), .ZN(n886) );
  NAND2_X1 U597 ( .A1(G125), .A2(n886), .ZN(n546) );
  NAND2_X1 U598 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U599 ( .A1(n549), .A2(n548), .ZN(G160) );
  NAND2_X1 U600 ( .A1(G114), .A2(n885), .ZN(n551) );
  NAND2_X1 U601 ( .A1(G126), .A2(n886), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n551), .A2(n550), .ZN(n556) );
  NAND2_X1 U603 ( .A1(G102), .A2(n690), .ZN(n552) );
  XNOR2_X1 U604 ( .A(n552), .B(KEYINPUT90), .ZN(n554) );
  NAND2_X1 U605 ( .A1(G138), .A2(n695), .ZN(n553) );
  NAND2_X1 U606 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U607 ( .A1(n556), .A2(n555), .ZN(G164) );
  NAND2_X1 U608 ( .A1(G87), .A2(n557), .ZN(n558) );
  XNOR2_X1 U609 ( .A(n558), .B(KEYINPUT76), .ZN(n563) );
  NAND2_X1 U610 ( .A1(G49), .A2(n792), .ZN(n560) );
  NAND2_X1 U611 ( .A1(G74), .A2(G651), .ZN(n559) );
  NAND2_X1 U612 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U613 ( .A1(n796), .A2(n561), .ZN(n562) );
  NAND2_X1 U614 ( .A1(n563), .A2(n562), .ZN(G288) );
  NAND2_X1 U615 ( .A1(G75), .A2(n791), .ZN(n564) );
  XNOR2_X1 U616 ( .A(n564), .B(KEYINPUT80), .ZN(n571) );
  NAND2_X1 U617 ( .A1(G88), .A2(n795), .ZN(n566) );
  NAND2_X1 U618 ( .A1(G50), .A2(n792), .ZN(n565) );
  NAND2_X1 U619 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U620 ( .A1(G62), .A2(n796), .ZN(n567) );
  XNOR2_X1 U621 ( .A(KEYINPUT79), .B(n567), .ZN(n568) );
  NOR2_X1 U622 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U623 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U624 ( .A(KEYINPUT81), .B(n572), .ZN(G166) );
  INV_X1 U625 ( .A(G166), .ZN(G303) );
  NAND2_X1 U626 ( .A1(G64), .A2(n796), .ZN(n574) );
  NAND2_X1 U627 ( .A1(G52), .A2(n792), .ZN(n573) );
  NAND2_X1 U628 ( .A1(n574), .A2(n573), .ZN(n579) );
  NAND2_X1 U629 ( .A1(G90), .A2(n795), .ZN(n576) );
  NAND2_X1 U630 ( .A1(G77), .A2(n791), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U632 ( .A(KEYINPUT9), .B(n577), .Z(n578) );
  NOR2_X1 U633 ( .A1(n579), .A2(n578), .ZN(G171) );
  NAND2_X1 U634 ( .A1(G91), .A2(n795), .ZN(n581) );
  NAND2_X1 U635 ( .A1(G65), .A2(n796), .ZN(n580) );
  NAND2_X1 U636 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U637 ( .A1(G53), .A2(n792), .ZN(n582) );
  XNOR2_X1 U638 ( .A(KEYINPUT65), .B(n582), .ZN(n583) );
  NOR2_X1 U639 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U640 ( .A1(n791), .A2(G78), .ZN(n585) );
  NAND2_X1 U641 ( .A1(n586), .A2(n585), .ZN(G299) );
  NAND2_X1 U642 ( .A1(n791), .A2(G73), .ZN(n588) );
  XNOR2_X1 U643 ( .A(KEYINPUT78), .B(KEYINPUT2), .ZN(n587) );
  XNOR2_X1 U644 ( .A(n588), .B(n587), .ZN(n595) );
  NAND2_X1 U645 ( .A1(G86), .A2(n795), .ZN(n590) );
  NAND2_X1 U646 ( .A1(G48), .A2(n792), .ZN(n589) );
  NAND2_X1 U647 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U648 ( .A1(G61), .A2(n796), .ZN(n591) );
  XNOR2_X1 U649 ( .A(KEYINPUT77), .B(n591), .ZN(n592) );
  NOR2_X1 U650 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U651 ( .A1(n595), .A2(n594), .ZN(G305) );
  NAND2_X1 U652 ( .A1(G85), .A2(n795), .ZN(n597) );
  NAND2_X1 U653 ( .A1(G60), .A2(n796), .ZN(n596) );
  NAND2_X1 U654 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U655 ( .A1(G72), .A2(n791), .ZN(n599) );
  NAND2_X1 U656 ( .A1(G47), .A2(n792), .ZN(n598) );
  NAND2_X1 U657 ( .A1(n599), .A2(n598), .ZN(n600) );
  OR2_X1 U658 ( .A1(n601), .A2(n600), .ZN(G290) );
  NAND2_X1 U659 ( .A1(G160), .A2(G40), .ZN(n710) );
  NOR2_X1 U660 ( .A1(G164), .A2(G1384), .ZN(n711) );
  INV_X1 U661 ( .A(n711), .ZN(n602) );
  NAND2_X1 U662 ( .A1(G8), .A2(n670), .ZN(n735) );
  NOR2_X1 U663 ( .A1(G1976), .A2(G288), .ZN(n606) );
  NAND2_X1 U664 ( .A1(n606), .A2(KEYINPUT33), .ZN(n603) );
  NOR2_X1 U665 ( .A1(n735), .A2(n603), .ZN(n604) );
  XOR2_X1 U666 ( .A(KEYINPUT103), .B(n604), .Z(n688) );
  NOR2_X1 U667 ( .A1(G1971), .A2(G303), .ZN(n605) );
  NOR2_X1 U668 ( .A1(n606), .A2(n605), .ZN(n989) );
  NOR2_X1 U669 ( .A1(G2084), .A2(n670), .ZN(n655) );
  NAND2_X1 U670 ( .A1(G8), .A2(n655), .ZN(n668) );
  NOR2_X1 U671 ( .A1(G1966), .A2(n735), .ZN(n666) );
  XNOR2_X1 U672 ( .A(G2078), .B(KEYINPUT25), .ZN(n954) );
  NOR2_X1 U673 ( .A1(n670), .A2(n954), .ZN(n608) );
  AND2_X1 U674 ( .A1(n670), .A2(G1961), .ZN(n607) );
  NOR2_X1 U675 ( .A1(n608), .A2(n607), .ZN(n654) );
  NAND2_X1 U676 ( .A1(G171), .A2(n654), .ZN(n653) );
  NAND2_X1 U677 ( .A1(G56), .A2(n796), .ZN(n609) );
  XOR2_X1 U678 ( .A(KEYINPUT14), .B(n609), .Z(n615) );
  NAND2_X1 U679 ( .A1(n795), .A2(G81), .ZN(n610) );
  XNOR2_X1 U680 ( .A(n610), .B(KEYINPUT12), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G68), .A2(n791), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U683 ( .A(KEYINPUT13), .B(n613), .Z(n614) );
  NOR2_X1 U684 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U685 ( .A1(n792), .A2(G43), .ZN(n616) );
  NAND2_X1 U686 ( .A1(n617), .A2(n616), .ZN(n991) );
  INV_X1 U687 ( .A(G1996), .ZN(n845) );
  XOR2_X1 U688 ( .A(n618), .B(KEYINPUT26), .Z(n620) );
  NAND2_X1 U689 ( .A1(n670), .A2(G1341), .ZN(n619) );
  NAND2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U691 ( .A1(n991), .A2(n621), .ZN(n636) );
  NAND2_X1 U692 ( .A1(n796), .A2(G66), .ZN(n622) );
  XOR2_X1 U693 ( .A(KEYINPUT67), .B(n622), .Z(n624) );
  NAND2_X1 U694 ( .A1(n795), .A2(G92), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U696 ( .A(KEYINPUT68), .B(n625), .ZN(n629) );
  NAND2_X1 U697 ( .A1(G79), .A2(n791), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G54), .A2(n792), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U701 ( .A(KEYINPUT15), .B(n630), .Z(n977) );
  NAND2_X1 U702 ( .A1(n636), .A2(n977), .ZN(n634) );
  NOR2_X1 U703 ( .A1(G2067), .A2(n670), .ZN(n632) );
  INV_X1 U704 ( .A(n670), .ZN(n639) );
  NOR2_X1 U705 ( .A1(n639), .A2(G1348), .ZN(n631) );
  NOR2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n635), .B(KEYINPUT98), .ZN(n638) );
  OR2_X1 U709 ( .A1(n636), .A2(n977), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n645) );
  INV_X1 U711 ( .A(G299), .ZN(n978) );
  NAND2_X1 U712 ( .A1(n670), .A2(G1956), .ZN(n642) );
  NAND2_X1 U713 ( .A1(n639), .A2(G2072), .ZN(n640) );
  XOR2_X1 U714 ( .A(KEYINPUT27), .B(n640), .Z(n641) );
  NAND2_X1 U715 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(KEYINPUT97), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n978), .A2(n646), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n649) );
  NOR2_X1 U719 ( .A1(n978), .A2(n646), .ZN(n647) );
  XOR2_X1 U720 ( .A(n647), .B(KEYINPUT28), .Z(n648) );
  NAND2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n653), .A2(n652), .ZN(n664) );
  NOR2_X1 U723 ( .A1(G171), .A2(n654), .ZN(n661) );
  NOR2_X1 U724 ( .A1(n666), .A2(n655), .ZN(n656) );
  XOR2_X1 U725 ( .A(KEYINPUT99), .B(n656), .Z(n657) );
  NAND2_X1 U726 ( .A1(G8), .A2(n657), .ZN(n658) );
  XNOR2_X1 U727 ( .A(KEYINPUT30), .B(n658), .ZN(n659) );
  NOR2_X1 U728 ( .A1(G168), .A2(n659), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT31), .B(n662), .Z(n663) );
  NAND2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n669) );
  INV_X1 U732 ( .A(n669), .ZN(n665) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n680) );
  NAND2_X1 U735 ( .A1(n669), .A2(G286), .ZN(n676) );
  NOR2_X1 U736 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n671), .B(KEYINPUT100), .ZN(n673) );
  NOR2_X1 U738 ( .A1(n735), .A2(G1971), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U740 ( .A1(n674), .A2(G303), .ZN(n675) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U742 ( .A1(G8), .A2(n677), .ZN(n678) );
  XNOR2_X1 U743 ( .A(n678), .B(KEYINPUT32), .ZN(n679) );
  NAND2_X1 U744 ( .A1(n680), .A2(n679), .ZN(n731) );
  NAND2_X1 U745 ( .A1(n989), .A2(n731), .ZN(n681) );
  XNOR2_X1 U746 ( .A(KEYINPUT101), .B(n681), .ZN(n684) );
  NAND2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n981) );
  INV_X1 U748 ( .A(n735), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n981), .A2(n682), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n685), .A2(KEYINPUT33), .ZN(n686) );
  XNOR2_X1 U752 ( .A(n686), .B(KEYINPUT102), .ZN(n687) );
  NOR2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n728) );
  XOR2_X1 U754 ( .A(G1981), .B(G305), .Z(n992) );
  XNOR2_X1 U755 ( .A(KEYINPUT91), .B(G1986), .ZN(n689) );
  XNOR2_X1 U756 ( .A(n689), .B(G290), .ZN(n975) );
  INV_X1 U757 ( .A(n690), .ZN(n691) );
  INV_X1 U758 ( .A(n691), .ZN(n890) );
  NAND2_X1 U759 ( .A1(G95), .A2(n890), .ZN(n694) );
  NAND2_X1 U760 ( .A1(G107), .A2(n885), .ZN(n692) );
  XOR2_X1 U761 ( .A(KEYINPUT95), .B(n692), .Z(n693) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n699) );
  BUF_X1 U763 ( .A(n695), .Z(n889) );
  NAND2_X1 U764 ( .A1(G131), .A2(n889), .ZN(n697) );
  NAND2_X1 U765 ( .A1(G119), .A2(n886), .ZN(n696) );
  NAND2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n882) );
  INV_X1 U768 ( .A(G1991), .ZN(n844) );
  NOR2_X1 U769 ( .A1(n882), .A2(n844), .ZN(n709) );
  NAND2_X1 U770 ( .A1(G117), .A2(n885), .ZN(n701) );
  NAND2_X1 U771 ( .A1(G129), .A2(n886), .ZN(n700) );
  NAND2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U773 ( .A1(n890), .A2(G105), .ZN(n702) );
  XOR2_X1 U774 ( .A(KEYINPUT38), .B(n702), .Z(n703) );
  NOR2_X1 U775 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U776 ( .A1(n889), .A2(G141), .ZN(n705) );
  NAND2_X1 U777 ( .A1(n706), .A2(n705), .ZN(n866) );
  NAND2_X1 U778 ( .A1(G1996), .A2(n866), .ZN(n707) );
  XOR2_X1 U779 ( .A(KEYINPUT96), .B(n707), .Z(n708) );
  NOR2_X1 U780 ( .A1(n709), .A2(n708), .ZN(n935) );
  NAND2_X1 U781 ( .A1(n975), .A2(n935), .ZN(n712) );
  NOR2_X1 U782 ( .A1(n711), .A2(n710), .ZN(n752) );
  NAND2_X1 U783 ( .A1(n712), .A2(n752), .ZN(n725) );
  NAND2_X1 U784 ( .A1(n889), .A2(G140), .ZN(n713) );
  XNOR2_X1 U785 ( .A(KEYINPUT93), .B(n713), .ZN(n716) );
  NAND2_X1 U786 ( .A1(G104), .A2(n890), .ZN(n714) );
  XOR2_X1 U787 ( .A(KEYINPUT92), .B(n714), .Z(n715) );
  NOR2_X1 U788 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U789 ( .A(KEYINPUT34), .B(n717), .ZN(n722) );
  NAND2_X1 U790 ( .A1(G116), .A2(n885), .ZN(n719) );
  NAND2_X1 U791 ( .A1(G128), .A2(n886), .ZN(n718) );
  NAND2_X1 U792 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U793 ( .A(KEYINPUT35), .B(n720), .ZN(n721) );
  NAND2_X1 U794 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U795 ( .A(n723), .B(KEYINPUT36), .ZN(n724) );
  XOR2_X1 U796 ( .A(KEYINPUT94), .B(n724), .Z(n898) );
  XNOR2_X1 U797 ( .A(G2067), .B(KEYINPUT37), .ZN(n740) );
  NOR2_X1 U798 ( .A1(n898), .A2(n740), .ZN(n937) );
  NAND2_X1 U799 ( .A1(n937), .A2(n752), .ZN(n747) );
  NAND2_X1 U800 ( .A1(n725), .A2(n747), .ZN(n739) );
  INV_X1 U801 ( .A(n739), .ZN(n726) );
  AND2_X1 U802 ( .A1(n992), .A2(n726), .ZN(n727) );
  NAND2_X1 U803 ( .A1(n728), .A2(n727), .ZN(n757) );
  NOR2_X1 U804 ( .A1(G2090), .A2(G303), .ZN(n729) );
  NAND2_X1 U805 ( .A1(G8), .A2(n729), .ZN(n730) );
  NAND2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n732) );
  AND2_X1 U807 ( .A1(n732), .A2(n735), .ZN(n737) );
  NOR2_X1 U808 ( .A1(G1981), .A2(G305), .ZN(n733) );
  XOR2_X1 U809 ( .A(n733), .B(KEYINPUT24), .Z(n734) );
  NOR2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U811 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U812 ( .A1(n739), .A2(n738), .ZN(n755) );
  NAND2_X1 U813 ( .A1(n898), .A2(n740), .ZN(n939) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n866), .ZN(n929) );
  INV_X1 U815 ( .A(n935), .ZN(n743) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n741) );
  AND2_X1 U817 ( .A1(n844), .A2(n882), .ZN(n925) );
  NOR2_X1 U818 ( .A1(n741), .A2(n925), .ZN(n742) );
  NOR2_X1 U819 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U820 ( .A1(n929), .A2(n744), .ZN(n745) );
  XNOR2_X1 U821 ( .A(KEYINPUT39), .B(n745), .ZN(n746) );
  XNOR2_X1 U822 ( .A(n746), .B(KEYINPUT104), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n939), .A2(n749), .ZN(n750) );
  XOR2_X1 U825 ( .A(KEYINPUT105), .B(n750), .Z(n751) );
  NAND2_X1 U826 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U827 ( .A(KEYINPUT106), .B(n753), .Z(n754) );
  NOR2_X1 U828 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U829 ( .A1(n757), .A2(n756), .ZN(n760) );
  INV_X1 U830 ( .A(KEYINPUT107), .ZN(n758) );
  INV_X1 U831 ( .A(G96), .ZN(G221) );
  AND2_X1 U832 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U833 ( .A1(G123), .A2(n886), .ZN(n761) );
  XOR2_X1 U834 ( .A(KEYINPUT18), .B(n761), .Z(n767) );
  NAND2_X1 U835 ( .A1(n885), .A2(G111), .ZN(n762) );
  XNOR2_X1 U836 ( .A(n762), .B(KEYINPUT72), .ZN(n764) );
  NAND2_X1 U837 ( .A1(G99), .A2(n890), .ZN(n763) );
  NAND2_X1 U838 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U839 ( .A(KEYINPUT73), .B(n765), .Z(n766) );
  NOR2_X1 U840 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U841 ( .A1(n889), .A2(G135), .ZN(n768) );
  NAND2_X1 U842 ( .A1(n769), .A2(n768), .ZN(n926) );
  XNOR2_X1 U843 ( .A(G2096), .B(n926), .ZN(n770) );
  OR2_X1 U844 ( .A1(G2100), .A2(n770), .ZN(G156) );
  INV_X1 U845 ( .A(G120), .ZN(G236) );
  INV_X1 U846 ( .A(G69), .ZN(G235) );
  INV_X1 U847 ( .A(G108), .ZN(G238) );
  INV_X1 U848 ( .A(G171), .ZN(G301) );
  NAND2_X1 U849 ( .A1(G7), .A2(G661), .ZN(n771) );
  XOR2_X1 U850 ( .A(n771), .B(KEYINPUT10), .Z(n923) );
  NAND2_X1 U851 ( .A1(n923), .A2(G567), .ZN(n772) );
  XOR2_X1 U852 ( .A(KEYINPUT11), .B(n772), .Z(G234) );
  INV_X1 U853 ( .A(G860), .ZN(n779) );
  NOR2_X1 U854 ( .A1(n991), .A2(n779), .ZN(n773) );
  XOR2_X1 U855 ( .A(KEYINPUT66), .B(n773), .Z(G153) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n775) );
  OR2_X1 U857 ( .A1(n977), .A2(G868), .ZN(n774) );
  NAND2_X1 U858 ( .A1(n775), .A2(n774), .ZN(G284) );
  INV_X1 U859 ( .A(G868), .ZN(n806) );
  NAND2_X1 U860 ( .A1(n978), .A2(n806), .ZN(n776) );
  XNOR2_X1 U861 ( .A(n776), .B(KEYINPUT71), .ZN(n778) );
  NOR2_X1 U862 ( .A1(n806), .A2(G286), .ZN(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n779), .A2(G559), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n780), .A2(n977), .ZN(n781) );
  XNOR2_X1 U866 ( .A(n781), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U867 ( .A1(G868), .A2(n991), .ZN(n784) );
  NAND2_X1 U868 ( .A1(n977), .A2(G868), .ZN(n782) );
  NOR2_X1 U869 ( .A1(G559), .A2(n782), .ZN(n783) );
  NOR2_X1 U870 ( .A1(n784), .A2(n783), .ZN(G282) );
  XNOR2_X1 U871 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n786) );
  XNOR2_X1 U872 ( .A(G288), .B(KEYINPUT82), .ZN(n785) );
  XNOR2_X1 U873 ( .A(n786), .B(n785), .ZN(n787) );
  XNOR2_X1 U874 ( .A(G290), .B(n787), .ZN(n789) );
  XOR2_X1 U875 ( .A(G299), .B(G166), .Z(n788) );
  XNOR2_X1 U876 ( .A(n789), .B(n788), .ZN(n790) );
  XNOR2_X1 U877 ( .A(n790), .B(G305), .ZN(n802) );
  NAND2_X1 U878 ( .A1(G80), .A2(n791), .ZN(n794) );
  NAND2_X1 U879 ( .A1(G55), .A2(n792), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n800) );
  NAND2_X1 U881 ( .A1(G93), .A2(n795), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G67), .A2(n796), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U884 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U885 ( .A(n801), .B(KEYINPUT75), .ZN(n831) );
  XNOR2_X1 U886 ( .A(n802), .B(n831), .ZN(n904) );
  NAND2_X1 U887 ( .A1(G559), .A2(n977), .ZN(n803) );
  XNOR2_X1 U888 ( .A(n803), .B(n991), .ZN(n830) );
  XNOR2_X1 U889 ( .A(KEYINPUT84), .B(n830), .ZN(n804) );
  XNOR2_X1 U890 ( .A(n904), .B(n804), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n805), .A2(G868), .ZN(n808) );
  NAND2_X1 U892 ( .A1(n806), .A2(n831), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n808), .A2(n807), .ZN(G295) );
  NAND2_X1 U894 ( .A1(G2078), .A2(G2084), .ZN(n809) );
  XOR2_X1 U895 ( .A(KEYINPUT20), .B(n809), .Z(n810) );
  NAND2_X1 U896 ( .A1(G2090), .A2(n810), .ZN(n811) );
  XNOR2_X1 U897 ( .A(KEYINPUT21), .B(n811), .ZN(n812) );
  NAND2_X1 U898 ( .A1(n812), .A2(G2072), .ZN(n813) );
  XOR2_X1 U899 ( .A(KEYINPUT85), .B(n813), .Z(G158) );
  XNOR2_X1 U900 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U901 ( .A1(G235), .A2(G236), .ZN(n814) );
  XOR2_X1 U902 ( .A(KEYINPUT88), .B(n814), .Z(n815) );
  NOR2_X1 U903 ( .A1(G238), .A2(n815), .ZN(n816) );
  NAND2_X1 U904 ( .A1(G57), .A2(n816), .ZN(n834) );
  NAND2_X1 U905 ( .A1(G567), .A2(n834), .ZN(n817) );
  XNOR2_X1 U906 ( .A(n817), .B(KEYINPUT89), .ZN(n824) );
  NAND2_X1 U907 ( .A1(G132), .A2(G82), .ZN(n818) );
  XNOR2_X1 U908 ( .A(n818), .B(KEYINPUT22), .ZN(n819) );
  XNOR2_X1 U909 ( .A(n819), .B(KEYINPUT86), .ZN(n820) );
  NOR2_X1 U910 ( .A1(G218), .A2(n820), .ZN(n821) );
  XNOR2_X1 U911 ( .A(n821), .B(KEYINPUT87), .ZN(n822) );
  OR2_X1 U912 ( .A1(G221), .A2(n822), .ZN(n835) );
  AND2_X1 U913 ( .A1(G2106), .A2(n835), .ZN(n823) );
  NOR2_X1 U914 ( .A1(n824), .A2(n823), .ZN(G319) );
  INV_X1 U915 ( .A(G319), .ZN(n826) );
  NAND2_X1 U916 ( .A1(G661), .A2(G483), .ZN(n825) );
  NOR2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n829) );
  NAND2_X1 U918 ( .A1(n829), .A2(G36), .ZN(G176) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n923), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U921 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(G188) );
  NOR2_X1 U925 ( .A1(n830), .A2(G860), .ZN(n833) );
  XOR2_X1 U926 ( .A(n831), .B(KEYINPUT74), .Z(n832) );
  XNOR2_X1 U927 ( .A(n833), .B(n832), .ZN(G145) );
  INV_X1 U928 ( .A(G132), .ZN(G219) );
  INV_X1 U929 ( .A(G82), .ZN(G220) );
  NOR2_X1 U930 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  XOR2_X1 U932 ( .A(G2100), .B(G2096), .Z(n837) );
  XNOR2_X1 U933 ( .A(KEYINPUT42), .B(G2678), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U935 ( .A(KEYINPUT43), .B(G2090), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U938 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U939 ( .A(G2078), .B(G2084), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(G227) );
  XNOR2_X1 U941 ( .A(n844), .B(G1976), .ZN(n847) );
  XOR2_X1 U942 ( .A(n845), .B(G1971), .Z(n846) );
  XNOR2_X1 U943 ( .A(n847), .B(n846), .ZN(n857) );
  XOR2_X1 U944 ( .A(KEYINPUT108), .B(G2474), .Z(n849) );
  XNOR2_X1 U945 ( .A(G1981), .B(KEYINPUT110), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U947 ( .A(G1986), .B(G1956), .Z(n851) );
  XNOR2_X1 U948 ( .A(G1966), .B(G1961), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U950 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U951 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G136), .A2(n889), .ZN(n864) );
  NAND2_X1 U955 ( .A1(n885), .A2(G112), .ZN(n859) );
  NAND2_X1 U956 ( .A1(G100), .A2(n890), .ZN(n858) );
  NAND2_X1 U957 ( .A1(n859), .A2(n858), .ZN(n862) );
  NAND2_X1 U958 ( .A1(n886), .A2(G124), .ZN(n860) );
  XOR2_X1 U959 ( .A(KEYINPUT44), .B(n860), .Z(n861) );
  NOR2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n865), .B(KEYINPUT111), .ZN(G162) );
  XNOR2_X1 U963 ( .A(n866), .B(G162), .ZN(n868) );
  XNOR2_X1 U964 ( .A(G160), .B(G164), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U966 ( .A(KEYINPUT115), .B(KEYINPUT48), .Z(n870) );
  XNOR2_X1 U967 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U969 ( .A(n872), .B(n871), .Z(n884) );
  NAND2_X1 U970 ( .A1(n889), .A2(G139), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G103), .A2(n890), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U973 ( .A(KEYINPUT112), .B(n875), .ZN(n881) );
  NAND2_X1 U974 ( .A1(G115), .A2(n885), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G127), .A2(n886), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U977 ( .A(KEYINPUT47), .B(n878), .ZN(n879) );
  XNOR2_X1 U978 ( .A(KEYINPUT113), .B(n879), .ZN(n880) );
  NOR2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n941) );
  XNOR2_X1 U980 ( .A(n882), .B(n941), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n900) );
  NAND2_X1 U982 ( .A1(G118), .A2(n885), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G130), .A2(n886), .ZN(n887) );
  NAND2_X1 U984 ( .A1(n888), .A2(n887), .ZN(n895) );
  NAND2_X1 U985 ( .A1(n889), .A2(G142), .ZN(n892) );
  NAND2_X1 U986 ( .A1(G106), .A2(n890), .ZN(n891) );
  NAND2_X1 U987 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U988 ( .A(n893), .B(KEYINPUT45), .Z(n894) );
  NOR2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U990 ( .A(n896), .B(n926), .ZN(n897) );
  XOR2_X1 U991 ( .A(n898), .B(n897), .Z(n899) );
  XNOR2_X1 U992 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U993 ( .A1(G37), .A2(n901), .ZN(G395) );
  XNOR2_X1 U994 ( .A(n991), .B(KEYINPUT116), .ZN(n903) );
  XOR2_X1 U995 ( .A(G301), .B(n977), .Z(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n906) );
  XOR2_X1 U997 ( .A(n904), .B(G286), .Z(n905) );
  XNOR2_X1 U998 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U999 ( .A1(G37), .A2(n907), .ZN(G397) );
  XOR2_X1 U1000 ( .A(G2451), .B(G2430), .Z(n909) );
  XNOR2_X1 U1001 ( .A(G2438), .B(G2443), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n909), .B(n908), .ZN(n915) );
  XOR2_X1 U1003 ( .A(G2435), .B(G2454), .Z(n911) );
  XNOR2_X1 U1004 ( .A(G1341), .B(G1348), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n913) );
  XOR2_X1 U1006 ( .A(G2446), .B(G2427), .Z(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1008 ( .A(n915), .B(n914), .Z(n916) );
  NAND2_X1 U1009 ( .A1(G14), .A2(n916), .ZN(n922) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n922), .ZN(n919) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G57), .ZN(G237) );
  INV_X1 U1018 ( .A(n922), .ZN(G401) );
  INV_X1 U1019 ( .A(n923), .ZN(G223) );
  XOR2_X1 U1020 ( .A(G2084), .B(G160), .Z(n924) );
  NOR2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n927) );
  NAND2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n933) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1025 ( .A(KEYINPUT51), .B(n930), .Z(n931) );
  XNOR2_X1 U1026 ( .A(n931), .B(KEYINPUT117), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(n938), .B(KEYINPUT118), .ZN(n940) );
  NAND2_X1 U1031 ( .A1(n940), .A2(n939), .ZN(n946) );
  XOR2_X1 U1032 ( .A(G2072), .B(n941), .Z(n943) );
  XOR2_X1 U1033 ( .A(G164), .B(G2078), .Z(n942) );
  NOR2_X1 U1034 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1035 ( .A(KEYINPUT50), .B(n944), .Z(n945) );
  NOR2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n947), .ZN(n949) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1039 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1040 ( .A1(n950), .A2(G29), .ZN(n1031) );
  XNOR2_X1 U1041 ( .A(G2090), .B(G35), .ZN(n967) );
  XOR2_X1 U1042 ( .A(G1991), .B(G25), .Z(n951) );
  NAND2_X1 U1043 ( .A1(n951), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(n952), .B(KEYINPUT119), .ZN(n961) );
  XOR2_X1 U1045 ( .A(G27), .B(KEYINPUT121), .Z(n953) );
  XNOR2_X1 U1046 ( .A(n954), .B(n953), .ZN(n956) );
  XOR2_X1 U1047 ( .A(G2072), .B(G33), .Z(n955) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(KEYINPUT122), .B(G1996), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G32), .B(n957), .ZN(n958) );
  NOR2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n964) );
  XNOR2_X1 U1053 ( .A(KEYINPUT120), .B(G2067), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(G26), .B(n962), .ZN(n963) );
  NOR2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n965), .ZN(n966) );
  NOR2_X1 U1057 ( .A1(n967), .A2(n966), .ZN(n970) );
  XOR2_X1 U1058 ( .A(G2084), .B(G34), .Z(n968) );
  XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(n968), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1061 ( .A(KEYINPUT55), .B(n971), .Z(n973) );
  INV_X1 U1062 ( .A(G29), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1064 ( .A1(G11), .A2(n974), .ZN(n1029) );
  INV_X1 U1065 ( .A(G16), .ZN(n1025) );
  XOR2_X1 U1066 ( .A(n1025), .B(KEYINPUT56), .Z(n1001) );
  XOR2_X1 U1067 ( .A(G301), .B(G1961), .Z(n976) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n987) );
  XNOR2_X1 U1069 ( .A(n977), .B(G1348), .ZN(n985) );
  XNOR2_X1 U1070 ( .A(G1956), .B(KEYINPUT124), .ZN(n979) );
  XOR2_X1 U1071 ( .A(n979), .B(n978), .Z(n983) );
  NAND2_X1 U1072 ( .A1(G1971), .A2(G303), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(KEYINPUT125), .B(n990), .ZN(n999) );
  XNOR2_X1 U1079 ( .A(n991), .B(G1341), .ZN(n997) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G168), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(n994), .B(KEYINPUT123), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(KEYINPUT57), .B(n995), .ZN(n996) );
  NOR2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1027) );
  XOR2_X1 U1087 ( .A(G1986), .B(G24), .Z(n1005) );
  XNOR2_X1 U1088 ( .A(G1971), .B(G22), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(G23), .B(G1976), .ZN(n1002) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(n1007), .B(n1006), .ZN(n1020) );
  XOR2_X1 U1094 ( .A(G1348), .B(KEYINPUT59), .Z(n1008) );
  XNOR2_X1 U1095 ( .A(G4), .B(n1008), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(G20), .B(G1956), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G1981), .B(G6), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(n1015), .B(KEYINPUT60), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(KEYINPUT126), .B(G1961), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(G5), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(G21), .B(G1966), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1032), .ZN(G150) );
  INV_X1 U1115 ( .A(G150), .ZN(G311) );
endmodule

