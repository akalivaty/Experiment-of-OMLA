

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592;

  XNOR2_X2 U323 ( .A(KEYINPUT65), .B(n416), .ZN(n459) );
  OR2_X1 U324 ( .A1(n381), .A2(n380), .ZN(n382) );
  NOR2_X1 U325 ( .A1(n510), .A2(n537), .ZN(n347) );
  BUF_X1 U326 ( .A(n533), .Z(n555) );
  XOR2_X1 U327 ( .A(n346), .B(n345), .Z(n571) );
  NOR2_X1 U328 ( .A1(n577), .A2(n576), .ZN(n581) );
  XNOR2_X1 U329 ( .A(G78GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U330 ( .A(n314), .B(G148GAT), .ZN(n446) );
  INV_X1 U331 ( .A(KEYINPUT31), .ZN(n315) );
  NAND2_X1 U332 ( .A1(n415), .A2(n522), .ZN(n416) );
  XNOR2_X1 U333 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U334 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U335 ( .A(n434), .B(n433), .Z(n536) );
  XNOR2_X1 U336 ( .A(n456), .B(G197GAT), .ZN(n457) );
  XNOR2_X1 U337 ( .A(n458), .B(n457), .ZN(G1352GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n292) );
  XNOR2_X1 U339 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n291) );
  XNOR2_X1 U340 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U341 ( .A(G169GAT), .B(n293), .Z(n434) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n294), .B(G92GAT), .ZN(n374) );
  XOR2_X1 U344 ( .A(n374), .B(KEYINPUT100), .Z(n296) );
  NAND2_X1 U345 ( .A1(G226GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n299) );
  XNOR2_X1 U347 ( .A(G218GAT), .B(G204GAT), .ZN(n297) );
  XOR2_X1 U348 ( .A(G176GAT), .B(G64GAT), .Z(n311) );
  XNOR2_X1 U349 ( .A(n297), .B(n311), .ZN(n298) );
  XOR2_X1 U350 ( .A(n299), .B(n298), .Z(n303) );
  XNOR2_X1 U351 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n300), .B(KEYINPUT92), .ZN(n445) );
  XNOR2_X1 U353 ( .A(G8GAT), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U354 ( .A(n301), .B(G211GAT), .ZN(n353) );
  XNOR2_X1 U355 ( .A(n445), .B(n353), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U357 ( .A(n434), .B(n304), .Z(n501) );
  INV_X1 U358 ( .A(n501), .ZN(n524) );
  XNOR2_X1 U359 ( .A(G71GAT), .B(G57GAT), .ZN(n310) );
  INV_X1 U360 ( .A(KEYINPUT13), .ZN(n305) );
  NAND2_X1 U361 ( .A1(n305), .A2(KEYINPUT67), .ZN(n308) );
  INV_X1 U362 ( .A(KEYINPUT67), .ZN(n306) );
  NAND2_X1 U363 ( .A1(n306), .A2(KEYINPUT13), .ZN(n307) );
  NAND2_X1 U364 ( .A1(n308), .A2(n307), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n354) );
  XNOR2_X1 U366 ( .A(n354), .B(n311), .ZN(n313) );
  AND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n446), .B(KEYINPUT69), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U372 ( .A(KEYINPUT68), .B(KEYINPUT72), .Z(n320) );
  XNOR2_X1 U373 ( .A(G120GAT), .B(G92GAT), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n330) );
  XOR2_X1 U376 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n324) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(G85GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U379 ( .A(G99GAT), .B(n325), .Z(n378) );
  XOR2_X1 U380 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n327) );
  XNOR2_X1 U381 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U383 ( .A(n378), .B(n328), .Z(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n582) );
  XOR2_X1 U385 ( .A(n582), .B(KEYINPUT64), .Z(n331) );
  XOR2_X1 U386 ( .A(KEYINPUT41), .B(n331), .Z(n561) );
  INV_X1 U387 ( .A(n561), .ZN(n510) );
  XOR2_X1 U388 ( .A(G22GAT), .B(G141GAT), .Z(n333) );
  XNOR2_X1 U389 ( .A(G169GAT), .B(G15GAT), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U391 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n335) );
  XNOR2_X1 U392 ( .A(G197GAT), .B(G8GAT), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n346) );
  XOR2_X1 U395 ( .A(G29GAT), .B(G43GAT), .Z(n339) );
  XNOR2_X1 U396 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n365) );
  XOR2_X1 U398 ( .A(n365), .B(KEYINPUT29), .Z(n341) );
  NAND2_X1 U399 ( .A1(G229GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U401 ( .A(G113GAT), .B(G1GAT), .Z(n404) );
  XOR2_X1 U402 ( .A(n342), .B(n404), .Z(n344) );
  XNOR2_X1 U403 ( .A(G50GAT), .B(G36GAT), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n345) );
  INV_X1 U405 ( .A(n571), .ZN(n537) );
  XNOR2_X1 U406 ( .A(n347), .B(KEYINPUT46), .ZN(n381) );
  XOR2_X1 U407 ( .A(KEYINPUT14), .B(KEYINPUT83), .Z(n349) );
  XNOR2_X1 U408 ( .A(KEYINPUT15), .B(KEYINPUT12), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n364) );
  XOR2_X1 U410 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n351) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U413 ( .A(n352), .B(KEYINPUT82), .Z(n356) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U416 ( .A(KEYINPUT81), .B(G64GAT), .Z(n358) );
  XOR2_X1 U417 ( .A(G15GAT), .B(G127GAT), .Z(n426) );
  XOR2_X1 U418 ( .A(G22GAT), .B(G155GAT), .Z(n438) );
  XNOR2_X1 U419 ( .A(n426), .B(n438), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U421 ( .A(n360), .B(n359), .Z(n362) );
  XNOR2_X1 U422 ( .A(G1GAT), .B(G78GAT), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n492) );
  XOR2_X1 U425 ( .A(n492), .B(KEYINPUT110), .Z(n573) );
  XOR2_X1 U426 ( .A(KEYINPUT11), .B(n365), .Z(n367) );
  NAND2_X1 U427 ( .A1(G232GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U429 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n369) );
  XNOR2_X1 U430 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U432 ( .A(n371), .B(n370), .Z(n376) );
  XOR2_X1 U433 ( .A(G162GAT), .B(KEYINPUT76), .Z(n373) );
  XNOR2_X1 U434 ( .A(G50GAT), .B(G218GAT), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n450) );
  XNOR2_X1 U436 ( .A(n450), .B(n374), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n567) );
  INV_X1 U439 ( .A(n567), .ZN(n379) );
  OR2_X1 U440 ( .A1(n573), .A2(n379), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n382), .B(KEYINPUT47), .ZN(n387) );
  XNOR2_X1 U442 ( .A(KEYINPUT78), .B(n567), .ZN(n577) );
  XNOR2_X1 U443 ( .A(KEYINPUT36), .B(n577), .ZN(n589) );
  NOR2_X1 U444 ( .A1(n589), .A2(n492), .ZN(n383) );
  XNOR2_X1 U445 ( .A(KEYINPUT45), .B(n383), .ZN(n384) );
  NAND2_X1 U446 ( .A1(n384), .A2(n582), .ZN(n385) );
  NOR2_X1 U447 ( .A1(n571), .A2(n385), .ZN(n386) );
  NOR2_X1 U448 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n388), .B(KEYINPUT48), .ZN(n533) );
  NOR2_X1 U450 ( .A1(n524), .A2(n533), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n389), .B(KEYINPUT54), .ZN(n415) );
  XOR2_X1 U452 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n391) );
  XNOR2_X1 U453 ( .A(KEYINPUT94), .B(KEYINPUT99), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U455 ( .A(G57GAT), .B(KEYINPUT95), .Z(n393) );
  XNOR2_X1 U456 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U458 ( .A(n395), .B(n394), .Z(n400) );
  XOR2_X1 U459 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n397) );
  NAND2_X1 U460 ( .A1(G225GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U462 ( .A(KEYINPUT98), .B(n398), .ZN(n399) );
  XNOR2_X1 U463 ( .A(n400), .B(n399), .ZN(n408) );
  XOR2_X1 U464 ( .A(G85GAT), .B(G155GAT), .Z(n402) );
  XNOR2_X1 U465 ( .A(G127GAT), .B(G148GAT), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U467 ( .A(n403), .B(G162GAT), .Z(n406) );
  XNOR2_X1 U468 ( .A(n404), .B(G29GAT), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U470 ( .A(n408), .B(n407), .Z(n414) );
  XOR2_X1 U471 ( .A(G120GAT), .B(KEYINPUT84), .Z(n410) );
  XNOR2_X1 U472 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n425) );
  XOR2_X1 U474 ( .A(G141GAT), .B(KEYINPUT3), .Z(n411) );
  XOR2_X1 U475 ( .A(KEYINPUT2), .B(n411), .Z(n451) );
  INV_X1 U476 ( .A(n451), .ZN(n412) );
  XOR2_X1 U477 ( .A(n425), .B(n412), .Z(n413) );
  XOR2_X1 U478 ( .A(n414), .B(n413), .Z(n522) );
  XOR2_X1 U479 ( .A(G71GAT), .B(G99GAT), .Z(n418) );
  XNOR2_X1 U480 ( .A(G43GAT), .B(G190GAT), .ZN(n417) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U482 ( .A(G176GAT), .B(KEYINPUT87), .Z(n420) );
  XNOR2_X1 U483 ( .A(G113GAT), .B(KEYINPUT85), .ZN(n419) );
  XNOR2_X1 U484 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U485 ( .A(n422), .B(n421), .Z(n432) );
  XOR2_X1 U486 ( .A(G183GAT), .B(KEYINPUT89), .Z(n424) );
  XNOR2_X1 U487 ( .A(KEYINPUT20), .B(KEYINPUT88), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U489 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U490 ( .A1(G227GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U494 ( .A(KEYINPUT93), .B(KEYINPUT24), .Z(n436) );
  XNOR2_X1 U495 ( .A(G106GAT), .B(KEYINPUT23), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U497 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U500 ( .A(KEYINPUT22), .B(KEYINPUT90), .Z(n442) );
  XNOR2_X1 U501 ( .A(G211GAT), .B(KEYINPUT91), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U503 ( .A(n444), .B(n443), .Z(n448) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n452) );
  XOR2_X1 U507 ( .A(n452), .B(n451), .Z(n477) );
  NOR2_X1 U508 ( .A1(n536), .A2(n477), .ZN(n453) );
  XOR2_X1 U509 ( .A(KEYINPUT26), .B(n453), .Z(n454) );
  XNOR2_X1 U510 ( .A(KEYINPUT101), .B(n454), .ZN(n552) );
  NAND2_X1 U511 ( .A1(n459), .A2(n552), .ZN(n455) );
  XNOR2_X1 U512 ( .A(KEYINPUT126), .B(n455), .ZN(n590) );
  INV_X1 U513 ( .A(n590), .ZN(n585) );
  NAND2_X1 U514 ( .A1(n585), .A2(n571), .ZN(n458) );
  XOR2_X1 U515 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n456) );
  NAND2_X1 U516 ( .A1(n459), .A2(n477), .ZN(n463) );
  XOR2_X1 U517 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n461) );
  INV_X1 U518 ( .A(KEYINPUT55), .ZN(n460) );
  INV_X1 U519 ( .A(n536), .ZN(n526) );
  NOR2_X2 U520 ( .A1(n464), .A2(n526), .ZN(n575) );
  AND2_X1 U521 ( .A1(n575), .A2(n561), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n466) );
  XNOR2_X1 U523 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n468), .B(n467), .ZN(G1349GAT) );
  NAND2_X1 U526 ( .A1(n571), .A2(n582), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n469), .B(KEYINPUT75), .ZN(n496) );
  INV_X1 U528 ( .A(n522), .ZN(n498) );
  NAND2_X1 U529 ( .A1(n536), .A2(n501), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n477), .A2(n470), .ZN(n471) );
  XOR2_X1 U531 ( .A(KEYINPUT25), .B(n471), .Z(n473) );
  XNOR2_X1 U532 ( .A(KEYINPUT27), .B(n501), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n552), .A2(n476), .ZN(n472) );
  NAND2_X1 U534 ( .A1(n473), .A2(n472), .ZN(n474) );
  XOR2_X1 U535 ( .A(KEYINPUT102), .B(n474), .Z(n475) );
  NOR2_X1 U536 ( .A1(n498), .A2(n475), .ZN(n479) );
  AND2_X1 U537 ( .A1(n476), .A2(n498), .ZN(n553) );
  XOR2_X1 U538 ( .A(KEYINPUT28), .B(n477), .Z(n507) );
  INV_X1 U539 ( .A(n507), .ZN(n529) );
  NAND2_X1 U540 ( .A1(n553), .A2(n529), .ZN(n534) );
  NOR2_X1 U541 ( .A1(n536), .A2(n534), .ZN(n478) );
  NOR2_X1 U542 ( .A1(n479), .A2(n478), .ZN(n491) );
  INV_X1 U543 ( .A(n492), .ZN(n586) );
  NAND2_X1 U544 ( .A1(n577), .A2(n586), .ZN(n480) );
  XNOR2_X1 U545 ( .A(KEYINPUT16), .B(n480), .ZN(n481) );
  NOR2_X1 U546 ( .A1(n491), .A2(n481), .ZN(n482) );
  XOR2_X1 U547 ( .A(KEYINPUT103), .B(n482), .Z(n511) );
  NAND2_X1 U548 ( .A1(n496), .A2(n511), .ZN(n489) );
  NOR2_X1 U549 ( .A1(n522), .A2(n489), .ZN(n483) );
  XOR2_X1 U550 ( .A(G1GAT), .B(n483), .Z(n484) );
  XNOR2_X1 U551 ( .A(KEYINPUT34), .B(n484), .ZN(G1324GAT) );
  NOR2_X1 U552 ( .A1(n524), .A2(n489), .ZN(n485) );
  XOR2_X1 U553 ( .A(KEYINPUT104), .B(n485), .Z(n486) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U555 ( .A1(n526), .A2(n489), .ZN(n488) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U557 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  NOR2_X1 U558 ( .A1(n529), .A2(n489), .ZN(n490) );
  XOR2_X1 U559 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  XOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .Z(n500) );
  XOR2_X1 U561 ( .A(KEYINPUT37), .B(KEYINPUT105), .Z(n495) );
  NOR2_X1 U562 ( .A1(n491), .A2(n589), .ZN(n493) );
  NAND2_X1 U563 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U564 ( .A(n495), .B(n494), .ZN(n521) );
  NAND2_X1 U565 ( .A1(n496), .A2(n521), .ZN(n497) );
  XOR2_X1 U566 ( .A(KEYINPUT38), .B(n497), .Z(n508) );
  NAND2_X1 U567 ( .A1(n498), .A2(n508), .ZN(n499) );
  XNOR2_X1 U568 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NAND2_X1 U569 ( .A1(n508), .A2(n501), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n502), .B(KEYINPUT106), .ZN(n503) );
  XNOR2_X1 U571 ( .A(G36GAT), .B(n503), .ZN(G1329GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n505) );
  NAND2_X1 U573 ( .A1(n536), .A2(n508), .ZN(n504) );
  XNOR2_X1 U574 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U575 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NAND2_X1 U576 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U578 ( .A1(n571), .A2(n510), .ZN(n520) );
  NAND2_X1 U579 ( .A1(n511), .A2(n520), .ZN(n517) );
  NOR2_X1 U580 ( .A1(n522), .A2(n517), .ZN(n512) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n512), .Z(n513) );
  XNOR2_X1 U582 ( .A(KEYINPUT42), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U583 ( .A1(n524), .A2(n517), .ZN(n514) );
  XOR2_X1 U584 ( .A(KEYINPUT108), .B(n514), .Z(n515) );
  XNOR2_X1 U585 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NOR2_X1 U586 ( .A1(n526), .A2(n517), .ZN(n516) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n529), .A2(n517), .ZN(n519) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U590 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U591 ( .A1(n521), .A2(n520), .ZN(n528) );
  NOR2_X1 U592 ( .A1(n522), .A2(n528), .ZN(n523) );
  XOR2_X1 U593 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U594 ( .A1(n524), .A2(n528), .ZN(n525) );
  XOR2_X1 U595 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U596 ( .A1(n526), .A2(n528), .ZN(n527) );
  XOR2_X1 U597 ( .A(G99GAT), .B(n527), .Z(G1338GAT) );
  NOR2_X1 U598 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U599 ( .A(KEYINPUT109), .B(KEYINPUT44), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U602 ( .A1(n555), .A2(n534), .ZN(n535) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n547) );
  NOR2_X1 U604 ( .A1(n537), .A2(n547), .ZN(n538) );
  XOR2_X1 U605 ( .A(G113GAT), .B(n538), .Z(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n540) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(n542) );
  NOR2_X1 U609 ( .A1(n510), .A2(n547), .ZN(n541) );
  XOR2_X1 U610 ( .A(n542), .B(n541), .Z(n543) );
  XNOR2_X1 U611 ( .A(KEYINPUT111), .B(n543), .ZN(G1341GAT) );
  INV_X1 U612 ( .A(n547), .ZN(n544) );
  NAND2_X1 U613 ( .A1(n573), .A2(n544), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n545), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  NOR2_X1 U616 ( .A1(n547), .A2(n577), .ZN(n551) );
  XOR2_X1 U617 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n549) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT115), .ZN(n548) );
  XNOR2_X1 U619 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n571), .A2(n565), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT116), .ZN(n557) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(n557), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n559) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U629 ( .A(KEYINPUT52), .B(n560), .Z(n563) );
  NAND2_X1 U630 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n586), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U634 ( .A(n565), .ZN(n566) );
  NOR2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n569) );
  XNOR2_X1 U636 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U638 ( .A(G162GAT), .B(n570), .ZN(G1347GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n571), .ZN(n572) );
  XNOR2_X1 U640 ( .A(G169GAT), .B(n572), .ZN(G1348GAT) );
  NAND2_X1 U641 ( .A1(n573), .A2(n575), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U643 ( .A(n575), .ZN(n576) );
  XNOR2_X1 U644 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(KEYINPUT124), .ZN(n579) );
  XNOR2_X1 U646 ( .A(KEYINPUT125), .B(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1351GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  OR2_X1 U649 ( .A1(n590), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U651 ( .A(G211GAT), .B(KEYINPUT127), .Z(n588) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

