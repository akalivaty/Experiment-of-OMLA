//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n450, new_n452, new_n453,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n563, new_n564, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n449));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  INV_X1    g026(.A(new_n450), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n452), .A2(G567), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(G234));
  NAND2_X1  g029(.A1(new_n452), .A2(G2106), .ZN(G217));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  INV_X1    g035(.A(G2106), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OAI22_X1  g037(.A1(new_n457), .A2(new_n461), .B1(new_n462), .B2(new_n458), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT67), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n472), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n466), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT70), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n473), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n472), .A2(new_n466), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G138), .B(new_n466), .C1(new_n470), .C2(new_n471), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT4), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n484), .B2(G126), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  OR2_X1    g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n498), .A2(new_n499), .B1(KEYINPUT6), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(new_n500), .B2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT71), .A3(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n501), .A2(new_n502), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n502), .B1(new_n501), .B2(new_n507), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G88), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(KEYINPUT6), .B2(new_n500), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n507), .A2(G50), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT72), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n498), .A2(new_n499), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n517), .A2(new_n500), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n511), .A2(new_n515), .A3(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT75), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  AND2_X1   g098(.A1(G63), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n523), .B1(new_n516), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n505), .A2(KEYINPUT71), .A3(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT71), .B1(new_n505), .B2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n513), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT74), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n507), .A2(new_n530), .A3(new_n513), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G51), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n510), .A2(G89), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n525), .A2(new_n533), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AND2_X1   g112(.A1(KEYINPUT5), .A2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(KEYINPUT5), .A2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n532), .A2(G52), .B1(G651), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n526), .A2(new_n527), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n538), .A2(new_n539), .B1(new_n505), .B2(G651), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT73), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n501), .A2(new_n502), .A3(new_n507), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n546), .A2(G90), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n543), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  AND3_X1   g125(.A1(new_n507), .A2(new_n530), .A3(new_n513), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n530), .B1(new_n507), .B2(new_n513), .ZN(new_n552));
  OAI21_X1  g127(.A(G43), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n546), .A2(G81), .A3(new_n547), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n540), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n553), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(new_n510), .A2(G91), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n507), .A2(G53), .A3(new_n513), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  XNOR2_X1  g144(.A(KEYINPUT76), .B(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n540), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n566), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G299));
  OAI21_X1  g149(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n575));
  INV_X1    g150(.A(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n528), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n510), .B2(G87), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G288));
  NAND3_X1  g154(.A1(new_n546), .A2(G86), .A3(new_n547), .ZN(new_n580));
  INV_X1    g155(.A(new_n528), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n540), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n581), .A2(G48), .B1(new_n584), .B2(G651), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n580), .A2(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n540), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g166(.A(KEYINPUT77), .B(new_n587), .C1(new_n540), .C2(new_n588), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n591), .A2(G651), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(G47), .B1(new_n551), .B2(new_n552), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n546), .A2(G85), .A3(new_n547), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n593), .A2(new_n594), .A3(new_n595), .A4(KEYINPUT78), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G290));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(G301), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n540), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n532), .A2(G54), .B1(G651), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n546), .A2(G92), .A3(new_n547), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(KEYINPUT79), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n546), .A2(new_n610), .A3(G92), .A4(new_n547), .ZN(new_n611));
  AND3_X1   g186(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n609), .B1(new_n608), .B2(new_n611), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(KEYINPUT80), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(KEYINPUT80), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n602), .B1(new_n617), .B2(new_n601), .ZN(G284));
  AOI21_X1  g193(.A(new_n602), .B1(new_n617), .B2(new_n601), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n573), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(G868), .B2(new_n573), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND3_X1  g199(.A1(new_n615), .A2(new_n623), .A3(new_n616), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n484), .A2(G123), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT81), .Z(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(G111), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G2105), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(new_n473), .B2(G135), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n468), .A2(new_n476), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n636), .A2(new_n641), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT83), .Z(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n650), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(G14), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NOR2_X1   g237(.A1(G2072), .A2(G2078), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n444), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n665), .B2(KEYINPUT84), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(KEYINPUT84), .B2(new_n665), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n664), .B(KEYINPUT17), .ZN(new_n670));
  INV_X1    g245(.A(new_n662), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n667), .B(new_n669), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n669), .A2(new_n664), .A3(new_n671), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n671), .A3(new_n668), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n683), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT20), .Z(new_n687));
  AOI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n680), .C2(new_n684), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT85), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(G229));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G32), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n484), .A2(G129), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT93), .Z(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT94), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT26), .ZN(new_n704));
  AOI22_X1  g279(.A1(G105), .A2(new_n468), .B1(new_n473), .B2(G141), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n701), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n699), .B1(new_n707), .B2(new_n698), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT27), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1996), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n473), .A2(G139), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT91), .Z(new_n712));
  NAND3_X1  g287(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT25), .Z(new_n714));
  AOI22_X1  g289(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n466), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(new_n698), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n698), .B2(G33), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G20), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT23), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n573), .B2(new_n721), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n720), .A2(new_n442), .B1(G1956), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n560), .A2(new_n721), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n721), .B2(G19), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G171), .A2(new_n721), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G5), .B2(new_n721), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  AOI22_X1  g306(.A1(G1341), .A2(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n710), .A2(new_n725), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G34), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n734), .B2(KEYINPUT24), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(KEYINPUT24), .B2(new_n734), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n481), .B2(new_n698), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2084), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G35), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G162), .B2(G29), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT29), .B(G2090), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G27), .A2(G29), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G164), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(new_n443), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n738), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  OAI22_X1  g321(.A1(new_n720), .A2(new_n442), .B1(G1341), .B2(new_n728), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n698), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n473), .A2(G140), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n484), .A2(G128), .ZN(new_n752));
  OR2_X1    g327(.A1(G104), .A2(G2105), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n753), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT89), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n750), .B1(new_n759), .B2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2067), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G1956), .B2(new_n724), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n733), .A2(new_n746), .A3(new_n747), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n617), .A2(new_n721), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G4), .B2(new_n721), .ZN(new_n765));
  INV_X1    g340(.A(G1348), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT30), .B(G28), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(new_n698), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n769), .B(new_n771), .C1(new_n635), .C2(new_n698), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n721), .A2(G21), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G168), .B2(new_n721), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n772), .B1(new_n774), .B2(G1966), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n775), .B1(new_n731), .B2(new_n730), .C1(G1966), .C2(new_n774), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT95), .Z(new_n777));
  NAND4_X1  g352(.A1(new_n763), .A2(new_n767), .A3(new_n768), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT36), .ZN(new_n779));
  NOR2_X1   g354(.A1(G25), .A2(G29), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n473), .A2(G131), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n484), .A2(G119), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n466), .A2(G107), .ZN(new_n783));
  OAI21_X1  g358(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n781), .B(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT86), .Z(new_n786));
  AOI21_X1  g361(.A(new_n780), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT35), .B(G1991), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT87), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n787), .B(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(G16), .A2(G24), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G290), .B2(new_n721), .ZN(new_n792));
  INV_X1    g367(.A(G1986), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n793), .B2(new_n792), .ZN(new_n797));
  NOR2_X1   g372(.A1(G6), .A2(G16), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n580), .A2(new_n585), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT32), .ZN(new_n801));
  INV_X1    g376(.A(G1981), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n721), .A2(G23), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n578), .B2(new_n721), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT33), .B(G1976), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n721), .A2(G22), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G166), .B2(new_n721), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n807), .B1(G1971), .B2(new_n809), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n803), .B(new_n810), .C1(G1971), .C2(new_n809), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT88), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT34), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n797), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n811), .B(KEYINPUT88), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n779), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n815), .A2(new_n779), .A3(new_n817), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n778), .B1(new_n819), .B2(new_n820), .ZN(G311));
  INV_X1    g396(.A(new_n778), .ZN(new_n822));
  INV_X1    g397(.A(new_n820), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n818), .ZN(G150));
  OAI21_X1  g399(.A(G55), .B1(new_n551), .B2(new_n552), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n546), .A2(G93), .A3(new_n547), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n500), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n825), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G860), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT37), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n617), .A2(G559), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT38), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n532), .A2(G43), .B1(G651), .B2(new_n557), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n828), .B1(new_n532), .B2(G55), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n554), .A4(new_n826), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n830), .A2(new_n559), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT38), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n617), .A2(new_n840), .A3(G559), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n834), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n839), .B1(new_n834), .B2(new_n841), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT96), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g421(.A(KEYINPUT96), .B(new_n845), .C1(new_n842), .C2(new_n843), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n844), .B2(new_n845), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n832), .B1(new_n849), .B2(new_n851), .ZN(G145));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n481), .A2(KEYINPUT97), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n481), .A2(KEYINPUT97), .ZN(new_n856));
  OAI21_X1  g431(.A(G162), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n856), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n858), .A2(new_n488), .A3(new_n854), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n635), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n857), .A2(new_n859), .A3(new_n630), .A4(new_n634), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n759), .A2(G164), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n759), .A2(G164), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n706), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n707), .A3(new_n864), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n718), .ZN(new_n871));
  INV_X1    g446(.A(new_n786), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n484), .A2(G130), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n466), .A2(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n473), .A2(KEYINPUT98), .A3(G142), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT98), .B1(new_n473), .B2(G142), .ZN(new_n877));
  OAI221_X1 g452(.A(new_n873), .B1(new_n874), .B2(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(new_n638), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n638), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n872), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n786), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n881), .A2(new_n883), .A3(new_n885), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n867), .B(new_n869), .C1(new_n712), .C2(new_n716), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n871), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n871), .A2(new_n889), .B1(new_n887), .B2(new_n888), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n863), .B(new_n890), .C1(new_n891), .C2(KEYINPUT101), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(KEYINPUT101), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n853), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n863), .A2(new_n890), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n891), .A2(KEYINPUT101), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n896), .A2(new_n897), .A3(KEYINPUT102), .A4(new_n893), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n871), .A2(new_n889), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n887), .A2(new_n888), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n863), .B1(new_n902), .B2(new_n890), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(G37), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(G395));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n608), .A2(new_n611), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT10), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n573), .B1(new_n912), .B2(new_n606), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n573), .B(new_n606), .C1(new_n612), .C2(new_n613), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n908), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n614), .A2(G299), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(KEYINPUT105), .A3(new_n914), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n839), .B(KEYINPUT104), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n920), .A2(new_n615), .A3(new_n623), .A4(new_n616), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n837), .A2(new_n838), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT104), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n625), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n919), .A2(new_n921), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n921), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n913), .B2(new_n915), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n914), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT106), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n919), .A2(new_n921), .A3(new_n924), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n926), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n935));
  NAND2_X1  g510(.A1(G303), .A2(new_n799), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n511), .A2(G305), .A3(new_n515), .A4(new_n518), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n598), .A2(new_n578), .A3(new_n599), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n578), .B1(new_n598), .B2(new_n599), .ZN(new_n940));
  OAI211_X1 g515(.A(KEYINPUT107), .B(new_n938), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT107), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(new_n938), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT107), .B1(new_n939), .B2(new_n940), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n947), .B(new_n926), .C1(new_n932), .C2(new_n933), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n935), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n935), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(G868), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n830), .A2(new_n601), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(G295));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n952), .ZN(G331));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT109), .B1(new_n543), .B2(new_n548), .ZN(new_n956));
  OAI21_X1  g531(.A(G52), .B1(new_n551), .B2(new_n552), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n542), .A2(G651), .ZN(new_n958));
  AND4_X1   g533(.A1(KEYINPUT109), .A2(new_n957), .A3(new_n548), .A4(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n922), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n838), .B(new_n837), .C1(new_n956), .C2(new_n959), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(G286), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(G168), .A3(new_n962), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n929), .A2(new_n964), .A3(new_n930), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT110), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n961), .A2(G168), .A3(new_n962), .ZN(new_n968));
  AOI21_X1  g543(.A(G168), .B1(new_n961), .B2(new_n962), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n929), .A4(new_n930), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n916), .B(new_n918), .C1(new_n968), .C2(new_n969), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n967), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n946), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n917), .B(new_n914), .C1(new_n968), .C2(new_n969), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n946), .A2(new_n966), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G37), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n955), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n946), .B1(new_n966), .B2(new_n977), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT44), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n976), .A2(new_n980), .A3(new_n984), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n985), .B1(new_n982), .B2(new_n983), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n987), .A2(new_n988), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n988), .B1(new_n987), .B2(new_n992), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(G397));
  AOI21_X1  g570(.A(G1384), .B1(new_n491), .B2(new_n495), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(KEYINPUT45), .ZN(new_n997));
  INV_X1    g572(.A(G40), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n475), .A2(new_n479), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(G1996), .A3(new_n706), .ZN(new_n1002));
  XOR2_X1   g577(.A(new_n1002), .B(KEYINPUT112), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n759), .A2(G2067), .ZN(new_n1004));
  INV_X1    g579(.A(G2067), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n757), .A2(new_n1005), .A3(new_n758), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1004), .B(new_n1006), .C1(G1996), .C2(new_n706), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1003), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n786), .A2(new_n788), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n786), .A2(new_n788), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1001), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(G290), .B(G1986), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1012), .B1(new_n1001), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1976), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(G288), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n999), .B2(new_n996), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1016), .B(new_n1018), .C1(new_n1015), .C2(G288), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1018), .B1(new_n1015), .B2(G288), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT52), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n584), .A2(G651), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  OAI21_X1  g599(.A(G1981), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(G305), .B(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(KEYINPUT49), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(KEYINPUT49), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n1018), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n999), .B1(new_n1030), .B2(new_n996), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G2090), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n996), .A2(new_n1034), .A3(new_n1030), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n996), .A2(new_n1030), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT118), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1971), .ZN(new_n1039));
  INV_X1    g614(.A(G1384), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n999), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n996), .A2(KEYINPUT45), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1039), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1017), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(G166), .B2(new_n1017), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1048));
  NAND3_X1  g623(.A1(G303), .A2(G8), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1022), .B(new_n1029), .C1(new_n1045), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1049), .ZN(new_n1053));
  AOI22_X1  g628(.A1(G303), .A2(G8), .B1(KEYINPUT114), .B2(KEYINPUT55), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1047), .A2(KEYINPUT115), .A3(new_n1049), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n1058));
  AOI21_X1  g633(.A(G2090), .B1(new_n996), .B2(new_n1030), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1032), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1059), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT113), .B1(new_n1061), .B2(new_n1031), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1060), .A2(new_n1062), .A3(new_n1044), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1057), .A2(G8), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT116), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1057), .A2(new_n1066), .A3(G8), .A4(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1051), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n996), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT50), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(new_n999), .A3(new_n1036), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n731), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n997), .A2(new_n443), .A3(new_n999), .A4(new_n1041), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1073), .A2(new_n1074), .A3(KEYINPUT53), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT53), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1068), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n1081));
  INV_X1    g656(.A(G1966), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT119), .B(new_n1082), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1083));
  INV_X1    g658(.A(G2084), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1070), .A2(new_n1084), .A3(new_n999), .A4(new_n1036), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n997), .A2(new_n999), .A3(new_n1041), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT119), .B1(new_n1087), .B2(new_n1082), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(G168), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(G1966), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(G168), .A3(new_n1085), .A4(new_n1083), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G8), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT51), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1097), .A3(G8), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1081), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1081), .A3(new_n1098), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1080), .A2(new_n1100), .A3(KEYINPUT124), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n1068), .A3(new_n1079), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(new_n1099), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n573), .B(KEYINPUT57), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1032), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1108));
  INV_X1    g683(.A(G1956), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1092), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1107), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1000), .A2(new_n1069), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1071), .A2(new_n766), .B1(new_n1115), .B2(new_n1005), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n614), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1113), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1114), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(new_n1113), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1116), .A2(new_n614), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT60), .B1(new_n1122), .B2(new_n1117), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT58), .B(G1341), .ZN(new_n1124));
  OAI22_X1  g699(.A1(new_n1087), .A2(G1996), .B1(new_n1115), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n560), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT59), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1128), .A3(new_n560), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n614), .A2(KEYINPUT60), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1127), .A2(new_n1129), .B1(new_n1116), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1121), .A2(new_n1123), .A3(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1120), .A2(new_n1113), .A3(new_n1119), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1118), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1072), .A2(KEYINPUT123), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1071), .A2(new_n1138), .A3(new_n731), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1137), .B(new_n1139), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1078), .B1(G171), .B2(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1142));
  OR2_X1    g717(.A1(new_n1077), .A2(G171), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n1140), .B2(G171), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1141), .A2(new_n1142), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1135), .A2(new_n1136), .A3(new_n1068), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1022), .A2(new_n1029), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(G8), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1063), .A2(new_n1050), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1149), .A2(new_n1151), .A3(G168), .A4(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1029), .A2(new_n1015), .A3(new_n578), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(G1981), .B2(G305), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1154), .A2(KEYINPUT63), .B1(new_n1018), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1159));
  NOR2_X1   g734(.A1(G286), .A2(KEYINPUT63), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1151), .B(new_n1160), .C1(new_n1050), .C2(new_n1045), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1157), .B(new_n1158), .C1(new_n1162), .C2(new_n1148), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1156), .A2(new_n1018), .ZN(new_n1164));
  NOR4_X1   g739(.A1(new_n1148), .A2(new_n1152), .A3(new_n1150), .A4(G286), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT63), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1148), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT120), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1147), .A2(new_n1163), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1014), .B1(new_n1106), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1001), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1172), .B1(new_n1173), .B2(new_n1006), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1174), .A2(KEYINPUT125), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT46), .ZN(new_n1176));
  OR3_X1    g751(.A1(new_n1172), .A2(new_n1176), .A3(G1996), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1176), .B1(new_n1172), .B2(G1996), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n707), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1177), .B(new_n1178), .C1(new_n1172), .C2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1180), .B(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n1174), .B2(KEYINPUT125), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1172), .A2(G1986), .A3(G290), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT127), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1185), .A2(KEYINPUT48), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(KEYINPUT48), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1186), .A2(new_n1008), .A3(new_n1011), .A4(new_n1187), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1175), .A2(new_n1183), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1171), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g765(.A1(G227), .A2(new_n464), .ZN(new_n1192));
  NOR3_X1   g766(.A1(G229), .A2(G401), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n989), .A2(new_n991), .ZN(new_n1194));
  AND3_X1   g768(.A1(new_n1193), .A2(new_n905), .A3(new_n1194), .ZN(G308));
  NAND3_X1  g769(.A1(new_n1193), .A2(new_n905), .A3(new_n1194), .ZN(G225));
endmodule


