//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT65), .B(G20), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  INV_X1    g0030(.A(G264), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n209), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n213), .B(new_n220), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n229), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  AND2_X1   g0052(.A1(KEYINPUT65), .A2(G20), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT65), .A2(G20), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(KEYINPUT7), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT7), .ZN(new_n260));
  NOR4_X1   g0060(.A1(new_n256), .A2(new_n257), .A3(new_n260), .A4(G20), .ZN(new_n261));
  OAI21_X1  g0061(.A(G68), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT71), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n264), .B(G68), .C1(new_n259), .C2(new_n261), .ZN(new_n265));
  AND3_X1   g0065(.A1(KEYINPUT72), .A2(G58), .A3(G68), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT72), .B1(G58), .B2(G68), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n266), .A2(new_n267), .A3(new_n201), .ZN(new_n268));
  INV_X1    g0068(.A(G159), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n268), .A2(new_n207), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n263), .A2(KEYINPUT16), .A3(new_n265), .A4(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT16), .ZN(new_n275));
  INV_X1    g0075(.A(G68), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n255), .A2(new_n258), .A3(KEYINPUT7), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n207), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n260), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n276), .B1(new_n277), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n275), .B1(new_n284), .B2(new_n272), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT73), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(KEYINPUT73), .B(new_n275), .C1(new_n284), .C2(new_n272), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n217), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n274), .A2(new_n287), .A3(new_n288), .A4(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G13), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G1), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  XOR2_X1   g0095(.A(KEYINPUT8), .B(G58), .Z(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n290), .B1(new_n206), .B2(G20), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT68), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G41), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n279), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT68), .B1(new_n306), .B2(new_n217), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G223), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G1698), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n256), .B2(new_n257), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT74), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n280), .A2(new_n281), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(KEYINPUT74), .A3(new_n310), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(G226), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G87), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n308), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G45), .ZN(new_n322));
  AOI21_X1  g0122(.A(G1), .B1(new_n305), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n302), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G232), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(G274), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n301), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  INV_X1    g0129(.A(new_n326), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n324), .B2(G232), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n319), .B1(new_n313), .B2(new_n315), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n329), .B(new_n331), .C1(new_n332), .C2(new_n308), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n300), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n291), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(KEYINPUT17), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(KEYINPUT17), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT75), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(KEYINPUT75), .A3(KEYINPUT17), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(new_n331), .C1(new_n332), .C2(new_n308), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n321), .A2(new_n327), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(G169), .ZN(new_n345));
  INV_X1    g0145(.A(new_n300), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n291), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT18), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n341), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G1698), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n314), .A2(G226), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n314), .A2(G232), .A3(G1698), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n304), .A2(new_n307), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n330), .B1(new_n324), .B2(G238), .ZN(new_n358));
  XOR2_X1   g0158(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n359));
  AND3_X1   g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n359), .B1(new_n357), .B2(new_n358), .ZN(new_n361));
  OAI21_X1  g0161(.A(G169), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT70), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT14), .ZN(new_n364));
  INV_X1    g0164(.A(G238), .ZN(new_n365));
  OR3_X1    g0165(.A1(new_n302), .A2(new_n365), .A3(new_n323), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n326), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n356), .B2(new_n355), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n359), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT13), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n369), .B(G179), .C1(new_n370), .C2(new_n368), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT14), .ZN(new_n372));
  OAI221_X1 g0172(.A(G169), .B1(KEYINPUT70), .B2(new_n372), .C1(new_n360), .C2(new_n361), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n364), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n293), .A2(G20), .A3(new_n276), .ZN(new_n375));
  XOR2_X1   g0175(.A(new_n375), .B(KEYINPUT12), .Z(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(G68), .B2(new_n298), .ZN(new_n377));
  INV_X1    g0177(.A(new_n290), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n255), .A2(G33), .A3(G77), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n270), .A2(G50), .B1(G20), .B2(new_n276), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(KEYINPUT11), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(KEYINPUT11), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n377), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n374), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n296), .A2(new_n270), .B1(new_n219), .B2(G77), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n255), .A2(G33), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT15), .B(G87), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n290), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n298), .A2(G77), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n390), .B(new_n391), .C1(G77), .C2(new_n294), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n314), .A2(G238), .A3(G1698), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n314), .A2(G232), .A3(new_n351), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n393), .B(new_n394), .C1(new_n230), .C2(new_n314), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n356), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n330), .B1(new_n324), .B2(G244), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G169), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n396), .A2(new_n397), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(new_n342), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n392), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n296), .A2(G33), .A3(new_n255), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n270), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n290), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n294), .A2(new_n202), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n298), .B2(new_n202), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G223), .A2(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n351), .A2(G222), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n258), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G77), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n314), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n356), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g0216(.A(KEYINPUT67), .B(G226), .Z(new_n417));
  AOI21_X1  g0217(.A(new_n330), .B1(new_n324), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(new_n342), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n399), .B1(new_n416), .B2(new_n418), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n410), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n403), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n398), .A2(new_n329), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n401), .A2(new_n301), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n392), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n369), .B(G190), .C1(new_n370), .C2(new_n368), .ZN(new_n428));
  INV_X1    g0228(.A(new_n384), .ZN(new_n429));
  OAI21_X1  g0229(.A(G200), .B1(new_n360), .B2(new_n361), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n419), .A2(G200), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT9), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n410), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n407), .A2(KEYINPUT9), .A3(new_n409), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n416), .A2(G190), .A3(new_n418), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n433), .A2(new_n435), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT10), .ZN(new_n439));
  AND4_X1   g0239(.A1(new_n385), .A2(new_n427), .A3(new_n432), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n350), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT76), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n350), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT19), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n255), .B1(new_n446), .B2(new_n354), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n222), .A2(new_n224), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(G107), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n446), .B1(new_n387), .B2(new_n224), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n314), .A2(new_n255), .A3(G68), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n290), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n295), .A2(new_n388), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n206), .A2(G33), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n378), .A2(new_n294), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT78), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n294), .A2(new_n455), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT78), .B1(new_n459), .B2(new_n290), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(G87), .A3(new_n460), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n453), .A2(new_n454), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n302), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n322), .A2(G1), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n223), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n206), .A2(G45), .ZN(new_n466));
  INV_X1    g0266(.A(G274), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n463), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G244), .A2(G1698), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n365), .B2(G1698), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n314), .A2(new_n471), .B1(G33), .B2(G116), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n469), .B1(new_n308), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n301), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(G190), .B2(new_n473), .ZN(new_n475));
  INV_X1    g0275(.A(new_n388), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n458), .A2(new_n476), .A3(new_n460), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n453), .A2(new_n454), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n473), .A2(G169), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n342), .B2(new_n473), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n462), .A2(new_n475), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n314), .A2(new_n255), .A3(G87), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT22), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OR2_X1    g0285(.A1(new_n483), .A2(new_n484), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n487), .A2(G20), .B1(new_n488), .B2(new_n230), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n219), .A2(new_n488), .A3(new_n230), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT82), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n490), .B2(new_n491), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n485), .B(new_n486), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT24), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n490), .A2(new_n491), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT82), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n493), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(KEYINPUT24), .A3(new_n485), .A4(new_n486), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n498), .A2(new_n290), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n295), .A2(new_n230), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT25), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n458), .A2(new_n460), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(G107), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(KEYINPUT5), .A2(G41), .ZN(new_n509));
  NOR2_X1   g0309(.A1(KEYINPUT5), .A2(G41), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n464), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n463), .A2(new_n511), .ZN(new_n512));
  OR3_X1    g0312(.A1(new_n512), .A2(KEYINPUT83), .A3(new_n231), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n314), .A2(G257), .A3(G1698), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G294), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n314), .A2(G250), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n515), .C1(new_n516), .C2(G1698), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n356), .ZN(new_n518));
  INV_X1    g0318(.A(new_n511), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G274), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT83), .B1(new_n512), .B2(new_n231), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n513), .A2(new_n518), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n301), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(G190), .B2(new_n522), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n482), .B1(new_n508), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n520), .B1(new_n225), .B2(new_n512), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n258), .A2(new_n223), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n527), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n314), .A2(G244), .A3(new_n351), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT79), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT4), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT4), .B1(new_n529), .B2(new_n530), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n526), .B1(new_n533), .B2(new_n356), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT80), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI211_X1 g0336(.A(KEYINPUT80), .B(new_n526), .C1(new_n533), .C2(new_n356), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n399), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n526), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G283), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n516), .B2(new_n351), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n529), .A2(new_n530), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT4), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT4), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n539), .B1(new_n546), .B2(new_n308), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n458), .A2(G97), .A3(new_n460), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G97), .B2(new_n294), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n277), .A2(new_n283), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(G107), .B1(G77), .B2(new_n270), .ZN(new_n551));
  XNOR2_X1  g0351(.A(G97), .B(G107), .ZN(new_n552));
  OR2_X1    g0352(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n553));
  OR2_X1    g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n224), .A2(KEYINPUT6), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n554), .A2(new_n219), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n378), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n547), .A2(G179), .B1(new_n549), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI211_X1 g0360(.A(new_n558), .B(new_n549), .C1(new_n547), .C2(G200), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n547), .A2(KEYINPUT80), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n535), .B(new_n539), .C1(new_n546), .C2(new_n308), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(G190), .A3(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n538), .A2(new_n560), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT21), .ZN(new_n566));
  INV_X1    g0366(.A(new_n512), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(G270), .B1(G274), .B2(new_n519), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n314), .A2(G264), .A3(G1698), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n314), .A2(G257), .A3(new_n351), .ZN(new_n570));
  INV_X1    g0370(.A(G303), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n314), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n356), .ZN(new_n573));
  AOI211_X1 g0373(.A(new_n566), .B(new_n399), .C1(new_n568), .C2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n568), .A2(new_n573), .A3(G179), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n255), .B(new_n540), .C1(G33), .C2(new_n224), .ZN(new_n577));
  INV_X1    g0377(.A(G116), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n289), .A2(new_n217), .B1(G20), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT20), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(KEYINPUT20), .A3(new_n579), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n294), .A2(new_n578), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n456), .B2(new_n578), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT81), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n577), .A2(KEYINPUT20), .A3(new_n579), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT20), .B1(new_n577), .B2(new_n579), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n586), .B(KEYINPUT81), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n574), .A2(new_n576), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT81), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n568), .A2(new_n573), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(G190), .ZN(new_n597));
  AOI21_X1  g0397(.A(G200), .B1(new_n568), .B2(new_n573), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n595), .B(new_n590), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n399), .B1(new_n568), .B2(new_n573), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n595), .B2(new_n590), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n592), .B(new_n599), .C1(new_n602), .C2(KEYINPUT21), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n522), .A2(new_n342), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n522), .A2(G169), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n503), .A2(new_n507), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  AND4_X1   g0407(.A1(new_n445), .A2(new_n525), .A3(new_n565), .A4(new_n607), .ZN(G372));
  INV_X1    g0408(.A(new_n422), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n385), .B1(new_n431), .B2(new_n403), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT75), .B1(new_n335), .B2(KEYINPUT17), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT17), .ZN(new_n612));
  AOI211_X1 g0412(.A(new_n338), .B(new_n612), .C1(new_n291), .C2(new_n334), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n611), .A2(new_n613), .B1(KEYINPUT17), .B2(new_n335), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n349), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n439), .B(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n615), .B2(KEYINPUT84), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n609), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n445), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n600), .B1(new_n587), .B2(new_n591), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n596), .A2(KEYINPUT21), .A3(G169), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n575), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n595), .A2(new_n590), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n623), .A2(new_n566), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n503), .A2(new_n507), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n605), .B1(new_n342), .B2(new_n522), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n525), .A2(new_n565), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n538), .A2(new_n560), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT26), .B1(new_n633), .B2(new_n482), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n478), .A2(new_n480), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n538), .A2(new_n560), .A3(new_n481), .A4(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n621), .B1(new_n622), .B2(new_n639), .ZN(new_n640));
  XOR2_X1   g0440(.A(new_n640), .B(KEYINPUT86), .Z(G369));
  AND2_X1   g0441(.A1(new_n603), .A2(KEYINPUT87), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n255), .A2(new_n293), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n626), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n603), .B2(KEYINPUT87), .ZN(new_n650));
  OAI22_X1  g0450(.A1(new_n642), .A2(new_n650), .B1(new_n627), .B2(new_n649), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n651), .A2(G330), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n508), .A2(new_n524), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n628), .A2(new_n648), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(KEYINPUT88), .B2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n654), .A2(KEYINPUT88), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n630), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n630), .A2(new_n648), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT89), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n657), .A2(new_n659), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n627), .A2(new_n648), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n658), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n663), .A2(new_n668), .ZN(G399));
  INV_X1    g0469(.A(new_n210), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n206), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n448), .A2(G107), .A3(G116), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n672), .A2(new_n673), .B1(new_n216), .B2(new_n671), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT28), .Z(new_n675));
  NOR2_X1   g0475(.A1(new_n536), .A2(new_n537), .ZN(new_n676));
  INV_X1    g0476(.A(new_n473), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n677), .A2(new_n513), .A3(new_n518), .A4(new_n521), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n575), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT30), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n562), .A2(new_n679), .A3(KEYINPUT30), .A4(new_n563), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n677), .A2(G179), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n547), .A2(new_n522), .A3(new_n596), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n648), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT31), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT90), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n562), .A2(new_n679), .A3(new_n563), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n681), .A3(new_n683), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT90), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(KEYINPUT31), .A4(new_n648), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n685), .A2(new_n686), .ZN(new_n694));
  INV_X1    g0494(.A(new_n648), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n607), .A2(new_n525), .A3(new_n565), .A4(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n687), .A2(new_n693), .A3(new_n694), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n639), .B2(new_n648), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT91), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n627), .A2(new_n630), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n627), .B2(new_n630), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n525), .B(new_n565), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n637), .A2(new_n635), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n562), .A2(new_n563), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n559), .B1(new_n707), .B2(new_n399), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n636), .B1(new_n708), .B2(new_n481), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n648), .B1(new_n705), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n699), .B1(new_n701), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n675), .B1(new_n713), .B2(G1), .ZN(G364));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n651), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n219), .A2(new_n292), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G45), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n672), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n651), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n217), .B1(G20), .B2(new_n399), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n210), .A2(new_n314), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT92), .Z(new_n731));
  AOI22_X1  g0531(.A1(new_n731), .A2(G355), .B1(new_n578), .B2(new_n670), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n670), .A2(new_n314), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n248), .A2(new_n322), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n216), .A2(G45), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n729), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n255), .A2(G190), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n301), .A2(G179), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n230), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n219), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G97), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n739), .A2(G20), .A3(G190), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n745), .B(new_n314), .C1(new_n222), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n329), .A2(new_n301), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n219), .A2(G179), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n741), .B(new_n747), .C1(G50), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n738), .A2(G179), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n301), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(new_n301), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n755), .A2(G77), .B1(G68), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n738), .A2(new_n742), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n269), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT32), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n219), .A2(G179), .A3(G190), .A4(new_n301), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT93), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G58), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n751), .A2(new_n757), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT33), .B(G317), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n755), .A2(G311), .B1(new_n756), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n258), .B1(new_n746), .B2(new_n571), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n768), .A2(KEYINPUT94), .B1(new_n761), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n758), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(G329), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n740), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n773), .A2(G283), .B1(G294), .B2(new_n744), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G326), .A2(new_n750), .B1(new_n768), .B2(KEYINPUT94), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n767), .A2(new_n772), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n765), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n737), .B1(new_n777), .B2(new_n727), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n719), .B1(new_n726), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n721), .A2(new_n779), .ZN(G396));
  OR2_X1    g0580(.A1(new_n403), .A2(new_n648), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n392), .A2(new_n648), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n403), .B1(new_n426), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n639), .B2(new_n648), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n786), .A2(KEYINPUT96), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n695), .B(new_n784), .C1(new_n632), .C2(new_n638), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n786), .A2(KEYINPUT96), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n720), .B1(new_n790), .B2(new_n699), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n699), .B2(new_n790), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n756), .A2(G150), .B1(G137), .B2(new_n750), .ZN(new_n793));
  INV_X1    g0593(.A(G143), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n793), .B1(new_n794), .B2(new_n762), .C1(new_n269), .C2(new_n754), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT95), .B(KEYINPUT34), .Z(new_n796));
  XNOR2_X1  g0596(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n771), .A2(G132), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n773), .A2(G68), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n744), .A2(G58), .ZN(new_n800));
  INV_X1    g0600(.A(new_n746), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n258), .B1(new_n801), .B2(G50), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n798), .A2(new_n799), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n797), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n761), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G294), .A2(new_n805), .B1(new_n750), .B2(G303), .ZN(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n807), .B2(new_n758), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n756), .A2(G283), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n740), .A2(new_n222), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n314), .B1(new_n801), .B2(G107), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n809), .A2(new_n811), .A3(new_n745), .A4(new_n812), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n808), .B(new_n813), .C1(G116), .C2(new_n755), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n727), .B1(new_n804), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n727), .A2(new_n722), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n719), .B1(new_n414), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n815), .B(new_n817), .C1(new_n723), .C2(new_n784), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n792), .A2(new_n818), .ZN(G384));
  NOR2_X1   g0619(.A1(new_n717), .A2(new_n206), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n385), .A2(KEYINPUT99), .A3(new_n432), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n429), .A2(new_n695), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n385), .A2(KEYINPUT99), .A3(new_n432), .A4(new_n822), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n824), .A2(new_n784), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT104), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(KEYINPUT31), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n685), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n691), .B(new_n648), .C1(new_n827), .C2(KEYINPUT31), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n696), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT38), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n275), .A2(KEYINPUT100), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n265), .A2(new_n273), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n260), .B1(new_n314), .B2(new_n219), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n264), .B1(new_n840), .B2(G68), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n836), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n263), .A2(new_n265), .A3(new_n273), .A4(new_n835), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n290), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n346), .ZN(new_n845));
  INV_X1    g0645(.A(new_n646), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n347), .B(KEYINPUT18), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n847), .B1(new_n614), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n291), .A2(new_n346), .ZN(new_n850));
  INV_X1    g0650(.A(new_n345), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n846), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n335), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n845), .A2(new_n846), .B1(new_n291), .B2(new_n334), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n845), .A2(new_n851), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n834), .B1(new_n849), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n847), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n341), .B2(new_n349), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n857), .A2(new_n858), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n855), .B1(new_n864), .B2(new_n854), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT101), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n861), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(new_n861), .B2(new_n866), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n833), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n350), .A2(new_n853), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n852), .A2(new_n853), .A3(new_n335), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(new_n854), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n834), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n866), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n826), .A2(KEYINPUT40), .A3(new_n831), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n445), .A2(new_n831), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n882), .A2(new_n715), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n385), .A2(new_n648), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT39), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n876), .A2(new_n887), .A3(new_n866), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(new_n861), .B2(new_n866), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n886), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n824), .A2(new_n825), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n788), .B2(new_n781), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n868), .B2(new_n869), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n349), .A2(new_n646), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT102), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n891), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n894), .A2(KEYINPUT102), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n445), .A2(new_n701), .A3(new_n712), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n621), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n900), .B(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n820), .B1(new_n884), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n903), .B2(new_n884), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n219), .A2(G116), .A3(new_n218), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT35), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n909), .A2(KEYINPUT97), .B1(new_n908), .B2(new_n907), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(KEYINPUT97), .B2(new_n909), .ZN(new_n911));
  XNOR2_X1  g0711(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NOR4_X1   g0713(.A1(new_n215), .A2(new_n414), .A3(new_n266), .A4(new_n267), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n276), .A2(G50), .ZN(new_n915));
  OAI211_X1 g0715(.A(G1), .B(new_n292), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n905), .A2(new_n913), .A3(new_n916), .ZN(G367));
  INV_X1    g0717(.A(new_n727), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT46), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n746), .B2(new_n578), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n801), .A2(KEYINPUT46), .A3(G116), .ZN(new_n921));
  INV_X1    g0721(.A(new_n756), .ZN(new_n922));
  INV_X1    g0722(.A(G294), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n920), .B(new_n921), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(KEYINPUT109), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(KEYINPUT109), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT110), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n740), .A2(new_n224), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n314), .B(new_n928), .C1(G317), .C2(new_n771), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n927), .ZN(new_n931));
  INV_X1    g0731(.A(new_n744), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n932), .A2(new_n230), .B1(new_n749), .B2(new_n807), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n755), .B2(G283), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n931), .B(new_n934), .C1(new_n571), .C2(new_n762), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n932), .A2(new_n276), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G150), .B2(new_n805), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n794), .B2(new_n749), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT111), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  INV_X1    g0741(.A(G137), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n314), .B1(new_n228), .B2(new_n746), .C1(new_n758), .C2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(G77), .B2(new_n773), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n755), .A2(G50), .B1(G159), .B2(new_n756), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n941), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n930), .A2(new_n935), .B1(new_n940), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n918), .B1(new_n948), .B2(KEYINPUT47), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(KEYINPUT47), .B2(new_n948), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n244), .A2(new_n733), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n729), .B1(new_n670), .B2(new_n476), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n719), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n462), .A2(new_n695), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n481), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n635), .B2(new_n954), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n950), .B(new_n953), .C1(new_n725), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n718), .A2(G1), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n561), .A2(new_n564), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n648), .B1(new_n549), .B2(new_n558), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n633), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT106), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n708), .A2(new_n648), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(KEYINPUT44), .B1(new_n668), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n660), .A2(new_n665), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n659), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  INV_X1    g0768(.A(new_n964), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT45), .B1(new_n668), .B2(new_n964), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n668), .A2(new_n964), .A3(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n972), .A2(new_n976), .A3(new_n663), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n967), .A2(new_n969), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(new_n973), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n662), .B1(new_n980), .B2(new_n971), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT108), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n652), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n664), .A2(KEYINPUT107), .A3(new_n666), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n982), .B2(new_n652), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n664), .A2(new_n666), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n966), .A2(KEYINPUT107), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n984), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n988), .A3(new_n984), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n977), .A2(new_n981), .A3(new_n713), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n713), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n671), .B(KEYINPUT41), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n958), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n969), .A2(new_n966), .A3(KEYINPUT42), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT42), .B1(new_n969), .B2(new_n966), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n633), .B1(new_n962), .B2(new_n630), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n695), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT105), .Z(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1006), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1002), .A2(new_n1008), .A3(new_n1003), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n663), .B2(new_n969), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1007), .A2(new_n662), .A3(new_n964), .A4(new_n1009), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n957), .B1(new_n997), .B2(new_n1013), .ZN(G387));
  NAND2_X1  g0814(.A1(new_n992), .A2(new_n713), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n713), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n990), .A2(new_n1016), .A3(new_n991), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1017), .A3(new_n671), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n733), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n240), .B2(G45), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n673), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n731), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n296), .A2(new_n202), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT50), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n322), .B1(new_n276), .B2(new_n414), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1024), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1022), .A2(new_n1026), .B1(G107), .B2(new_n210), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n719), .B1(new_n1027), .B2(new_n728), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n755), .A2(G68), .B1(new_n296), .B2(new_n756), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT113), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n801), .A2(G77), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n744), .A2(new_n476), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n1032), .A3(new_n314), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n750), .A2(G159), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT112), .B(G150), .Z(new_n1035));
  OAI221_X1 g0835(.A(new_n1034), .B1(new_n202), .B2(new_n761), .C1(new_n758), .C2(new_n1035), .ZN(new_n1036));
  NOR4_X1   g0836(.A1(new_n1030), .A2(new_n928), .A3(new_n1033), .A4(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n756), .A2(G311), .B1(G322), .B2(new_n750), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n571), .B2(new_n754), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G317), .B2(new_n763), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT48), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT48), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G294), .A2(new_n801), .B1(new_n744), .B2(G283), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(G326), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n258), .B1(new_n740), .B2(new_n578), .C1(new_n1047), .C2(new_n758), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1037), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1028), .B1(new_n1051), .B2(new_n918), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT114), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1054), .A2(new_n1055), .B1(new_n664), .B2(new_n724), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n992), .B2(new_n958), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1018), .A2(new_n1057), .ZN(G393));
  NAND3_X1  g0858(.A1(new_n977), .A2(new_n981), .A3(new_n958), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n728), .B1(new_n224), .B2(new_n210), .C1(new_n1019), .C2(new_n251), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n720), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT115), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G311), .A2(new_n805), .B1(new_n750), .B2(G317), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT52), .Z(new_n1064));
  NOR2_X1   g0864(.A1(new_n754), .A2(new_n923), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n258), .B1(new_n932), .B2(new_n578), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1065), .A2(new_n741), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(G283), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n758), .A2(new_n769), .B1(new_n1068), .B2(new_n746), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT116), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n756), .A2(G303), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1064), .A2(new_n1067), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n314), .B1(new_n276), .B2(new_n746), .C1(new_n932), .C2(new_n414), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n810), .B(new_n1073), .C1(G143), .C2(new_n771), .ZN(new_n1074));
  INV_X1    g0874(.A(G150), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n761), .A2(new_n269), .B1(new_n749), .B2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n755), .A2(new_n296), .B1(G50), .B2(new_n756), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1074), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1072), .A2(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1062), .B1(new_n918), .B2(new_n1080), .C1(new_n964), .C2(new_n725), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n977), .A2(new_n981), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1015), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n993), .A2(new_n671), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1059), .B(new_n1081), .C1(new_n1084), .C2(new_n1085), .ZN(G390));
  OAI211_X1 g0886(.A(new_n888), .B(new_n890), .C1(new_n893), .C2(new_n885), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n781), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n711), .B2(new_n783), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n877), .B(new_n886), .C1(new_n892), .C2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n826), .A2(new_n697), .A3(G330), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1087), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n826), .A2(G330), .A3(new_n831), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n958), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n888), .A2(new_n890), .A3(new_n722), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1035), .A2(new_n746), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1101));
  AOI22_X1  g0901(.A1(new_n1100), .A2(new_n1101), .B1(G159), .B2(new_n744), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1101), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n258), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1102), .B(new_n1104), .C1(new_n922), .C2(new_n942), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n771), .A2(G125), .B1(G132), .B2(new_n805), .ZN(new_n1106));
  INV_X1    g0906(.A(G128), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1106), .B1(new_n202), .B2(new_n740), .C1(new_n1107), .C2(new_n749), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT54), .B(G143), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1105), .B(new_n1108), .C1(new_n755), .C2(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n771), .A2(G294), .B1(G116), .B2(new_n805), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1068), .B2(new_n749), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n258), .B1(new_n746), .B2(new_n222), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G77), .B2(new_n744), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n799), .B(new_n1115), .C1(new_n922), .C2(new_n230), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1113), .B(new_n1116), .C1(G97), .C2(new_n755), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n727), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n816), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1118), .B(new_n720), .C1(new_n296), .C2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1098), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1094), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n445), .A2(G330), .A3(new_n831), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n901), .A2(new_n1126), .A3(new_n621), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n831), .A2(G330), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT117), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n831), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n785), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n892), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1128), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n697), .A2(G330), .A3(new_n784), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n892), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1094), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n788), .A2(new_n781), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1127), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1125), .A2(new_n1141), .A3(new_n1092), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1142), .A2(new_n671), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1143), .A2(KEYINPUT118), .ZN(new_n1144));
  OAI21_X1  g0944(.A(KEYINPUT119), .B1(new_n1096), .B2(new_n1141), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(KEYINPUT118), .A3(new_n671), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1141), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT119), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(new_n1093), .C2(new_n1095), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1145), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1097), .B(new_n1122), .C1(new_n1144), .C2(new_n1150), .ZN(G378));
  INV_X1    g0951(.A(new_n1127), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1142), .A2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n849), .A2(new_n860), .A3(new_n834), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT38), .B1(new_n863), .B2(new_n865), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT101), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n861), .A2(new_n866), .A3(new_n867), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n832), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n871), .ZN(new_n1159));
  OAI211_X1 g0959(.A(G330), .B(new_n879), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n618), .A2(new_n422), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n410), .B2(new_n846), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n846), .A2(new_n410), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n618), .B2(new_n422), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  OR3_X1    g0965(.A1(new_n1162), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1160), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n872), .A2(G330), .A3(new_n1168), .A4(new_n879), .ZN(new_n1171));
  AND4_X1   g0971(.A1(new_n899), .A2(new_n1170), .A3(new_n898), .A4(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1170), .A2(new_n1171), .B1(new_n898), .B2(new_n899), .ZN(new_n1173));
  OAI211_X1 g0973(.A(KEYINPUT57), .B(new_n1153), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT122), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1153), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT57), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n900), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1170), .A2(new_n898), .A3(new_n1171), .A4(new_n899), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT122), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1182), .A2(new_n1183), .A3(KEYINPUT57), .A4(new_n1153), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1175), .A2(new_n1178), .A3(new_n671), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n750), .A2(G125), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n801), .A2(new_n1110), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n744), .A2(G150), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(G132), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n922), .A2(new_n1190), .B1(new_n754), .B2(new_n942), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1189), .B(new_n1191), .C1(G128), .C2(new_n805), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n279), .B(new_n305), .C1(new_n740), .C2(new_n269), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G124), .B2(new_n771), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n773), .A2(G58), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT121), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1031), .A2(new_n305), .A3(new_n258), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n758), .A2(new_n1068), .B1(new_n230), .B2(new_n761), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n936), .B(new_n1203), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n224), .B2(new_n922), .C1(new_n388), .C2(new_n754), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1202), .B(new_n1205), .C1(G116), .C2(new_n750), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G50), .B1(new_n279), .B2(new_n305), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n314), .B2(G41), .ZN(new_n1210));
  AND4_X1   g1010(.A1(new_n1198), .A2(new_n1207), .A3(new_n1208), .A4(new_n1210), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n720), .B1(G50), .B2(new_n1119), .C1(new_n1211), .C2(new_n918), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1169), .B2(new_n722), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1182), .B2(new_n958), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1185), .A2(new_n1214), .ZN(G375));
  AOI21_X1  g1015(.A(new_n719), .B1(new_n276), .B2(new_n816), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n756), .A2(G116), .B1(G294), .B2(new_n750), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n230), .B2(new_n754), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT124), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n314), .B1(new_n801), .B2(G97), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n1032), .C1(new_n740), .C2(new_n414), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n758), .A2(new_n571), .B1(new_n1068), .B2(new_n761), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n763), .A2(G137), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n922), .A2(new_n1109), .B1(new_n754), .B2(new_n1075), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n258), .B1(new_n801), .B2(G159), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1199), .B(new_n1226), .C1(new_n202), .C2(new_n932), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n758), .A2(new_n1107), .B1(new_n1190), .B2(new_n749), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1219), .A2(new_n1223), .B1(new_n1224), .B2(new_n1229), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1216), .B1(new_n918), .B2(new_n1230), .C1(new_n1134), .C2(new_n723), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n958), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT123), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT123), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1236), .A3(new_n958), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1232), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1135), .A2(new_n1140), .A3(new_n1127), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1147), .A2(new_n996), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(G381));
  NAND2_X1  g1041(.A1(new_n1097), .A2(new_n1122), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1144), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1150), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1185), .A2(new_n1245), .A3(new_n1214), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1018), .B(new_n1057), .C1(new_n721), .C2(new_n779), .ZN(new_n1247));
  OR3_X1    g1047(.A1(G390), .A2(G384), .A3(new_n1247), .ZN(new_n1248));
  OR4_X1    g1048(.A1(G387), .A2(new_n1246), .A3(G381), .A4(new_n1248), .ZN(G407));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G343), .C2(new_n1246), .ZN(G409));
  INV_X1    g1050(.A(G390), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1252), .A2(new_n1247), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G387), .B2(KEYINPUT126), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1247), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n995), .B1(new_n993), .B2(new_n713), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1012), .B(new_n1011), .C1(new_n1256), .C2(new_n958), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1255), .B1(new_n1257), .B2(new_n957), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1251), .B1(new_n1254), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G387), .A2(new_n1253), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT126), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1257), .B2(new_n957), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1260), .B(G390), .C1(new_n1262), .C2(new_n1253), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1259), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT127), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1264), .B(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1185), .A2(G378), .A3(new_n1214), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1214), .B1(new_n995), .B2(new_n1176), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1245), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n647), .A2(G213), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1239), .A2(KEYINPUT60), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1239), .A2(KEYINPUT60), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n671), .B(new_n1147), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1274), .A2(new_n1238), .A3(G384), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G384), .B1(new_n1274), .B2(new_n1238), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1270), .A2(new_n1271), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT125), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1270), .A2(KEYINPUT125), .A3(new_n1271), .A4(new_n1277), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT62), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n647), .A2(G213), .A3(G2897), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1277), .B(new_n1284), .Z(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT61), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1278), .A2(KEYINPUT62), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1266), .B1(new_n1282), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1280), .A2(new_n1290), .A3(new_n1281), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1278), .A2(new_n1290), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1286), .A4(new_n1264), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1289), .A2(new_n1293), .ZN(G405));
  OAI21_X1  g1094(.A(new_n1264), .B1(new_n1276), .B2(new_n1275), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1259), .A2(new_n1277), .A3(new_n1263), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(G375), .B(new_n1245), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1297), .B(new_n1298), .ZN(G402));
endmodule


