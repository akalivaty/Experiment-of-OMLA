//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G211gat), .B(G218gat), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n205));
  OR2_X1    g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT79), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n210));
  AOI211_X1 g009(.A(new_n210), .B(new_n205), .C1(new_n206), .C2(new_n207), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n204), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(KEYINPUT79), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT2), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G148gat), .ZN(new_n219));
  INV_X1    g018(.A(G148gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G141gat), .ZN(new_n221));
  OAI211_X1 g020(.A(KEYINPUT84), .B(new_n217), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G155gat), .B(G162gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G141gat), .B(G148gat), .Z(new_n226));
  NAND4_X1  g025(.A1(new_n226), .A2(KEYINPUT84), .A3(new_n223), .A4(new_n217), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT85), .B(KEYINPUT3), .Z(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT86), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT86), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n225), .A2(new_n227), .A3(new_n231), .A4(new_n228), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n215), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n225), .A2(new_n227), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n206), .A2(new_n207), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n210), .B1(new_n238), .B2(new_n205), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n203), .B1(new_n239), .B2(new_n213), .ZN(new_n240));
  INV_X1    g039(.A(new_n214), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n234), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n237), .B1(new_n242), .B2(new_n228), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n202), .B1(new_n235), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT29), .B1(new_n212), .B2(new_n214), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n236), .B1(new_n245), .B2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g045(.A(new_n202), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT29), .B1(new_n230), .B2(new_n232), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n246), .B(new_n247), .C1(new_n215), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT91), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n244), .A2(new_n249), .A3(KEYINPUT91), .ZN(new_n253));
  XNOR2_X1  g052(.A(G78gat), .B(G106gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT31), .B(G50gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  NAND3_X1  g055(.A1(new_n252), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT92), .B(G22gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n256), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n244), .A2(new_n249), .A3(KEYINPUT91), .A4(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n257), .B2(new_n260), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G225gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(G134gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G127gat), .ZN(new_n266));
  INV_X1    g065(.A(G127gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G134gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G113gat), .B(G120gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n269), .B1(new_n270), .B2(KEYINPUT1), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n266), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G120gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT69), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G120gat), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n275), .A2(new_n277), .A3(KEYINPUT70), .A4(G113gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(new_n274), .B2(G113gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT69), .B(G120gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(new_n282), .B2(G113gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n271), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n236), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n275), .A2(new_n277), .A3(G113gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n281), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n278), .A3(new_n273), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n289), .A2(new_n227), .A3(new_n225), .A4(new_n271), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n264), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n292));
  OR3_X1    g091(.A1(new_n291), .A2(KEYINPUT88), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT88), .B1(new_n291), .B2(new_n292), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n236), .A2(KEYINPUT3), .B1(new_n289), .B2(new_n271), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n233), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT4), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n289), .A2(KEYINPUT71), .A3(new_n271), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n301), .A2(KEYINPUT4), .A3(new_n237), .A4(new_n302), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n297), .A2(new_n264), .A3(new_n299), .A4(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT87), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n303), .A2(new_n299), .ZN(new_n307));
  INV_X1    g106(.A(new_n264), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(new_n233), .B2(new_n296), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT87), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n295), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n292), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n301), .A2(new_n237), .A3(new_n302), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n298), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n290), .A2(new_n298), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n311), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G1gat), .B(G29gat), .Z(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT0), .ZN(new_n322));
  XNOR2_X1  g121(.A(G57gat), .B(G85gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT6), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n304), .A2(new_n305), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n307), .A2(KEYINPUT87), .A3(new_n309), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n318), .B1(new_n331), .B2(new_n295), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(new_n324), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n329), .A2(new_n330), .B1(new_n294), .B2(new_n293), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n324), .B1(new_n312), .B2(new_n317), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT89), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT89), .ZN(new_n337));
  INV_X1    g136(.A(new_n335), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n311), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n336), .A2(new_n339), .A3(new_n327), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n333), .B1(new_n340), .B2(KEYINPUT90), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT90), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n336), .A2(new_n339), .A3(new_n342), .A4(new_n327), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n328), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G8gat), .B(G36gat), .Z(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT81), .ZN(new_n346));
  XNOR2_X1  g145(.A(G64gat), .B(G92gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n346), .B(new_n347), .Z(new_n348));
  INV_X1    g147(.A(new_n215), .ZN(new_n349));
  INV_X1    g148(.A(G226gat), .ZN(new_n350));
  INV_X1    g149(.A(G233gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n353));
  INV_X1    g152(.A(G183gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT27), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G183gat), .ZN(new_n357));
  INV_X1    g156(.A(G190gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n353), .B1(new_n359), .B2(KEYINPUT67), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT66), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT27), .B(G183gat), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(new_n358), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n360), .B1(new_n363), .B2(KEYINPUT67), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT67), .B1(new_n359), .B2(KEYINPUT66), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n353), .ZN(new_n366));
  NOR2_X1   g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT68), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n369), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT26), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n370), .A2(new_n372), .B1(G183gat), .B2(G190gat), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n364), .A2(new_n366), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n367), .A2(KEYINPUT23), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT23), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(G169gat), .B2(G176gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT65), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n375), .A2(new_n377), .A3(new_n378), .A4(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT24), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(G183gat), .A3(G190gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G183gat), .B(G190gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(new_n383), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n382), .B1(new_n386), .B2(KEYINPUT25), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n354), .A2(G190gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n358), .A2(G183gat), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n383), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n383), .A2(G183gat), .A3(G190gat), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT64), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n378), .B1(new_n367), .B2(KEYINPUT23), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n376), .A2(G169gat), .A3(G176gat), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n379), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT64), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n396), .B(new_n384), .C1(new_n385), .C2(new_n383), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n387), .B1(new_n398), .B2(new_n380), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n374), .A2(new_n399), .A3(KEYINPUT80), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n395), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n388), .A2(new_n389), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT24), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n396), .B1(new_n404), .B2(new_n384), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n380), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n387), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n364), .A2(new_n366), .A3(new_n373), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n401), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n352), .B1(new_n400), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n352), .A2(KEYINPUT29), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n412), .B1(new_n374), .B2(new_n399), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n349), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT80), .B1(new_n374), .B2(new_n399), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n391), .B1(new_n403), .B2(KEYINPUT24), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n416), .A2(new_n396), .B1(new_n417), .B2(new_n379), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT25), .B1(new_n418), .B2(new_n392), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n401), .B(new_n409), .C1(new_n419), .C2(new_n387), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n420), .A3(new_n412), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n374), .A2(new_n399), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n352), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n421), .A2(new_n349), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n348), .B1(new_n414), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n426));
  INV_X1    g225(.A(new_n352), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(new_n415), .B2(new_n420), .ZN(new_n428));
  INV_X1    g227(.A(new_n413), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n215), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n421), .A2(new_n349), .A3(new_n423), .ZN(new_n431));
  INV_X1    g230(.A(new_n348), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT30), .A4(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n425), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n430), .A2(new_n431), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n435), .A2(KEYINPUT82), .A3(KEYINPUT30), .A4(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(new_n436), .A3(KEYINPUT83), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n435), .A2(new_n432), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n263), .B1(new_n344), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n324), .B(KEYINPUT93), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n320), .A2(KEYINPUT96), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT96), .ZN(new_n448));
  INV_X1    g247(.A(new_n446), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n448), .B1(new_n332), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n336), .A2(new_n339), .A3(new_n327), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n328), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT37), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n430), .A2(new_n454), .A3(new_n431), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n349), .B1(new_n428), .B2(new_n429), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n421), .A2(new_n215), .A3(new_n423), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(KEYINPUT37), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n432), .A2(KEYINPUT38), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n441), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT37), .B1(new_n414), .B2(new_n424), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT97), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n348), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n454), .B1(new_n430), .B2(new_n431), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT97), .B1(new_n465), .B2(new_n432), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n466), .A3(new_n455), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n461), .B1(new_n467), .B2(KEYINPUT38), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n314), .A2(new_n297), .A3(new_n316), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n308), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT95), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n285), .A2(new_n264), .A3(new_n290), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT94), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n285), .A2(new_n290), .A3(KEYINPUT94), .A4(new_n264), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT39), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n472), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n473), .A2(new_n474), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(KEYINPUT95), .A3(KEYINPUT39), .A4(new_n476), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n471), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n315), .B1(new_n313), .B2(new_n298), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n264), .B1(new_n482), .B2(new_n297), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT39), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n446), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n481), .A2(new_n485), .A3(KEYINPUT40), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n450), .B2(new_n447), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n437), .A2(new_n443), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n263), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n469), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT72), .B1(new_n374), .B2(new_n399), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(new_n409), .C1(new_n419), .C2(new_n387), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n301), .A2(new_n302), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(G227gat), .A2(G233gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n422), .A2(new_n496), .A3(new_n498), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT32), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT33), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT73), .B(G71gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(G99gat), .ZN(new_n508));
  XOR2_X1   g307(.A(G15gat), .B(G43gat), .Z(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  NAND3_X1  g309(.A1(new_n504), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n510), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n503), .B(KEYINPUT32), .C1(new_n505), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT74), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n500), .A2(new_n502), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n515), .B(new_n516), .C1(new_n517), .C2(new_n501), .ZN(new_n518));
  INV_X1    g317(.A(new_n516), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n501), .B1(new_n500), .B2(new_n502), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT76), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n511), .A2(new_n518), .A3(new_n513), .A4(new_n521), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n514), .A2(new_n522), .A3(KEYINPUT76), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(KEYINPUT36), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n525), .B(KEYINPUT77), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n523), .A2(KEYINPUT78), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT78), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n522), .A3(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n529), .A2(new_n530), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  AND4_X1   g333(.A1(new_n445), .A2(new_n494), .A3(new_n528), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n340), .A2(KEYINPUT90), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(new_n326), .A3(new_n343), .ZN(new_n537));
  INV_X1    g336(.A(new_n328), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n263), .B1(new_n527), .B2(new_n526), .ZN(new_n540));
  INV_X1    g339(.A(new_n440), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT83), .B1(new_n434), .B2(new_n436), .ZN(new_n542));
  INV_X1    g341(.A(new_n443), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n529), .A2(new_n531), .A3(new_n533), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n257), .A2(new_n260), .ZN(new_n547));
  INV_X1    g346(.A(new_n258), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n551), .A2(new_n552), .A3(new_n437), .A4(new_n443), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(new_n453), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n545), .A2(KEYINPUT35), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n535), .A2(new_n555), .ZN(new_n556));
  OR3_X1    g355(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT99), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n557), .B2(new_n558), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n559), .A2(new_n562), .B1(G29gat), .B2(G36gat), .ZN(new_n563));
  XOR2_X1   g362(.A(G43gat), .B(G50gat), .Z(new_n564));
  INV_X1    g363(.A(KEYINPUT15), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n564), .A2(new_n565), .B1(new_n557), .B2(new_n560), .ZN(new_n568));
  NAND2_X1  g367(.A1(G29gat), .A2(G36gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT100), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT17), .ZN(new_n573));
  INV_X1    g372(.A(G8gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(G15gat), .B(G22gat), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n575), .A2(G1gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT101), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT16), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n575), .B1(new_n579), .B2(G1gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n578), .B(new_n581), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n571), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n573), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n572), .A2(new_n582), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT18), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n582), .B(new_n583), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n589), .B(KEYINPUT13), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n586), .A2(KEYINPUT18), .A3(new_n589), .A4(new_n587), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT102), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(KEYINPUT98), .B(KEYINPUT11), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT12), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n595), .A2(new_n598), .A3(new_n605), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n556), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(KEYINPUT105), .A2(G85gat), .A3(G92gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT7), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(G99gat), .A2(G106gat), .ZN(new_n615));
  INV_X1    g414(.A(G85gat), .ZN(new_n616));
  INV_X1    g415(.A(G92gat), .ZN(new_n617));
  AOI22_X1  g416(.A1(KEYINPUT8), .A2(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G99gat), .B(G106gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n573), .A2(new_n585), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT106), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n621), .ZN(new_n625));
  AND2_X1   g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n583), .A2(new_n625), .B1(KEYINPUT41), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n626), .A2(KEYINPUT41), .ZN(new_n631));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n630), .B(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT103), .ZN(new_n637));
  XOR2_X1   g436(.A(G57gat), .B(G64gat), .Z(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G71gat), .B(G78gat), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(G64gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(G57gat), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT104), .B(G57gat), .Z(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n642), .ZN(new_n645));
  INV_X1    g444(.A(new_n640), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n637), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT21), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n267), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n582), .B1(new_n649), .B2(new_n648), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G155gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G183gat), .B(G211gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n635), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(G230gat), .A2(G233gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n648), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n625), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n648), .B2(new_n621), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n666), .A2(new_n668), .A3(new_n625), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT10), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT10), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n665), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n665), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G120gat), .B(G148gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(G176gat), .B(G204gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n678), .B(new_n679), .Z(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n681), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n677), .A2(KEYINPUT108), .A3(new_n681), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n664), .A2(KEYINPUT109), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT109), .B1(new_n664), .B2(new_n687), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n610), .A2(new_n344), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  AND3_X1   g491(.A1(new_n610), .A2(new_n492), .A3(new_n690), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n574), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  AND4_X1   g494(.A1(new_n492), .A2(new_n610), .A3(new_n690), .A4(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT42), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n696), .A2(KEYINPUT42), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n697), .B2(new_n699), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(G1325gat));
  NAND2_X1  g501(.A1(new_n610), .A2(new_n690), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n534), .A2(new_n528), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G15gat), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n546), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n707), .A2(G15gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n703), .B2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT111), .Z(G1326gat));
  NOR2_X1   g509(.A1(new_n703), .A2(new_n551), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT43), .B(G22gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  INV_X1    g512(.A(new_n635), .ZN(new_n714));
  INV_X1    g513(.A(new_n687), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n714), .A2(new_n662), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n610), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n717), .A2(G29gat), .A3(new_n539), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT45), .Z(new_n719));
  OAI21_X1  g518(.A(new_n635), .B1(new_n535), .B2(new_n555), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n635), .C1(new_n535), .C2(new_n555), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n609), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n725), .A2(new_n715), .A3(new_n662), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n344), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G29gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n719), .A2(new_n729), .ZN(G1328gat));
  INV_X1    g529(.A(G36gat), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n610), .A2(new_n731), .A3(new_n492), .A4(new_n716), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT46), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n727), .B2(new_n492), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n733), .A2(new_n734), .ZN(G1329gat));
  NOR3_X1   g534(.A1(new_n717), .A2(G43gat), .A3(new_n707), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n727), .A2(new_n704), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(G43gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g538(.A1(new_n717), .A2(G50gat), .A3(new_n551), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n263), .A3(new_n726), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(G50gat), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g542(.A1(new_n556), .A2(new_n725), .A3(new_n664), .A4(new_n715), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n344), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(new_n644), .ZN(G1332gat));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n492), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT49), .B(G64gat), .Z(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1333gat));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n704), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n707), .A2(G71gat), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n751), .A2(G71gat), .B1(new_n744), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n744), .A2(new_n263), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NAND4_X1  g555(.A1(new_n556), .A2(new_n725), .A3(new_n663), .A4(new_n635), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n759), .A2(new_n616), .A3(new_n344), .A4(new_n715), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n609), .A2(new_n662), .A3(new_n687), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n722), .A2(new_n723), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT112), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n722), .A2(new_n764), .A3(new_n723), .A4(new_n761), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n344), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G85gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n760), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1336gat));
  AND3_X1   g569(.A1(new_n715), .A2(new_n617), .A3(new_n492), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT52), .B1(new_n759), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n762), .B1(new_n437), .B2(new_n443), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n617), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n763), .A2(new_n492), .A3(new_n765), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(KEYINPUT114), .A3(G92gat), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT114), .B1(new_n775), .B2(G92gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n757), .A2(KEYINPUT116), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n758), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n757), .A2(KEYINPUT116), .A3(KEYINPUT51), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n771), .B(KEYINPUT115), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n776), .A2(new_n777), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n774), .B1(new_n783), .B2(new_n784), .ZN(G1337gat));
  NAND3_X1  g584(.A1(new_n763), .A2(new_n704), .A3(new_n765), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G99gat), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n707), .A2(new_n687), .A3(G99gat), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT117), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n759), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1338gat));
  NOR3_X1   g590(.A1(new_n687), .A2(G106gat), .A3(new_n551), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n779), .A2(new_n780), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n779), .A2(KEYINPUT118), .A3(new_n780), .A4(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n763), .A2(new_n263), .A3(new_n765), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(G106gat), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT53), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n724), .A2(new_n263), .A3(new_n761), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT53), .B1(new_n801), .B2(G106gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n759), .A2(new_n792), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n803), .A2(KEYINPUT119), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(KEYINPUT119), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n800), .A2(new_n806), .ZN(G1339gat));
  NOR2_X1   g606(.A1(new_n588), .A2(new_n589), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n591), .A2(new_n593), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n604), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n608), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n676), .A2(new_n673), .ZN(new_n812));
  INV_X1    g611(.A(new_n665), .ZN(new_n813));
  INV_X1    g612(.A(new_n674), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(KEYINPUT54), .A3(new_n675), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n817), .B(new_n665), .C1(new_n672), .C2(new_n674), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT55), .A4(new_n681), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n682), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n682), .A2(new_n819), .A3(KEYINPUT120), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n816), .A2(new_n818), .A3(new_n681), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n822), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n635), .A2(new_n811), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n609), .A2(new_n823), .A3(new_n826), .A4(new_n822), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n715), .A2(new_n811), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n635), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n663), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n714), .A2(new_n662), .A3(new_n687), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n609), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n539), .A2(new_n492), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n835), .A2(new_n551), .A3(new_n546), .A4(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(G113gat), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n837), .A2(new_n838), .A3(new_n725), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n835), .A2(new_n836), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n540), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n609), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n839), .B1(new_n838), .B2(new_n842), .ZN(G1340gat));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n282), .A3(new_n715), .ZN(new_n844));
  OAI21_X1  g643(.A(G120gat), .B1(new_n837), .B2(new_n687), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1341gat));
  NAND3_X1  g645(.A1(new_n841), .A2(new_n267), .A3(new_n662), .ZN(new_n847));
  OAI21_X1  g646(.A(G127gat), .B1(new_n837), .B2(new_n663), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1342gat));
  NAND3_X1  g648(.A1(new_n841), .A2(new_n265), .A3(new_n635), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n837), .B2(new_n714), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n704), .A2(new_n551), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n218), .A3(new_n609), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n855), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n835), .A2(new_n263), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n705), .A2(new_n836), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n609), .A2(new_n826), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n831), .B1(new_n866), .B2(new_n820), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n714), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n662), .B1(new_n868), .B2(new_n828), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n834), .A2(new_n609), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n263), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n865), .B1(new_n871), .B2(KEYINPUT57), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n873), .B2(new_n725), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n859), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n861), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n874), .B(new_n859), .C1(new_n860), .C2(new_n855), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1344gat));
  NAND3_X1  g677(.A1(new_n858), .A2(new_n220), .A3(new_n715), .ZN(new_n879));
  INV_X1    g678(.A(new_n873), .ZN(new_n880));
  AOI211_X1 g679(.A(KEYINPUT59), .B(new_n220), .C1(new_n880), .C2(new_n715), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n688), .A2(new_n689), .A3(new_n609), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n863), .B(new_n263), .C1(new_n883), .C2(new_n869), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n865), .A2(new_n687), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n884), .B(new_n885), .C1(new_n862), .C2(new_n863), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n882), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n879), .B1(new_n881), .B2(new_n887), .ZN(G1345gat));
  NAND2_X1  g687(.A1(new_n662), .A2(G155gat), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT122), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(G155gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n857), .B2(new_n663), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n891), .A2(KEYINPUT123), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1346gat));
  AND3_X1   g697(.A1(new_n880), .A2(G162gat), .A3(new_n635), .ZN(new_n899));
  AOI21_X1  g698(.A(G162gat), .B1(new_n858), .B2(new_n635), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(G1347gat));
  NAND2_X1  g700(.A1(new_n539), .A2(new_n492), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n707), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n832), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n662), .B1(new_n904), .B2(new_n828), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n551), .B(new_n903), .C1(new_n905), .C2(new_n870), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT124), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n835), .A2(new_n908), .A3(new_n551), .A4(new_n903), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(G169gat), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n910), .A2(new_n911), .A3(new_n725), .ZN(new_n912));
  AND4_X1   g711(.A1(new_n539), .A2(new_n835), .A3(new_n492), .A4(new_n540), .ZN(new_n913));
  AOI21_X1  g712(.A(G169gat), .B1(new_n913), .B2(new_n609), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n912), .A2(new_n914), .ZN(G1348gat));
  OAI21_X1  g714(.A(G176gat), .B1(new_n910), .B2(new_n687), .ZN(new_n916));
  INV_X1    g715(.A(G176gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n913), .A2(new_n917), .A3(new_n715), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1349gat));
  NOR2_X1   g718(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n920));
  OAI21_X1  g719(.A(G183gat), .B1(new_n910), .B2(new_n663), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n913), .A2(new_n362), .A3(new_n662), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n923), .B(new_n924), .ZN(G1350gat));
  NAND3_X1  g724(.A1(new_n913), .A2(new_n358), .A3(new_n635), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n907), .A2(new_n909), .A3(new_n635), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n927), .A2(new_n928), .A3(G190gat), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n927), .B2(G190gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(KEYINPUT126), .B(new_n926), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1351gat));
  NOR2_X1   g734(.A1(new_n704), .A2(new_n902), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n862), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n937), .A2(new_n609), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n884), .B(new_n936), .C1(new_n862), .C2(new_n863), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n609), .A2(G197gat), .ZN(new_n940));
  OAI22_X1  g739(.A1(new_n938), .A2(G197gat), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(G1352gat));
  XOR2_X1   g741(.A(KEYINPUT127), .B(G204gat), .Z(new_n943));
  NAND3_X1  g742(.A1(new_n937), .A2(new_n715), .A3(new_n943), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n939), .A2(new_n687), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n945), .B(new_n946), .C1(new_n943), .C2(new_n947), .ZN(G1353gat));
  INV_X1    g747(.A(G211gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n937), .A2(new_n949), .A3(new_n662), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n939), .A2(new_n663), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT63), .B1(new_n951), .B2(G211gat), .ZN(new_n952));
  OAI211_X1 g751(.A(KEYINPUT63), .B(G211gat), .C1(new_n939), .C2(new_n663), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n950), .B1(new_n952), .B2(new_n954), .ZN(G1354gat));
  OAI21_X1  g754(.A(G218gat), .B1(new_n939), .B2(new_n714), .ZN(new_n956));
  INV_X1    g755(.A(G218gat), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n937), .A2(new_n957), .A3(new_n635), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1355gat));
endmodule


