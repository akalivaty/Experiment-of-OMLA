//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n578, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT71), .Z(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n462), .B1(new_n464), .B2(new_n460), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT69), .B1(new_n469), .B2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n468), .A2(new_n470), .A3(new_n460), .A4(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n465), .A2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(new_n473), .A2(KEYINPUT72), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(KEYINPUT72), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT3), .ZN(new_n485));
  AND2_X1   g060(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n486));
  AOI22_X1  g061(.A1(KEYINPUT69), .A2(new_n485), .B1(new_n486), .B2(new_n469), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n487), .A2(G2105), .A3(new_n468), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n483), .B1(new_n488), .B2(G124), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n480), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT4), .B1(new_n472), .B2(new_n492), .ZN(new_n493));
  XOR2_X1   g068(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n494));
  NAND4_X1  g069(.A1(new_n494), .A2(G138), .A3(new_n460), .A4(new_n463), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n468), .A2(new_n470), .A3(new_n471), .A4(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n503), .A2(new_n504), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n487), .A2(KEYINPUT73), .A3(new_n468), .A4(new_n502), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(new_n504), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n500), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT74), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n497), .B1(new_n509), .B2(new_n513), .ZN(G164));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT77), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n518), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G88), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n518), .A2(new_n521), .A3(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(new_n515), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT79), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n526), .A2(G89), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n538));
  INV_X1    g113(.A(new_n528), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n536), .B(new_n537), .C1(new_n541), .C2(KEYINPUT78), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n541), .A2(KEYINPUT78), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(G168));
  XNOR2_X1  g119(.A(KEYINPUT80), .B(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n526), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n528), .A2(G52), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n515), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(G171));
  NAND2_X1  g126(.A1(new_n526), .A2(G81), .ZN(new_n552));
  XOR2_X1   g127(.A(KEYINPUT81), .B(G43), .Z(new_n553));
  NAND2_X1  g128(.A1(new_n528), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n515), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT82), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(new_n524), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n525), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n539), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n528), .A2(new_n574), .A3(G53), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n571), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  XNOR2_X1  g152(.A(new_n550), .B(KEYINPUT83), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  NAND2_X1  g155(.A1(new_n526), .A2(G87), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n528), .A2(G49), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(new_n526), .A2(G86), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n528), .A2(G48), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n515), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n526), .A2(G85), .ZN(new_n590));
  XOR2_X1   g165(.A(KEYINPUT84), .B(G47), .Z(new_n591));
  NAND2_X1  g166(.A1(new_n528), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n515), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n590), .A2(new_n592), .A3(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(KEYINPUT85), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n526), .A2(G92), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n566), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n528), .A2(G54), .B1(G651), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(KEYINPUT86), .ZN(new_n608));
  AND3_X1   g183(.A1(new_n601), .A2(KEYINPUT86), .A3(new_n605), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n596), .A2(KEYINPUT85), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n598), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G284));
  XNOR2_X1  g189(.A(new_n613), .B(KEYINPUT87), .ZN(G321));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(G299), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G168), .B2(new_n616), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(G168), .B2(new_n616), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n610), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n557), .A2(new_n616), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n608), .A2(new_n609), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n622), .B1(new_n624), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g200(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n626));
  XNOR2_X1  g201(.A(G323), .B(new_n626), .ZN(G282));
  NOR2_X1   g202(.A1(new_n484), .A2(G2105), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n463), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  NAND2_X1  g206(.A1(KEYINPUT89), .A2(G2100), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n631), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(KEYINPUT89), .B2(G2100), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n633), .B1(new_n635), .B2(new_n632), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n479), .A2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n488), .A2(G123), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT90), .ZN(new_n639));
  OR2_X1    g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n640), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n637), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n642), .A2(G2096), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(G2096), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n636), .A2(new_n643), .A3(new_n644), .ZN(G156));
  XOR2_X1   g220(.A(G2443), .B(G2446), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT92), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2451), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT93), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2427), .B(G2430), .Z(new_n655));
  AOI21_X1  g230(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n650), .B(new_n657), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT91), .B(KEYINPUT16), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2454), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(G14), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n659), .ZN(G401));
  XOR2_X1   g239(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  INV_X1    g247(.A(new_n665), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n672), .B1(new_n668), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n682), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT20), .Z(new_n686));
  AOI211_X1 g261(.A(new_n684), .B(new_n686), .C1(new_n679), .C2(new_n683), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  OAI21_X1  g268(.A(KEYINPUT95), .B1(G95), .B2(G2105), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g270(.A1(KEYINPUT95), .A2(G95), .A3(G2105), .ZN(new_n696));
  OAI221_X1 g271(.A(G2104), .B1(G107), .B2(new_n460), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT96), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G119), .B2(new_n488), .ZN(new_n699));
  INV_X1    g274(.A(G131), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n478), .ZN(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n701), .S(G29), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT35), .B(G1991), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G24), .ZN(new_n705));
  XOR2_X1   g280(.A(G290), .B(KEYINPUT97), .Z(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G16), .ZN(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G6), .B(G305), .S(G16), .Z(new_n710));
  XOR2_X1   g285(.A(KEYINPUT32), .B(G1981), .Z(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  MUX2_X1   g287(.A(G23), .B(G288), .S(G16), .Z(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT33), .B(G1976), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n713), .B(new_n714), .Z(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1971), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n712), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n704), .B(new_n709), .C1(new_n721), .C2(KEYINPUT34), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(KEYINPUT34), .B2(new_n721), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT36), .ZN(new_n724));
  INV_X1    g299(.A(G34), .ZN(new_n725));
  AOI21_X1  g300(.A(G29), .B1(new_n725), .B2(KEYINPUT24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(KEYINPUT24), .B2(new_n725), .ZN(new_n727));
  INV_X1    g302(.A(G160), .ZN(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G2084), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  INV_X1    g308(.A(G28), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(KEYINPUT30), .ZN(new_n735));
  AOI21_X1  g310(.A(G29), .B1(new_n734), .B2(KEYINPUT30), .ZN(new_n736));
  OR2_X1    g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  NAND2_X1  g312(.A1(KEYINPUT31), .A2(G11), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n732), .A2(new_n733), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n558), .A2(new_n716), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n716), .B2(G19), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(G1341), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  NOR2_X1   g320(.A1(G171), .A2(new_n716), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G5), .B2(new_n716), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n740), .B(new_n744), .C1(new_n745), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n729), .A2(G33), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n479), .A2(G139), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT25), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n463), .A2(G127), .ZN(new_n753));
  INV_X1    g328(.A(G115), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(new_n484), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n752), .B1(new_n755), .B2(G2105), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n749), .B1(new_n757), .B2(new_n729), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(G2072), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n716), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1956), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n747), .A2(new_n745), .B1(new_n729), .B2(new_n642), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G1341), .B2(new_n743), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n748), .A2(new_n759), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G4), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n610), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1348), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n716), .A2(G21), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G168), .B2(new_n716), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(G1966), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n729), .A2(G26), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT28), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n479), .A2(G140), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n776));
  INV_X1    g351(.A(G116), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G2105), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n488), .B2(G128), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n774), .B1(new_n780), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2067), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n771), .A2(G1966), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n772), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n766), .A2(new_n769), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n729), .A2(G27), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G164), .B2(new_n729), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT99), .B(G2078), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n729), .A2(G35), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G162), .B2(new_n729), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT29), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n790), .B1(new_n793), .B2(G2090), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n729), .A2(G32), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n476), .A2(G141), .A3(new_n477), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT98), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n488), .A2(G129), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT26), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n801), .A2(new_n802), .B1(G105), .B2(new_n628), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n797), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n795), .B1(new_n807), .B2(new_n729), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT27), .Z(new_n809));
  AOI211_X1 g384(.A(new_n789), .B(new_n794), .C1(G1996), .C2(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(G1996), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n793), .A2(G2090), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT100), .Z(new_n813));
  NAND4_X1  g388(.A1(new_n785), .A2(new_n810), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n724), .A2(new_n814), .ZN(G311));
  INV_X1    g390(.A(G311), .ZN(G150));
  NAND2_X1  g391(.A1(new_n528), .A2(G55), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n526), .A2(G93), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n817), .B(new_n818), .C1(new_n515), .C2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT101), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT102), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n558), .B1(new_n820), .B2(new_n821), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n822), .B1(new_n820), .B2(new_n821), .ZN(new_n825));
  OR3_X1    g400(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n824), .B1(new_n823), .B2(new_n825), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n610), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n832));
  AOI21_X1  g407(.A(G860), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n832), .B2(new_n831), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n820), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n838));
  INV_X1    g413(.A(new_n780), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n797), .B2(new_n805), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n797), .A3(new_n805), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n512), .A2(new_n496), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n843), .ZN(new_n845));
  INV_X1    g420(.A(new_n842), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n840), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n757), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n844), .A2(new_n847), .A3(new_n757), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n701), .B(new_n630), .ZN(new_n853));
  INV_X1    g428(.A(G118), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(KEYINPUT103), .A3(G2105), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT103), .B1(new_n854), .B2(G2105), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n488), .A2(G130), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G142), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n478), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n853), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n838), .B1(new_n852), .B2(new_n863), .ZN(new_n864));
  AOI211_X1 g439(.A(KEYINPUT104), .B(new_n862), .C1(new_n850), .C2(new_n851), .ZN(new_n865));
  OAI22_X1  g440(.A1(new_n864), .A2(new_n865), .B1(new_n863), .B2(new_n852), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n490), .B(new_n728), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n642), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n852), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n868), .B1(new_n870), .B2(new_n862), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n852), .A2(new_n863), .ZN(new_n872));
  AOI21_X1  g447(.A(G37), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(KEYINPUT40), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT40), .B1(new_n869), .B2(new_n873), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(G395));
  NAND4_X1  g452(.A1(new_n610), .A2(new_n620), .A3(new_n826), .A4(new_n827), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n828), .B1(new_n623), .B2(G559), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  NAND2_X1  g456(.A1(G299), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n576), .A2(KEYINPUT105), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n607), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n606), .A2(new_n881), .A3(G299), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT106), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(KEYINPUT41), .A3(new_n885), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT41), .B1(new_n884), .B2(new_n885), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n878), .B(new_n879), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT42), .ZN(new_n894));
  XOR2_X1   g469(.A(G303), .B(G288), .Z(new_n895));
  XOR2_X1   g470(.A(G290), .B(G305), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n888), .A2(new_n899), .A3(new_n892), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n894), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n898), .B1(new_n894), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g477(.A(G868), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n820), .A2(new_n616), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(G295));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n904), .ZN(G331));
  XOR2_X1   g481(.A(new_n886), .B(KEYINPUT106), .Z(new_n907));
  NAND2_X1  g482(.A1(G168), .A2(new_n578), .ZN(new_n908));
  NAND2_X1  g483(.A1(G286), .A2(new_n550), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n828), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n908), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n826), .A3(new_n827), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n891), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n910), .A2(new_n912), .A3(new_n914), .A4(new_n889), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n907), .A2(new_n913), .B1(new_n915), .B2(KEYINPUT107), .ZN(new_n916));
  INV_X1    g491(.A(new_n913), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n890), .A2(new_n891), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n897), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n915), .B1(new_n917), .B2(new_n886), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n922), .B1(new_n923), .B2(new_n898), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n886), .B1(new_n910), .B2(new_n912), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n917), .B2(new_n918), .ZN(new_n928));
  AOI21_X1  g503(.A(G37), .B1(new_n928), .B2(new_n897), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n923), .A2(new_n898), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT43), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n921), .A2(new_n924), .A3(KEYINPUT43), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n925), .B1(new_n929), .B2(new_n930), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n936), .ZN(G397));
  NAND2_X1  g512(.A1(G303), .A2(G8), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  INV_X1    g514(.A(G1971), .ZN(new_n940));
  XOR2_X1   g515(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(G164), .B2(G1384), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n474), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n464), .A2(new_n460), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n944), .A2(new_n945), .A3(G40), .A4(new_n462), .ZN(new_n946));
  AOI21_X1  g521(.A(G1384), .B1(new_n512), .B2(new_n496), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT45), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n948), .B2(KEYINPUT112), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n950), .A3(KEYINPUT45), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n940), .B1(new_n943), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n510), .A2(new_n511), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT74), .B1(new_n954), .B2(new_n501), .ZN(new_n955));
  AOI211_X1 g530(.A(new_n508), .B(new_n500), .C1(new_n510), .C2(new_n511), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n496), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n843), .A2(new_n959), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n946), .B1(new_n961), .B2(KEYINPUT50), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n963), .A2(G2090), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n953), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G8), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n939), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI211_X1 g542(.A(KEYINPUT113), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n968));
  INV_X1    g543(.A(G40), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n465), .A2(new_n474), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n958), .B1(new_n957), .B2(new_n959), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n947), .B2(new_n958), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n968), .B(new_n970), .C1(new_n971), .C2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT124), .B(G1961), .ZN(new_n975));
  INV_X1    g550(.A(G2078), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n942), .A2(new_n976), .A3(new_n949), .A4(new_n951), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n974), .A2(new_n975), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n970), .B1(new_n947), .B2(KEYINPUT45), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n941), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n957), .A2(new_n959), .A3(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n970), .B(KEYINPUT116), .C1(new_n947), .C2(KEYINPUT45), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  OR3_X1    g561(.A1(new_n986), .A2(new_n978), .A3(G2078), .ZN(new_n987));
  AOI21_X1  g562(.A(G301), .B1(new_n979), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n953), .B1(new_n974), .B2(G2090), .ZN(new_n989));
  INV_X1    g564(.A(new_n939), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(G8), .A3(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(G305), .A2(G1981), .ZN(new_n992));
  NAND2_X1  g567(.A1(G305), .A2(G1981), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n961), .A2(new_n946), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(new_n966), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n992), .A2(KEYINPUT49), .A3(new_n993), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1976), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n998), .B1(new_n1001), .B2(G288), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT52), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT52), .B1(G288), .B2(new_n1001), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n998), .B(new_n1004), .C1(new_n1001), .C2(G288), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1000), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AND4_X1   g581(.A1(new_n967), .A2(new_n988), .A3(new_n991), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT126), .ZN(new_n1008));
  INV_X1    g583(.A(new_n973), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n509), .A2(new_n513), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1384), .B1(new_n1010), .B2(new_n496), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1011), .B2(new_n958), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1012), .A2(new_n731), .A3(new_n970), .A4(new_n968), .ZN(new_n1013));
  INV_X1    g588(.A(G1966), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n986), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n966), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT123), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(G168), .B2(new_n966), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT123), .B(G8), .C1(new_n542), .C2(new_n543), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1016), .A2(KEYINPUT51), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1015), .B1(new_n974), .B2(G2084), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1020), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n1022), .B2(new_n1020), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1021), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1007), .B(new_n1008), .C1(new_n1028), .C2(KEYINPUT62), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1022), .A2(new_n1020), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(KEYINPUT51), .C1(new_n1020), .C2(new_n1016), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1023), .A2(new_n1026), .A3(new_n1024), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT62), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n967), .A2(new_n991), .A3(new_n1006), .A4(new_n988), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT126), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1029), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT63), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n967), .A2(new_n991), .A3(new_n1006), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1016), .A2(G168), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n991), .A2(new_n1006), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1040), .A2(new_n1038), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n989), .A2(G8), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1042), .B(new_n1043), .C1(new_n990), .C2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1006), .A2(G8), .A3(new_n990), .A4(new_n989), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G288), .A2(G1976), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT114), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1000), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n992), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n998), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1046), .A2(KEYINPUT115), .A3(new_n1051), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n1041), .A2(new_n1045), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n576), .A2(KEYINPUT57), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n573), .A2(new_n575), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n571), .A2(KEYINPUT119), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n571), .A2(KEYINPUT119), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1062));
  OAI21_X1  g637(.A(new_n1057), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT56), .B(G2072), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n942), .A2(new_n951), .A3(new_n949), .A4(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n1066));
  INV_X1    g641(.A(G1956), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n963), .B2(new_n1067), .ZN(new_n1068));
  AOI211_X1 g643(.A(KEYINPUT117), .B(G1956), .C1(new_n960), .C2(new_n962), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1063), .B(new_n1065), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n997), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(G2067), .ZN(new_n1073));
  INV_X1    g648(.A(G1348), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n974), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  AOI211_X1 g653(.A(KEYINPUT120), .B(new_n1073), .C1(new_n974), .C2(new_n1074), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n610), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n970), .B1(new_n947), .B2(new_n958), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n1011), .B2(new_n958), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT117), .B1(new_n1083), .B2(G1956), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n963), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1063), .B1(new_n1086), .B2(new_n1065), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1071), .B1(new_n1081), .B2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1090));
  INV_X1    g665(.A(G1996), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n942), .A2(new_n1091), .A3(new_n949), .A4(new_n951), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT58), .B(G1341), .Z(new_n1093));
  NAND2_X1  g668(.A1(new_n1072), .A2(new_n1093), .ZN(new_n1094));
  AOI211_X1 g669(.A(new_n557), .B(new_n1090), .C1(new_n1092), .C2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1096));
  XOR2_X1   g671(.A(new_n1095), .B(new_n1096), .Z(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT122), .B1(new_n1087), .B2(new_n1071), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT61), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(KEYINPUT122), .B(KEYINPUT61), .C1(new_n1087), .C2(new_n1071), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT60), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n623), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT60), .B(new_n610), .C1(new_n1077), .C2(new_n1079), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1104), .B(new_n1105), .C1(KEYINPUT60), .C2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1089), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n961), .A2(new_n941), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(KEYINPUT53), .A3(new_n976), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n979), .B1(new_n952), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1109), .B1(new_n1112), .B2(G171), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n979), .A2(G301), .A3(new_n987), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1113), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1112), .A2(new_n578), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1109), .B1(new_n1119), .B2(new_n988), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1039), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .A4(new_n1028), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1037), .B(new_n1056), .C1(new_n1108), .C2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1110), .A2(new_n946), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n807), .A2(new_n1091), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n780), .B(G2067), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1124), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1124), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(G1996), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n807), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1130), .A2(KEYINPUT110), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(KEYINPUT110), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1127), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT111), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n701), .B(new_n703), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(G290), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n708), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1138), .B(KEYINPUT109), .Z(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n708), .B2(new_n1137), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1136), .B1(new_n1124), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1123), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1124), .B1(new_n1126), .B2(new_n806), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1129), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1145), .A2(KEYINPUT46), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(KEYINPUT46), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1144), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT47), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1139), .A2(new_n1124), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT48), .Z(new_n1151));
  OAI21_X1  g726(.A(new_n1149), .B1(new_n1136), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n703), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n701), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1134), .A2(new_n1154), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n780), .A2(G2067), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1128), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1143), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g734(.A1(new_n907), .A2(new_n913), .ZN(new_n1161));
  NAND2_X1  g735(.A1(new_n915), .A2(KEYINPUT107), .ZN(new_n1162));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n1163), .A2(new_n898), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n1164), .A2(new_n929), .A3(new_n925), .ZN(new_n1165));
  INV_X1    g739(.A(new_n930), .ZN(new_n1166));
  OAI21_X1  g740(.A(KEYINPUT43), .B1(new_n1166), .B2(new_n924), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g742(.A1(new_n869), .A2(new_n873), .ZN(new_n1169));
  INV_X1    g743(.A(G319), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n1170), .A2(G227), .ZN(new_n1171));
  XNOR2_X1  g745(.A(new_n1171), .B(KEYINPUT127), .ZN(new_n1172));
  NOR3_X1   g746(.A1(G229), .A2(G401), .A3(new_n1172), .ZN(new_n1173));
  AND3_X1   g747(.A1(new_n1168), .A2(new_n1169), .A3(new_n1173), .ZN(G308));
  NAND3_X1  g748(.A1(new_n1168), .A2(new_n1169), .A3(new_n1173), .ZN(G225));
endmodule


