//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT17), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT91), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT91), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT14), .ZN(new_n208));
  NAND2_X1  g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n208), .B(new_n209), .C1(KEYINPUT14), .C2(new_n207), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n210), .A2(new_n211), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n214), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OAI211_X1 g017(.A(KEYINPUT92), .B(new_n202), .C1(new_n216), .C2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n210), .B(new_n211), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n213), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n202), .A2(KEYINPUT92), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n202), .A2(KEYINPUT92), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n221), .A2(new_n215), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT98), .B(G85gat), .Z(new_n226));
  INV_X1    g025(.A(G92gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G85gat), .A2(G92gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT7), .ZN(new_n230));
  INV_X1    g029(.A(G99gat), .ZN(new_n231));
  INV_X1    g030(.A(G106gat), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT8), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n228), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G99gat), .B(G106gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n234), .B(new_n235), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n225), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n215), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(new_n236), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(G190gat), .B(G218gat), .Z(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n237), .A2(new_n243), .A3(new_n240), .A4(new_n241), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G134gat), .B(G162gat), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n236), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n219), .B2(new_n224), .ZN(new_n252));
  INV_X1    g051(.A(new_n241), .ZN(new_n253));
  NOR4_X1   g052(.A1(new_n252), .A2(new_n244), .A3(new_n239), .A4(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n250), .B1(new_n254), .B2(KEYINPUT99), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n245), .A2(KEYINPUT99), .A3(new_n246), .A4(new_n250), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G15gat), .B(G22gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT16), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n259), .B1(new_n260), .B2(G1gat), .ZN(new_n261));
  INV_X1    g060(.A(G8gat), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n262), .A2(KEYINPUT93), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n261), .B(new_n263), .C1(G1gat), .C2(new_n259), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(KEYINPUT93), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G64gat), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n267), .A2(G57gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT96), .B(G57gat), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n268), .B1(new_n269), .B2(G64gat), .ZN(new_n270));
  AND2_X1   g069(.A1(G71gat), .A2(G78gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(G71gat), .A2(G78gat), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n271), .B1(KEYINPUT9), .B2(new_n272), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n267), .A2(G57gat), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT9), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n271), .A2(new_n272), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n266), .B1(KEYINPUT21), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT97), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT19), .ZN(new_n283));
  XNOR2_X1  g082(.A(G127gat), .B(G155gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT20), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n283), .B(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n280), .A2(KEYINPUT21), .ZN(new_n287));
  XNOR2_X1  g086(.A(G183gat), .B(G211gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(G231gat), .A2(G233gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n287), .B(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n286), .B(new_n291), .Z(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G227gat), .ZN(new_n294));
  INV_X1    g093(.A(G233gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G183gat), .ZN(new_n298));
  OR3_X1    g097(.A1(new_n298), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT27), .B1(new_n298), .B2(KEYINPUT66), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT27), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(G183gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n298), .A2(KEYINPUT27), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT67), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n298), .A2(KEYINPUT27), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT67), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(G190gat), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n303), .B1(new_n312), .B2(new_n300), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT68), .ZN(new_n314));
  NOR2_X1   g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n317), .A2(KEYINPUT26), .ZN(new_n318));
  NAND2_X1  g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n320), .B1(new_n317), .B2(KEYINPUT26), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n318), .A2(new_n321), .B1(G183gat), .B2(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n323), .B(new_n303), .C1(new_n312), .C2(new_n300), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n314), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n326));
  INV_X1    g125(.A(G134gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(G127gat), .ZN(new_n328));
  INV_X1    g127(.A(G127gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(G134gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n326), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G113gat), .B(G120gat), .Z(new_n332));
  XOR2_X1   g131(.A(KEYINPUT72), .B(KEYINPUT1), .Z(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(G134gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n327), .A2(G127gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT71), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n331), .A2(new_n332), .A3(new_n333), .A4(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT70), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n328), .A2(KEYINPUT70), .ZN(new_n340));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n339), .B(new_n340), .C1(KEYINPUT1), .C2(new_n341), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n337), .A2(KEYINPUT73), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT73), .B1(new_n337), .B2(new_n342), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT64), .B1(new_n315), .B2(KEYINPUT23), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n315), .A2(KEYINPUT23), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT64), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n348), .B(new_n349), .C1(G169gat), .C2(G176gat), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n346), .A2(new_n319), .A3(new_n347), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(KEYINPUT24), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n298), .A2(new_n301), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(KEYINPUT24), .A3(new_n352), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n351), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT25), .B1(new_n351), .B2(KEYINPUT65), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n320), .B1(KEYINPUT23), .B2(new_n315), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT65), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n360), .A2(new_n361), .A3(new_n346), .A4(new_n350), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n360), .A2(new_n355), .A3(new_n346), .A4(new_n350), .ZN(new_n363));
  OAI211_X1 g162(.A(KEYINPUT25), .B(new_n362), .C1(new_n363), .C2(new_n353), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n325), .A2(new_n345), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n345), .B1(new_n325), .B2(new_n365), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n297), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT77), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n370), .B(new_n297), .C1(new_n366), .C2(new_n367), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT34), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  OR3_X1    g172(.A1(new_n368), .A2(KEYINPUT77), .A3(new_n372), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n325), .A2(new_n365), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n337), .A2(new_n342), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT73), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n337), .A2(KEYINPUT73), .A3(new_n342), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n325), .A2(new_n345), .A3(new_n365), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n296), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT74), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n383), .A2(new_n387), .A3(new_n296), .A4(new_n384), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G15gat), .B(G43gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(G71gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(G99gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT75), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT75), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT32), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n376), .B1(new_n389), .B2(new_n400), .ZN(new_n401));
  AOI211_X1 g200(.A(KEYINPUT76), .B(new_n399), .C1(new_n386), .C2(new_n388), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n366), .A2(new_n367), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n387), .B1(new_n404), .B2(new_n296), .ZN(new_n405));
  INV_X1    g204(.A(new_n388), .ZN(new_n406));
  OAI22_X1  g205(.A1(new_n405), .A2(new_n406), .B1(KEYINPUT32), .B2(new_n395), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n393), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n375), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n400), .B1(new_n405), .B2(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT76), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n376), .A3(new_n400), .ZN(new_n412));
  AND4_X1   g211(.A1(new_n408), .A2(new_n375), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT36), .ZN(new_n415));
  INV_X1    g214(.A(G148gat), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT83), .B1(new_n416), .B2(G141gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n418));
  INV_X1    g217(.A(G141gat), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(new_n419), .A3(G148gat), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n417), .B(new_n420), .C1(new_n419), .C2(G148gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422));
  INV_X1    g221(.A(G155gat), .ZN(new_n423));
  INV_X1    g222(.A(G162gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n422), .B1(new_n425), .B2(KEYINPUT2), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  AND2_X1   g226(.A1(G155gat), .A2(G162gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT82), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT82), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n425), .A2(new_n431), .A3(new_n422), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n422), .A2(KEYINPUT2), .ZN(new_n433));
  XNOR2_X1  g232(.A(G141gat), .B(G148gat), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n430), .B(new_n432), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n427), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT3), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n427), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n378), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n337), .A2(new_n427), .A3(new_n435), .A4(new_n342), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT4), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n436), .B1(new_n380), .B2(new_n381), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n440), .B(new_n443), .C1(new_n444), .C2(KEYINPUT4), .ZN(new_n445));
  NAND2_X1  g244(.A1(G225gat), .A2(G233gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n445), .A2(KEYINPUT5), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n440), .A2(new_n446), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n337), .A2(new_n342), .ZN(new_n451));
  INV_X1    g250(.A(new_n436), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT84), .B1(new_n441), .B2(KEYINPUT4), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT4), .B1(new_n345), .B2(new_n436), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n450), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n342), .A2(new_n337), .B1(new_n427), .B2(new_n435), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n447), .B1(new_n442), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT5), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n449), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n440), .A2(new_n446), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n454), .B1(new_n382), .B2(new_n452), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n455), .A2(new_n456), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n462), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(KEYINPUT85), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n448), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G1gat), .B(G29gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(KEYINPUT0), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(G57gat), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n473), .B(G85gat), .Z(new_n474));
  AOI21_X1  g273(.A(KEYINPUT6), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n448), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n456), .B(new_n455), .C1(new_n444), .C2(new_n454), .ZN(new_n477));
  AOI211_X1 g276(.A(new_n449), .B(new_n462), .C1(new_n477), .C2(new_n464), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT85), .B1(new_n467), .B2(new_n468), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n474), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(KEYINPUT6), .A3(new_n481), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G197gat), .B(G204gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT22), .ZN(new_n487));
  INV_X1    g286(.A(G211gat), .ZN(new_n488));
  INV_X1    g287(.A(G218gat), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G211gat), .B(G218gat), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n486), .A3(new_n490), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT78), .ZN(new_n497));
  NAND2_X1  g296(.A1(G226gat), .A2(G233gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT79), .B(KEYINPUT29), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n377), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n325), .B2(new_n365), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n377), .A2(new_n499), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT29), .B1(new_n325), .B2(new_n365), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n505), .B(new_n496), .C1(new_n499), .C2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G8gat), .B(G36gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(new_n267), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(new_n227), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n504), .A2(new_n507), .A3(new_n512), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT81), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n504), .A2(KEYINPUT81), .A3(new_n507), .A4(new_n512), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n504), .A2(KEYINPUT30), .A3(new_n507), .A4(new_n512), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n521), .B(KEYINPUT80), .Z(new_n522));
  NAND3_X1  g321(.A1(new_n485), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT86), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n494), .A2(new_n495), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT78), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n439), .A2(new_n501), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n438), .B1(new_n525), .B2(KEYINPUT29), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n436), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n497), .A2(KEYINPUT86), .A3(new_n527), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(G228gat), .A2(G233gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G228gat), .A2(G233gat), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT3), .B1(new_n496), .B2(new_n501), .ZN(new_n537));
  OAI221_X1 g336(.A(new_n536), .B1(new_n537), .B2(new_n452), .C1(new_n528), .C2(new_n496), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT31), .B(G50gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n540), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n535), .A2(new_n542), .A3(new_n538), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G78gat), .B(G106gat), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(G22gat), .Z(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(new_n546), .A3(new_n543), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n523), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n409), .B2(new_n413), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n415), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n470), .A2(KEYINPUT87), .A3(new_n474), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT87), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n480), .B2(new_n481), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n475), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n480), .A2(KEYINPUT6), .A3(new_n481), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n504), .A2(new_n561), .A3(new_n507), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n562), .A2(new_n511), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT29), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n499), .B1(new_n377), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n525), .B1(new_n565), .B2(new_n503), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n500), .B1(new_n325), .B2(new_n365), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n505), .B(new_n526), .C1(new_n499), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT38), .B1(new_n569), .B2(KEYINPUT37), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n563), .A2(new_n570), .B1(new_n516), .B2(new_n517), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n559), .A2(new_n560), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT88), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n563), .B1(new_n561), .B2(new_n508), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT38), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT88), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n559), .A2(new_n571), .A3(new_n576), .A4(new_n560), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n445), .A2(new_n447), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n442), .A2(new_n460), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n579), .B(KEYINPUT39), .C1(new_n447), .C2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n581), .B(new_n474), .C1(KEYINPUT39), .C2(new_n579), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT40), .Z(new_n583));
  NOR2_X1   g382(.A1(new_n556), .A2(new_n558), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n520), .A2(new_n522), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n550), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n578), .A2(KEYINPUT89), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT89), .B1(new_n578), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n555), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n408), .A2(new_n411), .A3(new_n412), .ZN(new_n591));
  INV_X1    g390(.A(new_n375), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n403), .A2(new_n408), .A3(new_n375), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n550), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n586), .A2(KEYINPUT35), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n559), .A2(new_n560), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n599));
  INV_X1    g398(.A(new_n523), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI211_X1 g402(.A(new_n258), .B(new_n293), .C1(new_n590), .C2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n221), .A2(new_n215), .A3(new_n266), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n266), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n225), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT18), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n266), .B1(new_n219), .B2(new_n224), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT18), .ZN(new_n612));
  INV_X1    g411(.A(new_n609), .ZN(new_n613));
  NOR4_X1   g412(.A1(new_n611), .A2(new_n612), .A3(new_n606), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n238), .A2(new_n607), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT94), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n616), .A3(new_n605), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n609), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n238), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(KEYINPUT94), .A3(new_n266), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n610), .A2(new_n614), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(KEYINPUT90), .B(G197gat), .Z(new_n625));
  XNOR2_X1  g424(.A(G113gat), .B(G141gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT11), .B(G169gat), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  INV_X1    g429(.A(KEYINPUT95), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n630), .B1(new_n610), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n225), .A2(new_n607), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n609), .A3(new_n605), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n612), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n634), .B1(new_n637), .B2(KEYINPUT95), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n608), .A2(KEYINPUT18), .A3(new_n609), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n622), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n228), .A2(new_n233), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n235), .B1(new_n644), .B2(new_n230), .ZN(new_n645));
  AND4_X1   g444(.A1(new_n235), .A2(new_n228), .A3(new_n230), .A4(new_n233), .ZN(new_n646));
  OAI22_X1  g445(.A1(new_n645), .A2(new_n646), .B1(new_n279), .B2(KEYINPUT100), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  INV_X1    g447(.A(new_n278), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n270), .A2(new_n273), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT100), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n274), .B2(new_n278), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n647), .B(new_n648), .C1(new_n654), .C2(new_n236), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n279), .A2(new_n648), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n251), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(G230gat), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n295), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  MUX2_X1   g461(.A(new_n654), .B(new_n651), .S(new_n236), .Z(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G120gat), .B(G148gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT101), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G176gat), .ZN(new_n667));
  INV_X1    g466(.A(G204gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n664), .B(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n643), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n604), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n485), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT102), .B(G1gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1324gat));
  INV_X1    g474(.A(new_n672), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n262), .B1(new_n676), .B2(new_n586), .ZN(new_n677));
  INV_X1    g476(.A(new_n586), .ZN(new_n678));
  NOR2_X1   g477(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n260), .A2(new_n262), .ZN(new_n680));
  NOR4_X1   g479(.A1(new_n672), .A2(new_n678), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT42), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(KEYINPUT42), .B2(new_n681), .ZN(G1325gat));
  NAND2_X1  g482(.A1(new_n415), .A2(new_n553), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n676), .A2(G15gat), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n414), .ZN(new_n686));
  AOI21_X1  g485(.A(G15gat), .B1(new_n676), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n685), .A2(new_n687), .ZN(G1326gat));
  NAND2_X1  g487(.A1(new_n548), .A2(new_n549), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n672), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  INV_X1    g491(.A(new_n258), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n693), .B1(new_n590), .B2(new_n603), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n292), .A2(new_n670), .A3(new_n643), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n483), .A2(new_n484), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n203), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n578), .A2(new_n587), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT89), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n578), .A2(KEYINPUT89), .A3(new_n587), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n554), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g503(.A(KEYINPUT44), .B(new_n258), .C1(new_n704), .C2(new_n602), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT103), .B1(new_n598), .B2(new_n601), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n689), .B1(new_n409), .B2(new_n413), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT35), .B1(new_n707), .B2(new_n523), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n693), .B1(new_n590), .B2(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n705), .B(new_n695), .C1(KEYINPUT44), .C2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G29gat), .B1(new_n714), .B2(new_n485), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n715), .ZN(G1328gat));
  NAND3_X1  g515(.A1(new_n696), .A2(new_n204), .A3(new_n586), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT46), .Z(new_n718));
  OAI21_X1  g517(.A(G36gat), .B1(new_n714), .B2(new_n678), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(G1329gat));
  INV_X1    g519(.A(new_n684), .ZN(new_n721));
  OAI21_X1  g520(.A(G43gat), .B1(new_n714), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(G43gat), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n696), .A2(new_n723), .A3(new_n686), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g525(.A(G50gat), .B1(new_n714), .B2(new_n689), .ZN(new_n727));
  INV_X1    g526(.A(G50gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n696), .A2(new_n728), .A3(new_n550), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n733), .B2(KEYINPUT48), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735));
  AOI211_X1 g534(.A(KEYINPUT105), .B(new_n735), .C1(new_n727), .C2(new_n732), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n730), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n733), .A2(new_n731), .A3(KEYINPUT48), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n702), .A2(new_n703), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n740), .A2(new_n555), .B1(new_n706), .B2(new_n711), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n741), .B2(new_n693), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n742), .A2(new_n550), .A3(new_n695), .A4(new_n705), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT104), .B1(new_n743), .B2(G50gat), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT105), .B1(new_n744), .B2(new_n735), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n738), .A2(new_n745), .A3(new_n727), .A4(new_n729), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n737), .A2(new_n746), .ZN(G1331gat));
  INV_X1    g546(.A(new_n670), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n292), .A2(new_n643), .A3(new_n693), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n741), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n697), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(new_n269), .Z(G1332gat));
  NAND2_X1  g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n750), .A2(new_n586), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT106), .Z(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1333gat));
  NAND2_X1  g556(.A1(new_n750), .A2(new_n684), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n414), .A2(G71gat), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n758), .A2(G71gat), .B1(new_n750), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n750), .A2(new_n550), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g562(.A1(new_n590), .A2(new_n712), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT44), .B1(new_n764), .B2(new_n258), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(KEYINPUT44), .B2(new_n694), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n485), .A2(new_n748), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n292), .A2(new_n642), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT98), .B(G85gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n708), .A2(new_n710), .A3(new_n709), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n710), .B1(new_n708), .B2(new_n709), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n258), .B(new_n768), .C1(new_n704), .C2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n764), .A2(KEYINPUT51), .A3(new_n258), .A4(new_n768), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n779), .A2(new_n778), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n780), .A2(new_n781), .A3(new_n226), .A4(new_n767), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n771), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(G1336gat));
  NAND4_X1  g584(.A1(new_n742), .A2(new_n670), .A3(new_n705), .A4(new_n768), .ZN(new_n786));
  OAI21_X1  g585(.A(G92gat), .B1(new_n786), .B2(new_n678), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n678), .A2(G92gat), .A3(new_n748), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n780), .A2(new_n781), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n788), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n777), .B2(new_n779), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n787), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT109), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n766), .A2(new_n670), .A3(new_n586), .A4(new_n768), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n793), .B1(new_n799), .B2(G92gat), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n797), .B(new_n798), .C1(new_n800), .C2(new_n790), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(G1337gat));
  OAI21_X1  g601(.A(G99gat), .B1(new_n786), .B2(new_n721), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n780), .A2(new_n781), .A3(new_n231), .A4(new_n686), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(new_n748), .ZN(G1338gat));
  OAI21_X1  g604(.A(G106gat), .B1(new_n786), .B2(new_n689), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n689), .A2(new_n748), .A3(G106gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n780), .A2(new_n781), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n777), .A2(new_n779), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n807), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n813), .B2(new_n809), .ZN(G1339gat));
  INV_X1    g613(.A(new_n669), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n655), .A2(new_n660), .A3(new_n657), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n662), .A2(KEYINPUT54), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n817), .B2(KEYINPUT110), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n662), .A2(KEYINPUT54), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n662), .A2(new_n820), .A3(KEYINPUT54), .A4(new_n816), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n818), .A2(KEYINPUT55), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n664), .A2(new_n669), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n817), .A2(KEYINPUT110), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n825), .A2(new_n669), .A3(new_n819), .A4(new_n821), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n826), .A2(KEYINPUT111), .A3(new_n827), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n824), .A2(new_n830), .A3(new_n642), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n617), .A2(new_n621), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n618), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n613), .B1(new_n611), .B2(new_n606), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n624), .A2(new_n634), .B1(new_n629), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n670), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT113), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n832), .A2(new_n841), .A3(new_n838), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n693), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n830), .A2(new_n837), .A3(new_n831), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n824), .A2(new_n258), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT112), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n831), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT111), .B1(new_n826), .B2(new_n827), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n258), .A2(new_n823), .A3(new_n822), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n837), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n846), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n843), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n293), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n749), .A2(new_n670), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n292), .B1(new_n843), .B2(new_n853), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT114), .B1(new_n860), .B2(new_n857), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(new_n697), .A3(new_n678), .A4(new_n595), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n643), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g664(.A1(new_n863), .A2(new_n748), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g666(.A1(new_n863), .A2(new_n293), .ZN(new_n868));
  XOR2_X1   g667(.A(KEYINPUT115), .B(G127gat), .Z(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(G1342gat));
  NOR2_X1   g669(.A1(new_n586), .A2(new_n693), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n862), .A2(new_n697), .A3(new_n871), .ZN(new_n872));
  AND2_X1   g671(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n872), .A2(new_n707), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n874), .B(new_n875), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n642), .A2(new_n419), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT118), .Z(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n859), .A2(new_n861), .A3(new_n697), .A4(new_n721), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n880), .B1(new_n882), .B2(new_n550), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n881), .A2(KEYINPUT119), .A3(new_n689), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n678), .B(new_n879), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n859), .A2(new_n861), .A3(new_n886), .A4(new_n550), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n824), .A2(new_n642), .A3(new_n828), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n838), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n693), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n853), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(KEYINPUT116), .A3(new_n293), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n846), .A2(new_n852), .B1(new_n889), .B2(new_n693), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n292), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n892), .A2(new_n895), .A3(new_n858), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT57), .B1(new_n896), .B2(new_n689), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n684), .A2(new_n485), .A3(new_n586), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n887), .A2(new_n897), .A3(new_n642), .A4(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT58), .B1(new_n899), .B2(G141gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n899), .A2(KEYINPUT117), .A3(G141gat), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT117), .B1(new_n899), .B2(G141gat), .ZN(new_n903));
  NOR4_X1   g702(.A1(new_n881), .A2(new_n689), .A3(new_n586), .A4(new_n878), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(G1344gat));
  NOR2_X1   g706(.A1(new_n748), .A2(G148gat), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n678), .B(new_n908), .C1(new_n883), .C2(new_n884), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n887), .A2(new_n897), .A3(new_n898), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n748), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(KEYINPUT59), .A3(new_n416), .ZN(new_n912));
  XNOR2_X1  g711(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n859), .A2(new_n861), .A3(new_n550), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT57), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n849), .A2(new_n850), .A3(new_n837), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n292), .B1(new_n890), .B2(new_n916), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n886), .B(new_n550), .C1(new_n857), .C2(new_n917), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n915), .A2(new_n670), .A3(new_n898), .A4(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n913), .B1(new_n919), .B2(G148gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n909), .B1(new_n912), .B2(new_n920), .ZN(G1345gat));
  NOR3_X1   g720(.A1(new_n910), .A2(new_n423), .A3(new_n293), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n678), .B(new_n292), .C1(new_n883), .C2(new_n884), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n423), .ZN(G1346gat));
  OAI211_X1 g723(.A(new_n424), .B(new_n871), .C1(new_n883), .C2(new_n884), .ZN(new_n925));
  OAI21_X1  g724(.A(G162gat), .B1(new_n910), .B2(new_n693), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n678), .A2(new_n697), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n859), .A2(new_n861), .A3(new_n595), .A4(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n643), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(G169gat), .Z(G1348gat));
  NOR2_X1   g730(.A1(new_n929), .A2(new_n748), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(G176gat), .Z(G1349gat));
  NOR2_X1   g732(.A1(new_n929), .A2(new_n293), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n307), .A2(new_n311), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(G183gat), .B1(new_n929), .B2(new_n293), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT121), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n940), .A2(KEYINPUT122), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT121), .B1(new_n934), .B2(new_n935), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n939), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n936), .B2(new_n937), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n941), .B1(new_n947), .B2(new_n943), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(new_n948), .ZN(G1350gat));
  XNOR2_X1  g748(.A(KEYINPUT61), .B(G190gat), .ZN(new_n950));
  NAND2_X1  g749(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n929), .A2(new_n693), .ZN(new_n952));
  MUX2_X1   g751(.A(new_n950), .B(new_n951), .S(new_n952), .Z(G1351gat));
  XNOR2_X1  g752(.A(KEYINPUT123), .B(G197gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n684), .A2(new_n697), .A3(new_n678), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n915), .A2(new_n918), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n954), .B1(new_n956), .B2(new_n643), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n859), .A2(new_n550), .A3(new_n861), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(new_n955), .ZN(new_n959));
  INV_X1    g758(.A(new_n954), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n642), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n957), .A2(new_n961), .ZN(G1352gat));
  NAND4_X1  g761(.A1(new_n958), .A2(new_n668), .A3(new_n670), .A4(new_n955), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT124), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n964), .A2(KEYINPUT124), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n915), .A2(new_n670), .A3(new_n918), .A4(new_n955), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n969), .A2(KEYINPUT125), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(KEYINPUT125), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n970), .A2(G204gat), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n968), .A2(new_n972), .ZN(G1353gat));
  NAND4_X1  g772(.A1(new_n915), .A2(new_n292), .A3(new_n918), .A4(new_n955), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G211gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT63), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n975), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n959), .A2(new_n488), .A3(new_n292), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n974), .A2(new_n977), .A3(new_n978), .A4(G211gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(G1354gat));
  NOR3_X1   g782(.A1(new_n956), .A2(new_n489), .A3(new_n693), .ZN(new_n984));
  AOI21_X1  g783(.A(G218gat), .B1(new_n959), .B2(new_n258), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n984), .A2(new_n985), .ZN(G1355gat));
endmodule


