

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U555 ( .A(n688), .B(n687), .ZN(n719) );
  XOR2_X1 U556 ( .A(KEYINPUT66), .B(n555), .Z(n896) );
  AND2_X1 U557 ( .A1(n764), .A2(n763), .ZN(n766) );
  XNOR2_X1 U558 ( .A(n744), .B(KEYINPUT90), .ZN(n747) );
  OR2_X1 U559 ( .A1(n686), .A2(n685), .ZN(n688) );
  INV_X1 U560 ( .A(KEYINPUT67), .ZN(n548) );
  XNOR2_X1 U561 ( .A(KEYINPUT28), .B(n746), .ZN(n518) );
  INV_X1 U562 ( .A(n767), .ZN(n722) );
  NOR2_X1 U563 ( .A1(n952), .A2(n733), .ZN(n734) );
  NOR2_X1 U564 ( .A1(n745), .A2(G299), .ZN(n727) );
  AND2_X1 U565 ( .A1(n747), .A2(n518), .ZN(n748) );
  INV_X1 U566 ( .A(KEYINPUT93), .ZN(n765) );
  XNOR2_X1 U567 ( .A(n766), .B(n765), .ZN(n773) );
  NAND2_X1 U568 ( .A1(n787), .A2(n786), .ZN(n809) );
  NAND2_X2 U569 ( .A1(n719), .A2(n718), .ZN(n767) );
  NOR2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n547) );
  INV_X1 U571 ( .A(G2105), .ZN(n554) );
  NOR2_X1 U572 ( .A1(G543), .A2(G651), .ZN(n632) );
  XNOR2_X1 U573 ( .A(n549), .B(n548), .ZN(n553) );
  NAND2_X1 U574 ( .A1(G91), .A2(n632), .ZN(n522) );
  XNOR2_X1 U575 ( .A(KEYINPUT1), .B(KEYINPUT71), .ZN(n520) );
  XOR2_X1 U576 ( .A(G651), .B(KEYINPUT68), .Z(n523) );
  NOR2_X1 U577 ( .A1(G543), .A2(n523), .ZN(n519) );
  XNOR2_X1 U578 ( .A(n520), .B(n519), .ZN(n646) );
  NAND2_X1 U579 ( .A1(G65), .A2(n646), .ZN(n521) );
  NAND2_X1 U580 ( .A1(n522), .A2(n521), .ZN(n529) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n641) );
  OR2_X1 U582 ( .A1(n641), .A2(n523), .ZN(n524) );
  XNOR2_X1 U583 ( .A(KEYINPUT69), .B(n524), .ZN(n635) );
  NAND2_X1 U584 ( .A1(n635), .A2(G78), .ZN(n527) );
  NOR2_X1 U585 ( .A1(n641), .A2(G651), .ZN(n525) );
  XNOR2_X1 U586 ( .A(KEYINPUT64), .B(n525), .ZN(n642) );
  NAND2_X1 U587 ( .A1(G53), .A2(n642), .ZN(n526) );
  NAND2_X1 U588 ( .A1(n527), .A2(n526), .ZN(n528) );
  OR2_X1 U589 ( .A1(n529), .A2(n528), .ZN(G299) );
  XOR2_X1 U590 ( .A(KEYINPUT99), .B(G2435), .Z(n531) );
  XNOR2_X1 U591 ( .A(G2430), .B(G2438), .ZN(n530) );
  XNOR2_X1 U592 ( .A(n531), .B(n530), .ZN(n538) );
  XOR2_X1 U593 ( .A(G2446), .B(G2454), .Z(n533) );
  XNOR2_X1 U594 ( .A(G2451), .B(G2443), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U596 ( .A(n534), .B(G2427), .Z(n536) );
  XNOR2_X1 U597 ( .A(G1348), .B(G1341), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U599 ( .A(n538), .B(n537), .ZN(n539) );
  AND2_X1 U600 ( .A1(n539), .A2(G14), .ZN(G401) );
  NAND2_X1 U601 ( .A1(n646), .A2(G64), .ZN(n541) );
  NAND2_X1 U602 ( .A1(G52), .A2(n642), .ZN(n540) );
  NAND2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n546) );
  NAND2_X1 U604 ( .A1(G90), .A2(n632), .ZN(n543) );
  NAND2_X1 U605 ( .A1(G77), .A2(n635), .ZN(n542) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(n544), .Z(n545) );
  NOR2_X1 U608 ( .A1(n546), .A2(n545), .ZN(G171) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U610 ( .A(G69), .ZN(G235) );
  INV_X1 U611 ( .A(G132), .ZN(G219) );
  INV_X1 U612 ( .A(G82), .ZN(G220) );
  XOR2_X2 U613 ( .A(KEYINPUT17), .B(n547), .Z(n903) );
  NAND2_X1 U614 ( .A1(n903), .A2(G137), .ZN(n549) );
  AND2_X1 U615 ( .A1(n554), .A2(G2104), .ZN(n901) );
  NAND2_X1 U616 ( .A1(G101), .A2(n901), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(KEYINPUT65), .ZN(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT23), .B(n551), .ZN(n552) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n686) );
  NOR2_X1 U620 ( .A1(G2104), .A2(n554), .ZN(n898) );
  NAND2_X1 U621 ( .A1(n898), .A2(G125), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G2105), .A2(G2104), .ZN(n555) );
  NAND2_X1 U623 ( .A1(G113), .A2(n896), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n683) );
  NOR2_X1 U625 ( .A1(n686), .A2(n683), .ZN(G160) );
  NAND2_X1 U626 ( .A1(G89), .A2(n632), .ZN(n558) );
  XOR2_X1 U627 ( .A(KEYINPUT75), .B(n558), .Z(n559) );
  XNOR2_X1 U628 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G76), .A2(n635), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n562), .B(KEYINPUT5), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n646), .A2(G63), .ZN(n564) );
  NAND2_X1 U633 ( .A1(G51), .A2(n642), .ZN(n563) );
  NAND2_X1 U634 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U635 ( .A(KEYINPUT6), .B(n565), .Z(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n568), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U640 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U641 ( .A(G223), .ZN(n841) );
  NAND2_X1 U642 ( .A1(n841), .A2(G567), .ZN(n570) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n572) );
  NAND2_X1 U645 ( .A1(G56), .A2(n646), .ZN(n571) );
  XNOR2_X1 U646 ( .A(n572), .B(n571), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n632), .A2(G81), .ZN(n573) );
  XNOR2_X1 U648 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U649 ( .A1(G68), .A2(n635), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U651 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U653 ( .A1(G43), .A2(n642), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n580), .A2(n579), .ZN(n952) );
  INV_X1 U655 ( .A(G860), .ZN(n595) );
  OR2_X1 U656 ( .A1(n952), .A2(n595), .ZN(G153) );
  INV_X1 U657 ( .A(G171), .ZN(G301) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n642), .A2(G54), .ZN(n581) );
  XNOR2_X1 U660 ( .A(n581), .B(KEYINPUT74), .ZN(n588) );
  NAND2_X1 U661 ( .A1(G66), .A2(n646), .ZN(n583) );
  NAND2_X1 U662 ( .A1(G79), .A2(n635), .ZN(n582) );
  NAND2_X1 U663 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U664 ( .A1(G92), .A2(n632), .ZN(n584) );
  XNOR2_X1 U665 ( .A(KEYINPUT73), .B(n584), .ZN(n585) );
  NOR2_X1 U666 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U668 ( .A(KEYINPUT15), .B(n589), .ZN(n965) );
  OR2_X1 U669 ( .A1(n965), .A2(G868), .ZN(n590) );
  NAND2_X1 U670 ( .A1(n591), .A2(n590), .ZN(G284) );
  INV_X1 U671 ( .A(G868), .ZN(n659) );
  XNOR2_X1 U672 ( .A(KEYINPUT76), .B(n659), .ZN(n592) );
  NOR2_X1 U673 ( .A1(G286), .A2(n592), .ZN(n594) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U675 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n595), .A2(G559), .ZN(n596) );
  NAND2_X1 U677 ( .A1(n596), .A2(n965), .ZN(n597) );
  XNOR2_X1 U678 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U679 ( .A1(G868), .A2(n952), .ZN(n600) );
  NAND2_X1 U680 ( .A1(G868), .A2(n965), .ZN(n598) );
  NOR2_X1 U681 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U682 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G99), .A2(n901), .ZN(n602) );
  NAND2_X1 U684 ( .A1(G111), .A2(n896), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n602), .A2(n601), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n898), .A2(G123), .ZN(n603) );
  XNOR2_X1 U687 ( .A(n603), .B(KEYINPUT18), .ZN(n605) );
  NAND2_X1 U688 ( .A1(G135), .A2(n903), .ZN(n604) );
  NAND2_X1 U689 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U690 ( .A(KEYINPUT77), .B(n606), .Z(n607) );
  NOR2_X1 U691 ( .A1(n608), .A2(n607), .ZN(n992) );
  XNOR2_X1 U692 ( .A(n992), .B(G2096), .ZN(n610) );
  INV_X1 U693 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U694 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U695 ( .A1(n965), .A2(G559), .ZN(n656) );
  XNOR2_X1 U696 ( .A(n952), .B(n656), .ZN(n611) );
  NOR2_X1 U697 ( .A1(n611), .A2(G860), .ZN(n618) );
  NAND2_X1 U698 ( .A1(G93), .A2(n632), .ZN(n613) );
  NAND2_X1 U699 ( .A1(G67), .A2(n646), .ZN(n612) );
  NAND2_X1 U700 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n635), .A2(G80), .ZN(n615) );
  NAND2_X1 U702 ( .A1(G55), .A2(n642), .ZN(n614) );
  NAND2_X1 U703 ( .A1(n615), .A2(n614), .ZN(n616) );
  OR2_X1 U704 ( .A1(n617), .A2(n616), .ZN(n658) );
  XOR2_X1 U705 ( .A(n618), .B(n658), .Z(G145) );
  NAND2_X1 U706 ( .A1(G88), .A2(n632), .ZN(n620) );
  NAND2_X1 U707 ( .A1(G75), .A2(n635), .ZN(n619) );
  NAND2_X1 U708 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n646), .A2(G62), .ZN(n622) );
  NAND2_X1 U710 ( .A1(G50), .A2(n642), .ZN(n621) );
  NAND2_X1 U711 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U712 ( .A1(n624), .A2(n623), .ZN(G166) );
  NAND2_X1 U713 ( .A1(G86), .A2(n632), .ZN(n626) );
  NAND2_X1 U714 ( .A1(G48), .A2(n642), .ZN(n625) );
  NAND2_X1 U715 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U716 ( .A1(n635), .A2(G73), .ZN(n627) );
  XOR2_X1 U717 ( .A(KEYINPUT2), .B(n627), .Z(n628) );
  NOR2_X1 U718 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U719 ( .A1(n646), .A2(G61), .ZN(n630) );
  NAND2_X1 U720 ( .A1(n631), .A2(n630), .ZN(G305) );
  NAND2_X1 U721 ( .A1(G85), .A2(n632), .ZN(n634) );
  NAND2_X1 U722 ( .A1(G47), .A2(n642), .ZN(n633) );
  NAND2_X1 U723 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U724 ( .A1(G72), .A2(n635), .ZN(n636) );
  XOR2_X1 U725 ( .A(KEYINPUT70), .B(n636), .Z(n637) );
  NOR2_X1 U726 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n646), .A2(G60), .ZN(n639) );
  NAND2_X1 U728 ( .A1(n640), .A2(n639), .ZN(G290) );
  NAND2_X1 U729 ( .A1(n641), .A2(G87), .ZN(n644) );
  NAND2_X1 U730 ( .A1(G49), .A2(n642), .ZN(n643) );
  NAND2_X1 U731 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U732 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U733 ( .A1(G651), .A2(G74), .ZN(n647) );
  NAND2_X1 U734 ( .A1(n648), .A2(n647), .ZN(G288) );
  XNOR2_X1 U735 ( .A(G166), .B(G299), .ZN(n655) );
  XOR2_X1 U736 ( .A(n658), .B(KEYINPUT78), .Z(n649) );
  XNOR2_X1 U737 ( .A(n649), .B(KEYINPUT19), .ZN(n652) );
  XOR2_X1 U738 ( .A(G290), .B(n952), .Z(n650) );
  XNOR2_X1 U739 ( .A(G305), .B(n650), .ZN(n651) );
  XNOR2_X1 U740 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U741 ( .A(n653), .B(G288), .ZN(n654) );
  XNOR2_X1 U742 ( .A(n655), .B(n654), .ZN(n849) );
  XNOR2_X1 U743 ( .A(n656), .B(n849), .ZN(n657) );
  NAND2_X1 U744 ( .A1(n657), .A2(G868), .ZN(n661) );
  NAND2_X1 U745 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U746 ( .A1(n661), .A2(n660), .ZN(G295) );
  XNOR2_X1 U747 ( .A(KEYINPUT20), .B(KEYINPUT80), .ZN(n664) );
  NAND2_X1 U748 ( .A1(G2084), .A2(G2078), .ZN(n662) );
  XNOR2_X1 U749 ( .A(n662), .B(KEYINPUT79), .ZN(n663) );
  XNOR2_X1 U750 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U753 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n668) );
  XNOR2_X1 U756 ( .A(KEYINPUT22), .B(n668), .ZN(n669) );
  NAND2_X1 U757 ( .A1(n669), .A2(G96), .ZN(n670) );
  NOR2_X1 U758 ( .A1(n670), .A2(G218), .ZN(n671) );
  XNOR2_X1 U759 ( .A(n671), .B(KEYINPUT81), .ZN(n847) );
  NAND2_X1 U760 ( .A1(n847), .A2(G2106), .ZN(n675) );
  NAND2_X1 U761 ( .A1(G120), .A2(G108), .ZN(n672) );
  NOR2_X1 U762 ( .A1(G235), .A2(n672), .ZN(n673) );
  NAND2_X1 U763 ( .A1(G57), .A2(n673), .ZN(n848) );
  NAND2_X1 U764 ( .A1(n848), .A2(G567), .ZN(n674) );
  NAND2_X1 U765 ( .A1(n675), .A2(n674), .ZN(n927) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U767 ( .A1(n927), .A2(n676), .ZN(n846) );
  NAND2_X1 U768 ( .A1(n846), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(G138), .A2(n903), .ZN(n678) );
  NAND2_X1 U770 ( .A1(G102), .A2(n901), .ZN(n677) );
  NAND2_X1 U771 ( .A1(n678), .A2(n677), .ZN(n682) );
  NAND2_X1 U772 ( .A1(n898), .A2(G126), .ZN(n680) );
  NAND2_X1 U773 ( .A1(G114), .A2(n896), .ZN(n679) );
  NAND2_X1 U774 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U775 ( .A1(n682), .A2(n681), .ZN(G164) );
  INV_X1 U776 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U777 ( .A(G1986), .B(G290), .ZN(n954) );
  INV_X1 U778 ( .A(n683), .ZN(n684) );
  NAND2_X1 U779 ( .A1(G40), .A2(n684), .ZN(n685) );
  INV_X1 U780 ( .A(KEYINPUT82), .ZN(n687) );
  INV_X1 U781 ( .A(n719), .ZN(n689) );
  NOR2_X1 U782 ( .A1(G164), .A2(G1384), .ZN(n718) );
  NOR2_X1 U783 ( .A1(n689), .A2(n718), .ZN(n836) );
  NAND2_X1 U784 ( .A1(n954), .A2(n836), .ZN(n824) );
  XNOR2_X1 U785 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NAND2_X1 U786 ( .A1(G140), .A2(n903), .ZN(n691) );
  NAND2_X1 U787 ( .A1(G104), .A2(n901), .ZN(n690) );
  NAND2_X1 U788 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U789 ( .A(KEYINPUT34), .B(n692), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n898), .A2(G128), .ZN(n694) );
  NAND2_X1 U791 ( .A1(G116), .A2(n896), .ZN(n693) );
  NAND2_X1 U792 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U793 ( .A(KEYINPUT83), .B(n695), .ZN(n696) );
  XNOR2_X1 U794 ( .A(KEYINPUT35), .B(n696), .ZN(n697) );
  NOR2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U796 ( .A(KEYINPUT36), .B(n699), .ZN(n916) );
  NOR2_X1 U797 ( .A1(n825), .A2(n916), .ZN(n989) );
  NAND2_X1 U798 ( .A1(n836), .A2(n989), .ZN(n833) );
  XNOR2_X1 U799 ( .A(n836), .B(KEYINPUT84), .ZN(n715) );
  NAND2_X1 U800 ( .A1(n898), .A2(G129), .ZN(n701) );
  NAND2_X1 U801 ( .A1(G117), .A2(n896), .ZN(n700) );
  NAND2_X1 U802 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U803 ( .A1(n901), .A2(G105), .ZN(n702) );
  XOR2_X1 U804 ( .A(KEYINPUT38), .B(n702), .Z(n703) );
  NOR2_X1 U805 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U806 ( .A1(n903), .A2(G141), .ZN(n705) );
  NAND2_X1 U807 ( .A1(n706), .A2(n705), .ZN(n882) );
  NAND2_X1 U808 ( .A1(G1996), .A2(n882), .ZN(n714) );
  NAND2_X1 U809 ( .A1(G95), .A2(n901), .ZN(n708) );
  NAND2_X1 U810 ( .A1(G107), .A2(n896), .ZN(n707) );
  NAND2_X1 U811 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U812 ( .A1(G131), .A2(n903), .ZN(n710) );
  NAND2_X1 U813 ( .A1(G119), .A2(n898), .ZN(n709) );
  NAND2_X1 U814 ( .A1(n710), .A2(n709), .ZN(n711) );
  OR2_X1 U815 ( .A1(n712), .A2(n711), .ZN(n883) );
  NAND2_X1 U816 ( .A1(G1991), .A2(n883), .ZN(n713) );
  NAND2_X1 U817 ( .A1(n714), .A2(n713), .ZN(n985) );
  NAND2_X1 U818 ( .A1(n715), .A2(n985), .ZN(n716) );
  XNOR2_X1 U819 ( .A(n716), .B(KEYINPUT85), .ZN(n829) );
  INV_X1 U820 ( .A(n829), .ZN(n717) );
  NAND2_X1 U821 ( .A1(n833), .A2(n717), .ZN(n822) );
  NAND2_X1 U822 ( .A1(G8), .A2(n767), .ZN(n793) );
  NOR2_X1 U823 ( .A1(G1981), .A2(G305), .ZN(n720) );
  XOR2_X1 U824 ( .A(n720), .B(KEYINPUT24), .Z(n721) );
  NOR2_X1 U825 ( .A1(n793), .A2(n721), .ZN(n820) );
  NAND2_X1 U826 ( .A1(n722), .A2(G2072), .ZN(n724) );
  INV_X1 U827 ( .A(KEYINPUT27), .ZN(n723) );
  XNOR2_X1 U828 ( .A(n724), .B(n723), .ZN(n726) );
  NAND2_X1 U829 ( .A1(G1956), .A2(n767), .ZN(n725) );
  NAND2_X1 U830 ( .A1(n726), .A2(n725), .ZN(n745) );
  XNOR2_X1 U831 ( .A(n727), .B(KEYINPUT89), .ZN(n743) );
  INV_X1 U832 ( .A(G1996), .ZN(n728) );
  NOR2_X1 U833 ( .A1(n767), .A2(n728), .ZN(n730) );
  INV_X1 U834 ( .A(KEYINPUT26), .ZN(n729) );
  XNOR2_X1 U835 ( .A(n730), .B(n729), .ZN(n732) );
  NAND2_X1 U836 ( .A1(n767), .A2(G1341), .ZN(n731) );
  NAND2_X1 U837 ( .A1(n732), .A2(n731), .ZN(n733) );
  OR2_X1 U838 ( .A1(n734), .A2(n965), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n965), .A2(n734), .ZN(n739) );
  INV_X1 U840 ( .A(G2067), .ZN(n932) );
  NOR2_X1 U841 ( .A1(n767), .A2(n932), .ZN(n735) );
  XOR2_X1 U842 ( .A(n735), .B(KEYINPUT88), .Z(n737) );
  NAND2_X1 U843 ( .A1(n767), .A2(G1348), .ZN(n736) );
  NAND2_X1 U844 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U845 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U846 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U847 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U848 ( .A1(G299), .A2(n745), .ZN(n746) );
  XNOR2_X1 U849 ( .A(n748), .B(KEYINPUT29), .ZN(n778) );
  XOR2_X1 U850 ( .A(G2078), .B(KEYINPUT86), .Z(n749) );
  XNOR2_X1 U851 ( .A(KEYINPUT25), .B(n749), .ZN(n938) );
  NOR2_X1 U852 ( .A1(n767), .A2(n938), .ZN(n750) );
  XNOR2_X1 U853 ( .A(n750), .B(KEYINPUT87), .ZN(n752) );
  INV_X1 U854 ( .A(G1961), .ZN(n1015) );
  NAND2_X1 U855 ( .A1(n1015), .A2(n767), .ZN(n751) );
  NAND2_X1 U856 ( .A1(n752), .A2(n751), .ZN(n757) );
  NAND2_X1 U857 ( .A1(G171), .A2(n757), .ZN(n777) );
  AND2_X1 U858 ( .A1(n777), .A2(G286), .ZN(n753) );
  NAND2_X1 U859 ( .A1(n778), .A2(n753), .ZN(n764) );
  INV_X1 U860 ( .A(G286), .ZN(n762) );
  NOR2_X1 U861 ( .A1(G1966), .A2(n793), .ZN(n783) );
  NOR2_X1 U862 ( .A1(G2084), .A2(n767), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n783), .A2(n776), .ZN(n754) );
  NAND2_X1 U864 ( .A1(G8), .A2(n754), .ZN(n755) );
  XNOR2_X1 U865 ( .A(KEYINPUT30), .B(n755), .ZN(n756) );
  NOR2_X1 U866 ( .A1(G168), .A2(n756), .ZN(n759) );
  NOR2_X1 U867 ( .A1(G171), .A2(n757), .ZN(n758) );
  NOR2_X1 U868 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U869 ( .A(KEYINPUT31), .B(n760), .ZN(n761) );
  XNOR2_X1 U870 ( .A(n761), .B(KEYINPUT91), .ZN(n780) );
  OR2_X1 U871 ( .A1(n762), .A2(n780), .ZN(n763) );
  NOR2_X1 U872 ( .A1(G1971), .A2(n793), .ZN(n769) );
  NOR2_X1 U873 ( .A1(G2090), .A2(n767), .ZN(n768) );
  NOR2_X1 U874 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U875 ( .A1(n770), .A2(G303), .ZN(n771) );
  XNOR2_X1 U876 ( .A(KEYINPUT94), .B(n771), .ZN(n772) );
  NAND2_X1 U877 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U878 ( .A1(G8), .A2(n774), .ZN(n775) );
  XNOR2_X1 U879 ( .A(n775), .B(KEYINPUT32), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G8), .A2(n776), .ZN(n785) );
  NAND2_X1 U881 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U882 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U883 ( .A(n781), .B(KEYINPUT92), .Z(n782) );
  NOR2_X1 U884 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U885 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U886 ( .A1(G2090), .A2(G303), .ZN(n788) );
  NAND2_X1 U887 ( .A1(G8), .A2(n788), .ZN(n789) );
  NAND2_X1 U888 ( .A1(n809), .A2(n789), .ZN(n790) );
  NAND2_X1 U889 ( .A1(n790), .A2(n793), .ZN(n818) );
  NOR2_X1 U890 ( .A1(G1971), .A2(G303), .ZN(n791) );
  XOR2_X1 U891 ( .A(n791), .B(KEYINPUT95), .Z(n792) );
  NOR2_X1 U892 ( .A1(KEYINPUT33), .A2(n792), .ZN(n807) );
  XOR2_X1 U893 ( .A(G1981), .B(G305), .Z(n966) );
  INV_X1 U894 ( .A(n966), .ZN(n806) );
  INV_X1 U895 ( .A(n793), .ZN(n795) );
  NAND2_X1 U896 ( .A1(n795), .A2(KEYINPUT33), .ZN(n799) );
  NOR2_X1 U897 ( .A1(G1976), .A2(G288), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n803), .A2(KEYINPUT96), .ZN(n794) );
  OR2_X1 U899 ( .A1(n799), .A2(n794), .ZN(n802) );
  INV_X1 U900 ( .A(KEYINPUT33), .ZN(n797) );
  NAND2_X1 U901 ( .A1(G1976), .A2(G288), .ZN(n955) );
  NAND2_X1 U902 ( .A1(n795), .A2(n955), .ZN(n796) );
  NAND2_X1 U903 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U904 ( .A1(n798), .A2(KEYINPUT96), .ZN(n800) );
  NAND2_X1 U905 ( .A1(n800), .A2(n799), .ZN(n801) );
  AND2_X1 U906 ( .A1(n802), .A2(n801), .ZN(n811) );
  INV_X1 U907 ( .A(n811), .ZN(n804) );
  INV_X1 U908 ( .A(n803), .ZN(n956) );
  OR2_X1 U909 ( .A1(n804), .A2(n956), .ZN(n805) );
  OR2_X1 U910 ( .A1(n806), .A2(n805), .ZN(n810) );
  AND2_X1 U911 ( .A1(n807), .A2(n810), .ZN(n808) );
  NAND2_X1 U912 ( .A1(n809), .A2(n808), .ZN(n816) );
  INV_X1 U913 ( .A(n810), .ZN(n814) );
  AND2_X1 U914 ( .A1(KEYINPUT96), .A2(n811), .ZN(n812) );
  AND2_X1 U915 ( .A1(n812), .A2(n966), .ZN(n813) );
  OR2_X1 U916 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U917 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U918 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U919 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n839) );
  NAND2_X1 U922 ( .A1(n825), .A2(n916), .ZN(n986) );
  NOR2_X1 U923 ( .A1(G1996), .A2(n882), .ZN(n826) );
  XOR2_X1 U924 ( .A(KEYINPUT97), .B(n826), .Z(n983) );
  NOR2_X1 U925 ( .A1(G1991), .A2(n883), .ZN(n988) );
  NOR2_X1 U926 ( .A1(G1986), .A2(G290), .ZN(n827) );
  NOR2_X1 U927 ( .A1(n988), .A2(n827), .ZN(n828) );
  NOR2_X1 U928 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U929 ( .A1(n983), .A2(n830), .ZN(n831) );
  XNOR2_X1 U930 ( .A(KEYINPUT39), .B(n831), .ZN(n832) );
  XNOR2_X1 U931 ( .A(n832), .B(KEYINPUT98), .ZN(n834) );
  NAND2_X1 U932 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U933 ( .A1(n986), .A2(n835), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U936 ( .A(KEYINPUT40), .B(n840), .ZN(G329) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n841), .ZN(G217) );
  INV_X1 U938 ( .A(G661), .ZN(n843) );
  NAND2_X1 U939 ( .A1(G2), .A2(G15), .ZN(n842) );
  NOR2_X1 U940 ( .A1(n843), .A2(n842), .ZN(n844) );
  XOR2_X1 U941 ( .A(KEYINPUT100), .B(n844), .Z(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U943 ( .A1(n846), .A2(n845), .ZN(G188) );
  XNOR2_X1 U944 ( .A(G120), .B(KEYINPUT101), .ZN(G236) );
  NOR2_X1 U945 ( .A1(n848), .A2(n847), .ZN(G325) );
  XOR2_X1 U946 ( .A(KEYINPUT102), .B(G325), .Z(G261) );
  XOR2_X1 U947 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  INV_X1 U949 ( .A(G96), .ZN(G221) );
  XOR2_X1 U950 ( .A(n849), .B(G286), .Z(n851) );
  XNOR2_X1 U951 ( .A(G171), .B(n965), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n852) );
  NOR2_X1 U953 ( .A1(G37), .A2(n852), .ZN(G397) );
  XOR2_X1 U954 ( .A(KEYINPUT104), .B(G2678), .Z(n854) );
  XNOR2_X1 U955 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U957 ( .A(KEYINPUT42), .B(G2090), .Z(n856) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U960 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U961 ( .A(G2096), .B(G2100), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n862) );
  XOR2_X1 U963 ( .A(G2084), .B(G2078), .Z(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U965 ( .A(G1976), .B(G1981), .Z(n864) );
  XNOR2_X1 U966 ( .A(G1966), .B(G1956), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U968 ( .A(n865), .B(KEYINPUT41), .Z(n867) );
  XNOR2_X1 U969 ( .A(G1996), .B(G1991), .ZN(n866) );
  XNOR2_X1 U970 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U971 ( .A(G2474), .B(G1971), .Z(n869) );
  XNOR2_X1 U972 ( .A(G1986), .B(G1961), .ZN(n868) );
  XNOR2_X1 U973 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U974 ( .A(n871), .B(n870), .ZN(G229) );
  XOR2_X1 U975 ( .A(KEYINPUT44), .B(KEYINPUT106), .Z(n873) );
  NAND2_X1 U976 ( .A1(G124), .A2(n898), .ZN(n872) );
  XNOR2_X1 U977 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n874), .B(KEYINPUT105), .ZN(n877) );
  NAND2_X1 U979 ( .A1(G100), .A2(n901), .ZN(n875) );
  XOR2_X1 U980 ( .A(KEYINPUT107), .B(n875), .Z(n876) );
  NAND2_X1 U981 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G136), .A2(n903), .ZN(n879) );
  NAND2_X1 U983 ( .A1(G112), .A2(n896), .ZN(n878) );
  NAND2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U985 ( .A1(n881), .A2(n880), .ZN(G162) );
  XNOR2_X1 U986 ( .A(G164), .B(n882), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n888) );
  XOR2_X1 U988 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n886) );
  XNOR2_X1 U989 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U990 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U991 ( .A(n888), .B(n887), .Z(n912) );
  NAND2_X1 U992 ( .A1(G139), .A2(n903), .ZN(n890) );
  NAND2_X1 U993 ( .A1(G103), .A2(n901), .ZN(n889) );
  NAND2_X1 U994 ( .A1(n890), .A2(n889), .ZN(n895) );
  NAND2_X1 U995 ( .A1(n898), .A2(G127), .ZN(n892) );
  NAND2_X1 U996 ( .A1(G115), .A2(n896), .ZN(n891) );
  NAND2_X1 U997 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U998 ( .A(KEYINPUT47), .B(n893), .Z(n894) );
  NOR2_X1 U999 ( .A1(n895), .A2(n894), .ZN(n977) );
  NAND2_X1 U1000 ( .A1(G118), .A2(n896), .ZN(n897) );
  XNOR2_X1 U1001 ( .A(n897), .B(KEYINPUT108), .ZN(n900) );
  NAND2_X1 U1002 ( .A1(G130), .A2(n898), .ZN(n899) );
  NAND2_X1 U1003 ( .A1(n900), .A2(n899), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(n901), .A2(G106), .ZN(n902) );
  XOR2_X1 U1005 ( .A(KEYINPUT109), .B(n902), .Z(n905) );
  NAND2_X1 U1006 ( .A1(n903), .A2(G142), .ZN(n904) );
  NAND2_X1 U1007 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1008 ( .A(KEYINPUT110), .B(n906), .Z(n907) );
  XNOR2_X1 U1009 ( .A(KEYINPUT45), .B(n907), .ZN(n908) );
  NOR2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(n977), .B(n910), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1013 ( .A(n913), .B(G162), .Z(n915) );
  XNOR2_X1 U1014 ( .A(G160), .B(n992), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(n915), .B(n914), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n918), .ZN(G395) );
  NOR2_X1 U1018 ( .A1(G401), .A2(n927), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G227), .A2(G229), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n919) );
  XNOR2_X1 U1021 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1022 ( .A(KEYINPUT49), .B(n921), .Z(n922) );
  NOR2_X1 U1023 ( .A1(G397), .A2(n922), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(n925), .A2(G395), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n926), .B(KEYINPUT115), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(n927), .ZN(G319) );
  INV_X1 U1029 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1030 ( .A(G25), .B(G1991), .ZN(n928) );
  XNOR2_X1 U1031 ( .A(n928), .B(KEYINPUT121), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(G1996), .B(G32), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(G33), .B(G2072), .ZN(n929) );
  NOR2_X1 U1034 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1035 ( .A1(G28), .A2(n931), .ZN(n935) );
  XOR2_X1 U1036 ( .A(KEYINPUT122), .B(n932), .Z(n933) );
  XNOR2_X1 U1037 ( .A(G26), .B(n933), .ZN(n934) );
  NOR2_X1 U1038 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(G27), .B(n938), .ZN(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(n941), .B(KEYINPUT123), .ZN(n942) );
  XNOR2_X1 U1043 ( .A(n942), .B(KEYINPUT53), .ZN(n945) );
  XOR2_X1 U1044 ( .A(G2084), .B(G34), .Z(n943) );
  XNOR2_X1 U1045 ( .A(KEYINPUT54), .B(n943), .ZN(n944) );
  NAND2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(G35), .B(G2090), .ZN(n946) );
  NOR2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1049 ( .A(KEYINPUT55), .B(n948), .ZN(n950) );
  INV_X1 U1050 ( .A(G29), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1052 ( .A1(n951), .A2(G11), .ZN(n976) );
  XOR2_X1 U1053 ( .A(KEYINPUT56), .B(G16), .Z(n974) );
  XNOR2_X1 U1054 ( .A(G1341), .B(n952), .ZN(n953) );
  NOR2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G171), .B(G1961), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(G299), .B(G1956), .ZN(n958) );
  XNOR2_X1 U1059 ( .A(G303), .B(G1971), .ZN(n957) );
  NOR2_X1 U1060 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G1348), .B(n965), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(G1966), .B(G168), .ZN(n967) );
  NAND2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(n968), .B(KEYINPUT57), .ZN(n969) );
  NAND2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n1007) );
  XNOR2_X1 U1072 ( .A(G164), .B(G2078), .ZN(n980) );
  XOR2_X1 U1073 ( .A(G2072), .B(n977), .Z(n978) );
  XNOR2_X1 U1074 ( .A(KEYINPUT119), .B(n978), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(n981), .B(KEYINPUT50), .ZN(n1001) );
  XOR2_X1 U1077 ( .A(G2090), .B(G162), .Z(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1079 ( .A(KEYINPUT51), .B(n984), .Z(n999) );
  INV_X1 U1080 ( .A(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n997) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G2084), .B(G160), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(KEYINPUT117), .B(n990), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(KEYINPUT118), .B(n995), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1091 ( .A(KEYINPUT52), .B(n1002), .Z(n1003) );
  NOR2_X1 U1092 ( .A1(KEYINPUT55), .A2(n1003), .ZN(n1004) );
  XOR2_X1 U1093 ( .A(KEYINPUT120), .B(n1004), .Z(n1005) );
  NAND2_X1 U1094 ( .A1(G29), .A2(n1005), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1035) );
  XOR2_X1 U1096 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n1014) );
  XNOR2_X1 U1097 ( .A(G1986), .B(G24), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G22), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(G1976), .B(KEYINPUT126), .Z(n1010) );
  XNOR2_X1 U1101 ( .A(G23), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(n1014), .B(n1013), .ZN(n1031) );
  XNOR2_X1 U1104 ( .A(G5), .B(n1015), .ZN(n1029) );
  XOR2_X1 U1105 ( .A(G1348), .B(KEYINPUT59), .Z(n1016) );
  XNOR2_X1 U1106 ( .A(G4), .B(n1016), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(G1981), .B(G6), .Z(n1019) );
  XOR2_X1 U1108 ( .A(G20), .B(KEYINPUT124), .Z(n1017) );
  XNOR2_X1 U1109 ( .A(n1017), .B(G1956), .ZN(n1018) );
  NAND2_X1 U1110 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  XNOR2_X1 U1111 ( .A(G19), .B(G1341), .ZN(n1020) );
  NOR2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1113 ( .A(n1022), .B(KEYINPUT125), .ZN(n1023) );
  NOR2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1115 ( .A(KEYINPUT60), .B(n1025), .Z(n1027) );
  XNOR2_X1 U1116 ( .A(G1966), .B(G21), .ZN(n1026) );
  NOR2_X1 U1117 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1119 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1120 ( .A(KEYINPUT61), .B(n1032), .Z(n1033) );
  NOR2_X1 U1121 ( .A1(G16), .A2(n1033), .ZN(n1034) );
  NOR2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1123 ( .A(n1036), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

