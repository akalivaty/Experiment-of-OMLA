

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751;

  INV_X1 U367 ( .A(n560), .ZN(n598) );
  BUF_X1 U368 ( .A(n655), .Z(n389) );
  XOR2_X1 U369 ( .A(G104), .B(G122), .Z(n442) );
  XNOR2_X1 U370 ( .A(G113), .B(G143), .ZN(n441) );
  XNOR2_X1 U371 ( .A(G131), .B(G140), .ZN(n443) );
  BUF_X1 U372 ( .A(G119), .Z(n390) );
  XNOR2_X1 U373 ( .A(G128), .B(KEYINPUT24), .ZN(n485) );
  XNOR2_X1 U374 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n454) );
  NAND2_X2 U375 ( .A1(G214), .A2(n429), .ZN(n668) );
  INV_X2 U376 ( .A(KEYINPUT64), .ZN(n401) );
  XNOR2_X2 U377 ( .A(n430), .B(KEYINPUT19), .ZN(n436) );
  XNOR2_X2 U378 ( .A(n351), .B(KEYINPUT32), .ZN(n748) );
  XNOR2_X2 U379 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n413) );
  XNOR2_X2 U380 ( .A(n427), .B(G902), .ZN(n603) );
  INV_X1 U381 ( .A(G953), .ZN(n550) );
  INV_X1 U382 ( .A(n389), .ZN(n535) );
  XOR2_X1 U383 ( .A(n486), .B(n485), .Z(n346) );
  NAND2_X2 U384 ( .A1(n352), .A2(n394), .ZN(n397) );
  AND2_X2 U385 ( .A1(n393), .A2(n399), .ZN(n352) );
  NOR2_X1 U386 ( .A1(n750), .A2(n751), .ZN(n577) );
  NOR2_X2 U387 ( .A1(G953), .A2(G237), .ZN(n499) );
  AND2_X1 U388 ( .A1(n368), .A2(n372), .ZN(n371) );
  AND2_X1 U389 ( .A1(n740), .A2(KEYINPUT65), .ZN(n369) );
  XNOR2_X1 U390 ( .A(n366), .B(n365), .ZN(n750) );
  BUF_X1 U391 ( .A(n531), .Z(n660) );
  INV_X2 U392 ( .A(n640), .ZN(n642) );
  XNOR2_X1 U393 ( .A(n531), .B(KEYINPUT101), .ZN(n565) );
  NAND2_X1 U394 ( .A1(n616), .A2(G472), .ZN(n364) );
  XNOR2_X1 U395 ( .A(KEYINPUT87), .B(n488), .ZN(n732) );
  INV_X1 U396 ( .A(KEYINPUT2), .ZN(n375) );
  NAND2_X1 U397 ( .A1(G902), .A2(G472), .ZN(n363) );
  INV_X1 U398 ( .A(KEYINPUT15), .ZN(n427) );
  INV_X1 U399 ( .A(G134), .ZN(n464) );
  XOR2_X2 U400 ( .A(G146), .B(G125), .Z(n447) );
  INV_X1 U401 ( .A(KEYINPUT40), .ZN(n365) );
  INV_X1 U402 ( .A(G472), .ZN(n361) );
  NAND2_X1 U403 ( .A1(n354), .A2(n353), .ZN(n568) );
  NAND2_X1 U404 ( .A1(n561), .A2(n350), .ZN(n349) );
  OR2_X2 U405 ( .A1(n362), .A2(n359), .ZN(n531) );
  NAND2_X1 U406 ( .A1(n364), .A2(n363), .ZN(n362) );
  XOR2_X1 U407 ( .A(KEYINPUT62), .B(n617), .Z(n618) );
  INV_X1 U408 ( .A(n651), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U410 ( .A(n440), .B(KEYINPUT21), .ZN(n651) );
  XOR2_X1 U411 ( .A(n622), .B(KEYINPUT59), .Z(n623) );
  AND2_X1 U412 ( .A1(n604), .A2(n403), .ZN(n370) );
  OR2_X1 U413 ( .A1(n604), .A2(n403), .ZN(n372) );
  NAND2_X1 U414 ( .A1(n361), .A2(n480), .ZN(n360) );
  XNOR2_X2 U415 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n484) );
  NAND2_X1 U416 ( .A1(G234), .A2(G237), .ZN(n431) );
  INV_X1 U417 ( .A(KEYINPUT77), .ZN(n367) );
  XNOR2_X1 U418 ( .A(KEYINPUT70), .B(G113), .ZN(n391) );
  XNOR2_X2 U419 ( .A(G104), .B(KEYINPUT76), .ZN(n419) );
  XOR2_X2 U420 ( .A(G107), .B(KEYINPUT88), .Z(n475) );
  XNOR2_X1 U421 ( .A(G137), .B(G116), .ZN(n500) );
  XOR2_X2 U422 ( .A(KEYINPUT96), .B(KEYINPUT94), .Z(n457) );
  XNOR2_X2 U423 ( .A(G116), .B(G107), .ZN(n418) );
  NOR2_X2 U424 ( .A1(n347), .A2(n676), .ZN(n514) );
  OR2_X2 U425 ( .A1(n347), .A2(n349), .ZN(n348) );
  NOR2_X1 U426 ( .A1(n347), .A2(n568), .ZN(n530) );
  OR2_X1 U427 ( .A1(n662), .A2(n347), .ZN(n536) );
  XNOR2_X2 U428 ( .A(n437), .B(KEYINPUT0), .ZN(n347) );
  XNOR2_X2 U429 ( .A(n348), .B(n384), .ZN(n392) );
  NAND2_X1 U430 ( .A1(n392), .A2(n381), .ZN(n351) );
  NAND2_X1 U431 ( .A1(n524), .A2(n748), .ZN(n546) );
  NAND2_X2 U432 ( .A1(n356), .A2(n371), .ZN(n402) );
  NAND2_X1 U433 ( .A1(n358), .A2(n370), .ZN(n357) );
  AND2_X2 U434 ( .A1(n357), .A2(n373), .ZN(n356) );
  INV_X1 U435 ( .A(n355), .ZN(n353) );
  INV_X1 U436 ( .A(n654), .ZN(n354) );
  XNOR2_X2 U437 ( .A(n355), .B(KEYINPUT1), .ZN(n655) );
  XNOR2_X1 U438 ( .A(n355), .B(KEYINPUT107), .ZN(n557) );
  XNOR2_X2 U439 ( .A(n482), .B(n481), .ZN(n355) );
  NAND2_X1 U440 ( .A1(n397), .A2(n740), .ZN(n358) );
  XNOR2_X2 U441 ( .A(n531), .B(n509), .ZN(n584) );
  NOR2_X1 U442 ( .A1(n616), .A2(n360), .ZN(n359) );
  XNOR2_X2 U443 ( .A(n507), .B(n506), .ZN(n616) );
  NAND2_X1 U444 ( .A1(n601), .A2(n642), .ZN(n366) );
  XNOR2_X2 U445 ( .A(n576), .B(KEYINPUT39), .ZN(n601) );
  AND2_X1 U446 ( .A1(n575), .A2(n560), .ZN(n578) );
  XNOR2_X1 U447 ( .A(n574), .B(n367), .ZN(n575) );
  NOR2_X1 U448 ( .A1(n606), .A2(n375), .ZN(n374) );
  NAND2_X1 U449 ( .A1(n397), .A2(n369), .ZN(n368) );
  NAND2_X1 U450 ( .A1(n374), .A2(n740), .ZN(n373) );
  XNOR2_X2 U451 ( .A(n376), .B(n420), .ZN(n720) );
  XNOR2_X2 U452 ( .A(n505), .B(n414), .ZN(n376) );
  XNOR2_X2 U453 ( .A(n377), .B(n391), .ZN(n505) );
  XNOR2_X2 U454 ( .A(n416), .B(n417), .ZN(n377) );
  XNOR2_X1 U455 ( .A(n439), .B(n438), .ZN(n494) );
  NAND2_X1 U456 ( .A1(n548), .A2(n400), .ZN(n399) );
  NAND2_X1 U457 ( .A1(n395), .A2(n398), .ZN(n394) );
  NOR2_X1 U458 ( .A1(n548), .A2(n400), .ZN(n398) );
  INV_X1 U459 ( .A(n547), .ZN(n405) );
  INV_X1 U460 ( .A(KEYINPUT44), .ZN(n409) );
  XNOR2_X1 U461 ( .A(n498), .B(n497), .ZN(n652) );
  INV_X1 U462 ( .A(KEYINPUT4), .ZN(n470) );
  INV_X1 U463 ( .A(G902), .ZN(n480) );
  XNOR2_X1 U464 ( .A(n390), .B(G110), .ZN(n490) );
  AND2_X2 U465 ( .A1(n396), .A2(n380), .ZN(n740) );
  XNOR2_X1 U466 ( .A(n594), .B(n385), .ZN(n396) );
  INV_X1 U467 ( .A(KEYINPUT80), .ZN(n400) );
  OR2_X1 U468 ( .A1(G237), .A2(G902), .ZN(n429) );
  XNOR2_X1 U469 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n421) );
  INV_X1 U470 ( .A(KEYINPUT45), .ZN(n406) );
  NAND2_X1 U471 ( .A1(n705), .A2(n480), .ZN(n482) );
  BUF_X1 U472 ( .A(n652), .Z(n388) );
  XNOR2_X1 U473 ( .A(KEYINPUT93), .B(KEYINPUT5), .ZN(n502) );
  XNOR2_X1 U474 ( .A(KEYINPUT7), .B(KEYINPUT95), .ZN(n456) );
  NAND2_X1 U475 ( .A1(n575), .A2(n378), .ZN(n576) );
  XNOR2_X1 U476 ( .A(n487), .B(n346), .ZN(n492) );
  AND2_X1 U477 ( .A1(n612), .A2(G953), .ZN(n718) );
  NAND2_X1 U478 ( .A1(n516), .A2(n515), .ZN(n518) );
  INV_X1 U479 ( .A(n581), .ZN(n404) );
  XNOR2_X1 U480 ( .A(KEYINPUT38), .B(n598), .ZN(n378) );
  NAND2_X1 U481 ( .A1(G210), .A2(n429), .ZN(n379) );
  AND2_X1 U482 ( .A1(n602), .A2(n650), .ZN(n380) );
  AND2_X1 U483 ( .A1(n521), .A2(n520), .ZN(n381) );
  AND2_X1 U484 ( .A1(n508), .A2(n565), .ZN(n382) );
  AND2_X1 U485 ( .A1(n526), .A2(n525), .ZN(n383) );
  XOR2_X1 U486 ( .A(n469), .B(n468), .Z(n384) );
  XOR2_X1 U487 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n385) );
  XNOR2_X2 U488 ( .A(n402), .B(n401), .ZN(n386) );
  NOR2_X2 U489 ( .A1(n655), .A2(n654), .ZN(n510) );
  BUF_X1 U490 ( .A(n436), .Z(n387) );
  NAND2_X1 U491 ( .A1(n546), .A2(KEYINPUT44), .ZN(n544) );
  NOR2_X1 U492 ( .A1(n573), .A2(n572), .ZN(n574) );
  AND2_X2 U493 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X2 U494 ( .A(n507), .B(n479), .ZN(n705) );
  NAND2_X1 U495 ( .A1(n392), .A2(n383), .ZN(n528) );
  NAND2_X1 U496 ( .A1(n392), .A2(n382), .ZN(n522) );
  NAND2_X1 U497 ( .A1(n605), .A2(n400), .ZN(n393) );
  INV_X1 U498 ( .A(n605), .ZN(n395) );
  XNOR2_X2 U499 ( .A(n402), .B(n401), .ZN(n700) );
  INV_X1 U500 ( .A(KEYINPUT65), .ZN(n403) );
  NAND2_X1 U501 ( .A1(n404), .A2(n387), .ZN(n639) );
  NAND2_X1 U502 ( .A1(n405), .A2(n409), .ZN(n408) );
  XNOR2_X2 U503 ( .A(n407), .B(n406), .ZN(n605) );
  NAND2_X1 U504 ( .A1(n410), .A2(n408), .ZN(n407) );
  XNOR2_X1 U505 ( .A(n545), .B(n411), .ZN(n410) );
  INV_X1 U506 ( .A(KEYINPUT82), .ZN(n411) );
  NOR2_X1 U507 ( .A1(n532), .A2(n660), .ZN(n412) );
  XNOR2_X1 U508 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n414) );
  OR2_X1 U509 ( .A1(n554), .A2(n435), .ZN(n415) );
  AND2_X1 U510 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U511 ( .A(KEYINPUT90), .B(KEYINPUT20), .ZN(n438) );
  INV_X1 U512 ( .A(n569), .ZN(n570) );
  BUF_X1 U513 ( .A(n676), .Z(n685) );
  BUF_X1 U514 ( .A(n616), .Z(n617) );
  XNOR2_X1 U515 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X2 U516 ( .A(KEYINPUT71), .B(G119), .ZN(n416) );
  XNOR2_X2 U517 ( .A(G101), .B(KEYINPUT3), .ZN(n417) );
  XNOR2_X1 U518 ( .A(n418), .B(G122), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n419), .B(G110), .ZN(n473) );
  XNOR2_X1 U520 ( .A(n459), .B(n473), .ZN(n420) );
  XOR2_X1 U521 ( .A(n447), .B(KEYINPUT18), .Z(n425) );
  XNOR2_X2 U522 ( .A(G143), .B(G128), .ZN(n465) );
  NAND2_X1 U523 ( .A1(G224), .A2(n550), .ZN(n422) );
  XNOR2_X1 U524 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U525 ( .A(n465), .B(n423), .ZN(n424) );
  XNOR2_X1 U526 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U527 ( .A(n720), .B(n426), .ZN(n607) );
  NOR2_X1 U528 ( .A1(n607), .A2(n603), .ZN(n428) );
  XNOR2_X1 U529 ( .A(n428), .B(n379), .ZN(n559) );
  NAND2_X1 U530 ( .A1(n559), .A2(n668), .ZN(n430) );
  XNOR2_X1 U531 ( .A(n431), .B(KEYINPUT14), .ZN(n432) );
  NAND2_X1 U532 ( .A1(G952), .A2(n432), .ZN(n684) );
  NOR2_X1 U533 ( .A1(G953), .A2(n684), .ZN(n554) );
  NAND2_X1 U534 ( .A1(n432), .A2(G902), .ZN(n433) );
  XNOR2_X1 U535 ( .A(KEYINPUT86), .B(n433), .ZN(n549) );
  XOR2_X1 U536 ( .A(G898), .B(KEYINPUT84), .Z(n725) );
  NAND2_X1 U537 ( .A1(n725), .A2(G953), .ZN(n434) );
  XOR2_X1 U538 ( .A(KEYINPUT85), .B(n434), .Z(n719) );
  NOR2_X1 U539 ( .A1(n549), .A2(n719), .ZN(n435) );
  NAND2_X1 U540 ( .A1(n436), .A2(n415), .ZN(n437) );
  INV_X1 U541 ( .A(n603), .ZN(n548) );
  NAND2_X1 U542 ( .A1(n548), .A2(G234), .ZN(n439) );
  NAND2_X1 U543 ( .A1(n494), .A2(G221), .ZN(n440) );
  XNOR2_X1 U544 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U545 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n444) );
  XNOR2_X1 U546 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U547 ( .A(n446), .B(n445), .Z(n451) );
  INV_X1 U548 ( .A(n447), .ZN(n448) );
  XNOR2_X1 U549 ( .A(KEYINPUT10), .B(n448), .ZN(n731) );
  AND2_X1 U550 ( .A1(n499), .A2(G214), .ZN(n449) );
  XNOR2_X1 U551 ( .A(n731), .B(n449), .ZN(n450) );
  XNOR2_X1 U552 ( .A(n451), .B(n450), .ZN(n622) );
  NAND2_X1 U553 ( .A1(n622), .A2(n480), .ZN(n453) );
  XOR2_X1 U554 ( .A(KEYINPUT13), .B(G475), .Z(n452) );
  XNOR2_X1 U555 ( .A(n453), .B(n452), .ZN(n537) );
  NAND2_X1 U556 ( .A1(n550), .A2(G234), .ZN(n455) );
  XNOR2_X1 U557 ( .A(n455), .B(n454), .ZN(n483) );
  NAND2_X1 U558 ( .A1(n483), .A2(G217), .ZN(n463) );
  XOR2_X1 U559 ( .A(KEYINPUT9), .B(KEYINPUT97), .Z(n461) );
  XNOR2_X1 U560 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U561 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U562 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U563 ( .A(n463), .B(n462), .ZN(n466) );
  XNOR2_X2 U564 ( .A(n465), .B(n464), .ZN(n472) );
  XNOR2_X1 U565 ( .A(n472), .B(n466), .ZN(n709) );
  NAND2_X1 U566 ( .A1(n709), .A2(n480), .ZN(n467) );
  XNOR2_X1 U567 ( .A(n467), .B(G478), .ZN(n539) );
  NOR2_X1 U568 ( .A1(n537), .A2(n539), .ZN(n561) );
  XOR2_X1 U569 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n469) );
  XNOR2_X1 U570 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n468) );
  XNOR2_X1 U571 ( .A(n470), .B(G131), .ZN(n471) );
  XNOR2_X2 U572 ( .A(n472), .B(n471), .ZN(n735) );
  XNOR2_X2 U573 ( .A(n735), .B(G146), .ZN(n507) );
  XNOR2_X2 U574 ( .A(G137), .B(G140), .ZN(n488) );
  XNOR2_X1 U575 ( .A(n732), .B(n473), .ZN(n478) );
  NAND2_X1 U576 ( .A1(G227), .A2(n550), .ZN(n474) );
  XNOR2_X1 U577 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U578 ( .A(n476), .B(G101), .ZN(n477) );
  XNOR2_X1 U579 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U580 ( .A(KEYINPUT69), .B(G469), .ZN(n481) );
  NAND2_X1 U581 ( .A1(G221), .A2(n483), .ZN(n487) );
  INV_X1 U582 ( .A(n484), .ZN(n486) );
  INV_X1 U583 ( .A(n488), .ZN(n489) );
  XNOR2_X1 U584 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U585 ( .A(n493), .B(n731), .ZN(n714) );
  NOR2_X1 U586 ( .A1(n714), .A2(G902), .ZN(n498) );
  XOR2_X1 U587 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n496) );
  NAND2_X1 U588 ( .A1(G217), .A2(n494), .ZN(n495) );
  XOR2_X1 U589 ( .A(n496), .B(n495), .Z(n497) );
  INV_X1 U590 ( .A(n388), .ZN(n519) );
  NOR2_X1 U591 ( .A1(n535), .A2(n519), .ZN(n508) );
  NAND2_X1 U592 ( .A1(n499), .A2(G210), .ZN(n501) );
  XNOR2_X1 U593 ( .A(n501), .B(n500), .ZN(n503) );
  XNOR2_X1 U594 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U595 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U596 ( .A(n522), .B(G110), .ZN(G12) );
  OR2_X2 U597 ( .A1(n652), .A2(n651), .ZN(n654) );
  XNOR2_X1 U598 ( .A(KEYINPUT99), .B(KEYINPUT6), .ZN(n509) );
  NAND2_X1 U599 ( .A1(n510), .A2(n584), .ZN(n513) );
  XNOR2_X1 U600 ( .A(KEYINPUT102), .B(KEYINPUT33), .ZN(n511) );
  XNOR2_X1 U601 ( .A(n511), .B(KEYINPUT83), .ZN(n512) );
  XNOR2_X1 U602 ( .A(n513), .B(n512), .ZN(n676) );
  XNOR2_X1 U603 ( .A(n514), .B(n413), .ZN(n516) );
  NAND2_X1 U604 ( .A1(n539), .A2(n537), .ZN(n580) );
  INV_X1 U605 ( .A(n580), .ZN(n515) );
  XNOR2_X1 U606 ( .A(KEYINPUT81), .B(KEYINPUT35), .ZN(n517) );
  XNOR2_X2 U607 ( .A(n518), .B(n517), .ZN(n523) );
  XNOR2_X1 U608 ( .A(n523), .B(G122), .ZN(G24) );
  XOR2_X1 U609 ( .A(KEYINPUT78), .B(n584), .Z(n521) );
  NOR2_X1 U610 ( .A1(n389), .A2(n519), .ZN(n520) );
  NOR2_X1 U611 ( .A1(n535), .A2(n388), .ZN(n526) );
  INV_X1 U612 ( .A(n584), .ZN(n525) );
  INV_X1 U613 ( .A(KEYINPUT100), .ZN(n527) );
  XNOR2_X1 U614 ( .A(n528), .B(n527), .ZN(n747) );
  INV_X1 U615 ( .A(KEYINPUT92), .ZN(n529) );
  XNOR2_X1 U616 ( .A(n530), .B(n529), .ZN(n532) );
  INV_X1 U617 ( .A(n660), .ZN(n533) );
  NOR2_X1 U618 ( .A1(n533), .A2(n654), .ZN(n534) );
  NAND2_X1 U619 ( .A1(n535), .A2(n534), .ZN(n662) );
  XNOR2_X1 U620 ( .A(n536), .B(KEYINPUT31), .ZN(n646) );
  NOR2_X1 U621 ( .A1(n412), .A2(n646), .ZN(n541) );
  INV_X1 U622 ( .A(n537), .ZN(n538) );
  OR2_X1 U623 ( .A1(n539), .A2(n538), .ZN(n640) );
  AND2_X1 U624 ( .A1(n539), .A2(n538), .ZN(n645) );
  NOR2_X1 U625 ( .A1(n642), .A2(n645), .ZN(n540) );
  XNOR2_X1 U626 ( .A(KEYINPUT98), .B(n540), .ZN(n672) );
  NOR2_X1 U627 ( .A1(n541), .A2(n672), .ZN(n542) );
  NOR2_X1 U628 ( .A1(n747), .A2(n542), .ZN(n543) );
  NAND2_X1 U629 ( .A1(n544), .A2(n543), .ZN(n545) );
  BUF_X1 U630 ( .A(n546), .Z(n547) );
  OR2_X1 U631 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U632 ( .A1(G900), .A2(n551), .ZN(n552) );
  XOR2_X1 U633 ( .A(KEYINPUT103), .B(n552), .Z(n553) );
  NOR2_X1 U634 ( .A1(n554), .A2(n553), .ZN(n569) );
  NOR2_X1 U635 ( .A1(n651), .A2(n569), .ZN(n555) );
  NAND2_X1 U636 ( .A1(n388), .A2(n555), .ZN(n587) );
  NOR2_X1 U637 ( .A1(n565), .A2(n587), .ZN(n556) );
  XNOR2_X1 U638 ( .A(n556), .B(KEYINPUT28), .ZN(n558) );
  NAND2_X1 U639 ( .A1(n558), .A2(n557), .ZN(n581) );
  BUF_X1 U640 ( .A(n559), .Z(n560) );
  NAND2_X1 U641 ( .A1(n378), .A2(n668), .ZN(n673) );
  INV_X1 U642 ( .A(n561), .ZN(n671) );
  NOR2_X1 U643 ( .A1(n673), .A2(n671), .ZN(n563) );
  XNOR2_X1 U644 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n562) );
  XNOR2_X1 U645 ( .A(n563), .B(n562), .ZN(n686) );
  NOR2_X1 U646 ( .A1(n581), .A2(n686), .ZN(n564) );
  XNOR2_X1 U647 ( .A(n564), .B(KEYINPUT42), .ZN(n751) );
  INV_X1 U648 ( .A(n565), .ZN(n566) );
  NAND2_X1 U649 ( .A1(n566), .A2(n668), .ZN(n567) );
  XNOR2_X1 U650 ( .A(n567), .B(KEYINPUT30), .ZN(n573) );
  INV_X1 U651 ( .A(n568), .ZN(n571) );
  NAND2_X1 U652 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U653 ( .A(n577), .B(KEYINPUT46), .ZN(n593) );
  XOR2_X1 U654 ( .A(KEYINPUT106), .B(n578), .Z(n579) );
  NOR2_X1 U655 ( .A1(n580), .A2(n579), .ZN(n638) );
  NOR2_X1 U656 ( .A1(n672), .A2(n639), .ZN(n582) );
  XOR2_X1 U657 ( .A(KEYINPUT47), .B(n582), .Z(n583) );
  NOR2_X1 U658 ( .A1(n638), .A2(n583), .ZN(n591) );
  AND2_X1 U659 ( .A1(n642), .A2(n668), .ZN(n585) );
  NAND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n586) );
  OR2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n595) );
  NOR2_X1 U662 ( .A1(n598), .A2(n595), .ZN(n588) );
  XOR2_X1 U663 ( .A(KEYINPUT36), .B(n588), .Z(n589) );
  NOR2_X1 U664 ( .A1(n589), .A2(n389), .ZN(n648) );
  INV_X1 U665 ( .A(n648), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U667 ( .A(KEYINPUT104), .B(n595), .Z(n596) );
  NAND2_X1 U668 ( .A1(n596), .A2(n389), .ZN(n597) );
  XNOR2_X1 U669 ( .A(n597), .B(KEYINPUT43), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT105), .ZN(n746) );
  INV_X1 U672 ( .A(n746), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n601), .A2(n645), .ZN(n650) );
  NAND2_X1 U674 ( .A1(n603), .A2(KEYINPUT2), .ZN(n604) );
  BUF_X1 U675 ( .A(n605), .Z(n606) );
  NAND2_X1 U676 ( .A1(n386), .A2(G210), .ZN(n611) );
  BUF_X1 U677 ( .A(n607), .Z(n609) );
  XNOR2_X1 U678 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n611), .B(n610), .ZN(n613) );
  INV_X1 U680 ( .A(G952), .ZN(n612) );
  INV_X1 U681 ( .A(n718), .ZN(n625) );
  NAND2_X1 U682 ( .A1(n613), .A2(n625), .ZN(n615) );
  INV_X1 U683 ( .A(KEYINPUT56), .ZN(n614) );
  XNOR2_X1 U684 ( .A(n615), .B(n614), .ZN(G51) );
  NAND2_X1 U685 ( .A1(n700), .A2(G472), .ZN(n619) );
  XNOR2_X1 U686 ( .A(n619), .B(n618), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n620), .A2(n625), .ZN(n621) );
  XNOR2_X1 U688 ( .A(n621), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U689 ( .A1(n700), .A2(G475), .ZN(n624) );
  XNOR2_X1 U690 ( .A(n624), .B(n623), .ZN(n626) );
  NAND2_X1 U691 ( .A1(n626), .A2(n625), .ZN(n628) );
  INV_X1 U692 ( .A(KEYINPUT60), .ZN(n627) );
  XNOR2_X1 U693 ( .A(n628), .B(n627), .ZN(G60) );
  NAND2_X1 U694 ( .A1(n412), .A2(n642), .ZN(n629) );
  XNOR2_X1 U695 ( .A(n629), .B(G104), .ZN(G6) );
  XOR2_X1 U696 ( .A(KEYINPUT26), .B(KEYINPUT109), .Z(n631) );
  NAND2_X1 U697 ( .A1(n412), .A2(n645), .ZN(n630) );
  XNOR2_X1 U698 ( .A(n631), .B(n630), .ZN(n633) );
  XOR2_X1 U699 ( .A(G107), .B(KEYINPUT27), .Z(n632) );
  XNOR2_X1 U700 ( .A(n633), .B(n632), .ZN(G9) );
  INV_X1 U701 ( .A(n645), .ZN(n634) );
  NOR2_X1 U702 ( .A1(n634), .A2(n639), .ZN(n636) );
  XNOR2_X1 U703 ( .A(KEYINPUT110), .B(KEYINPUT29), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U705 ( .A(G128), .B(n637), .ZN(G30) );
  XOR2_X1 U706 ( .A(G143), .B(n638), .Z(G45) );
  NOR2_X1 U707 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U708 ( .A(G146), .B(n641), .Z(G48) );
  XOR2_X1 U709 ( .A(G113), .B(KEYINPUT111), .Z(n644) );
  NAND2_X1 U710 ( .A1(n646), .A2(n642), .ZN(n643) );
  XNOR2_X1 U711 ( .A(n644), .B(n643), .ZN(G15) );
  NAND2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U713 ( .A(n647), .B(G116), .ZN(G18) );
  XNOR2_X1 U714 ( .A(n648), .B(G125), .ZN(n649) );
  XNOR2_X1 U715 ( .A(n649), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U716 ( .A(G134), .B(n650), .ZN(G36) );
  XNOR2_X1 U717 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n681) );
  AND2_X1 U718 ( .A1(n388), .A2(n651), .ZN(n653) );
  XNOR2_X1 U719 ( .A(KEYINPUT49), .B(n653), .ZN(n659) );
  NAND2_X1 U720 ( .A1(n389), .A2(n654), .ZN(n656) );
  XNOR2_X1 U721 ( .A(n656), .B(KEYINPUT112), .ZN(n657) );
  XNOR2_X1 U722 ( .A(KEYINPUT50), .B(n657), .ZN(n658) );
  NAND2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n661) );
  NOR2_X1 U724 ( .A1(n661), .A2(n660), .ZN(n664) );
  INV_X1 U725 ( .A(n662), .ZN(n663) );
  NOR2_X1 U726 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U727 ( .A(n665), .B(KEYINPUT113), .ZN(n666) );
  XNOR2_X1 U728 ( .A(KEYINPUT51), .B(n666), .ZN(n667) );
  NOR2_X1 U729 ( .A1(n686), .A2(n667), .ZN(n679) );
  NOR2_X1 U730 ( .A1(n378), .A2(n668), .ZN(n669) );
  XNOR2_X1 U731 ( .A(n669), .B(KEYINPUT114), .ZN(n670) );
  NOR2_X1 U732 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U733 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U734 ( .A1(n675), .A2(n674), .ZN(n677) );
  NOR2_X1 U735 ( .A1(n677), .A2(n685), .ZN(n678) );
  NOR2_X1 U736 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U737 ( .A(n681), .B(n680), .ZN(n682) );
  XOR2_X1 U738 ( .A(KEYINPUT52), .B(n682), .Z(n683) );
  NOR2_X1 U739 ( .A1(n684), .A2(n683), .ZN(n689) );
  NOR2_X1 U740 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U741 ( .A(KEYINPUT117), .B(n687), .Z(n688) );
  NOR2_X1 U742 ( .A1(n689), .A2(n688), .ZN(n697) );
  INV_X1 U743 ( .A(n740), .ZN(n690) );
  NOR2_X1 U744 ( .A1(n606), .A2(n690), .ZN(n691) );
  NOR2_X1 U745 ( .A1(n691), .A2(KEYINPUT79), .ZN(n692) );
  XNOR2_X1 U746 ( .A(n692), .B(KEYINPUT2), .ZN(n695) );
  NAND2_X1 U747 ( .A1(n606), .A2(n740), .ZN(n693) );
  NAND2_X1 U748 ( .A1(n693), .A2(KEYINPUT79), .ZN(n694) );
  NAND2_X1 U749 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U750 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U751 ( .A1(n698), .A2(G953), .ZN(n699) );
  XNOR2_X1 U752 ( .A(n699), .B(KEYINPUT53), .ZN(G75) );
  BUF_X2 U753 ( .A(n386), .Z(n713) );
  NAND2_X1 U754 ( .A1(n713), .A2(G469), .ZN(n707) );
  XNOR2_X1 U755 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n701) );
  XNOR2_X1 U756 ( .A(n701), .B(KEYINPUT118), .ZN(n702) );
  XOR2_X1 U757 ( .A(n702), .B(KEYINPUT58), .Z(n703) );
  XNOR2_X1 U758 ( .A(n703), .B(KEYINPUT57), .ZN(n704) );
  XNOR2_X1 U759 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U761 ( .A1(n718), .A2(n708), .ZN(G54) );
  NAND2_X1 U762 ( .A1(n713), .A2(G478), .ZN(n711) );
  XNOR2_X1 U763 ( .A(n709), .B(KEYINPUT121), .ZN(n710) );
  XNOR2_X1 U764 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U765 ( .A1(n718), .A2(n712), .ZN(G63) );
  NAND2_X1 U766 ( .A1(n713), .A2(G217), .ZN(n716) );
  XNOR2_X1 U767 ( .A(n714), .B(KEYINPUT122), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n718), .A2(n717), .ZN(G66) );
  INV_X1 U770 ( .A(n719), .ZN(n722) );
  BUF_X1 U771 ( .A(n720), .Z(n721) );
  NOR2_X1 U772 ( .A1(n722), .A2(n721), .ZN(n730) );
  NOR2_X1 U773 ( .A1(n606), .A2(G953), .ZN(n727) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n723) );
  XOR2_X1 U775 ( .A(KEYINPUT61), .B(n723), .Z(n724) );
  NOR2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U777 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U778 ( .A(n728), .B(KEYINPUT123), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(G69) );
  XOR2_X1 U780 ( .A(n732), .B(n731), .Z(n733) );
  XNOR2_X1 U781 ( .A(KEYINPUT124), .B(n733), .ZN(n734) );
  XOR2_X1 U782 ( .A(n735), .B(n734), .Z(n739) );
  XNOR2_X1 U783 ( .A(n739), .B(G227), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U785 ( .A1(G953), .A2(n737), .ZN(n738) );
  XOR2_X1 U786 ( .A(KEYINPUT126), .B(n738), .Z(n744) );
  XNOR2_X1 U787 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U788 ( .A1(G953), .A2(n741), .ZN(n742) );
  XOR2_X1 U789 ( .A(KEYINPUT125), .B(n742), .Z(n743) );
  NOR2_X1 U790 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U791 ( .A(KEYINPUT127), .B(n745), .ZN(G72) );
  XOR2_X1 U792 ( .A(G140), .B(n746), .Z(G42) );
  XOR2_X1 U793 ( .A(n747), .B(G101), .Z(G3) );
  BUF_X1 U794 ( .A(n748), .Z(n749) );
  XNOR2_X1 U795 ( .A(n749), .B(n390), .ZN(G21) );
  XOR2_X1 U796 ( .A(n750), .B(G131), .Z(G33) );
  XOR2_X1 U797 ( .A(G137), .B(n751), .Z(G39) );
endmodule

