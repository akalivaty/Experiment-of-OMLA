

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U556 ( .A1(n611), .A2(n610), .ZN(n1018) );
  INV_X1 U557 ( .A(n669), .ZN(n648) );
  NOR2_X2 U558 ( .A1(n528), .A2(G2105), .ZN(n524) );
  NOR2_X2 U559 ( .A1(n609), .A2(n608), .ZN(n611) );
  NOR2_X1 U560 ( .A1(n1018), .A2(n617), .ZN(n618) );
  XNOR2_X1 U561 ( .A(G2104), .B(KEYINPUT67), .ZN(n528) );
  OR2_X2 U562 ( .A1(n756), .A2(n755), .ZN(n770) );
  BUF_X1 U563 ( .A(n653), .Z(n669) );
  NOR2_X1 U564 ( .A1(n661), .A2(n660), .ZN(n663) );
  INV_X1 U565 ( .A(KEYINPUT107), .ZN(n721) );
  XOR2_X1 U566 ( .A(G543), .B(KEYINPUT0), .Z(n584) );
  NOR2_X2 U567 ( .A1(n541), .A2(n540), .ZN(G160) );
  NOR2_X1 U568 ( .A1(n715), .A2(n684), .ZN(n521) );
  NOR2_X1 U569 ( .A1(n634), .A2(n633), .ZN(n635) );
  INV_X1 U570 ( .A(KEYINPUT31), .ZN(n662) );
  XNOR2_X1 U571 ( .A(n663), .B(n662), .ZN(n664) );
  INV_X1 U572 ( .A(KEYINPUT99), .ZN(n666) );
  XNOR2_X1 U573 ( .A(n667), .B(n666), .ZN(n678) );
  AND2_X1 U574 ( .A1(n702), .A2(n691), .ZN(n690) );
  INV_X1 U575 ( .A(KEYINPUT106), .ZN(n711) );
  INV_X1 U576 ( .A(KEYINPUT75), .ZN(n602) );
  XNOR2_X1 U577 ( .A(n602), .B(KEYINPUT12), .ZN(n603) );
  XNOR2_X1 U578 ( .A(n604), .B(n603), .ZN(n606) );
  NOR2_X1 U579 ( .A1(G164), .A2(G1384), .ZN(n742) );
  INV_X1 U580 ( .A(G651), .ZN(n546) );
  NAND2_X1 U581 ( .A1(n754), .A2(n763), .ZN(n755) );
  NOR2_X1 U582 ( .A1(G651), .A2(G543), .ZN(n803) );
  INV_X1 U583 ( .A(KEYINPUT23), .ZN(n536) );
  XNOR2_X1 U584 ( .A(KEYINPUT66), .B(n543), .ZN(n800) );
  XNOR2_X1 U585 ( .A(KEYINPUT70), .B(n548), .ZN(n799) );
  XNOR2_X1 U586 ( .A(n537), .B(n536), .ZN(n539) );
  XNOR2_X1 U587 ( .A(KEYINPUT17), .B(KEYINPUT69), .ZN(n523) );
  NOR2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n892) );
  NAND2_X1 U590 ( .A1(n892), .A2(G138), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n524), .B(KEYINPUT68), .ZN(n535) );
  INV_X1 U592 ( .A(n535), .ZN(n525) );
  INV_X2 U593 ( .A(n525), .ZN(n893) );
  NAND2_X1 U594 ( .A1(G102), .A2(n893), .ZN(n526) );
  NAND2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n532) );
  AND2_X1 U596 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  NAND2_X1 U597 ( .A1(G114), .A2(n897), .ZN(n530) );
  AND2_X1 U598 ( .A1(n528), .A2(G2105), .ZN(n900) );
  NAND2_X1 U599 ( .A1(G126), .A2(n900), .ZN(n529) );
  NAND2_X1 U600 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U601 ( .A1(n532), .A2(n531), .ZN(G164) );
  NAND2_X1 U602 ( .A1(G137), .A2(n892), .ZN(n534) );
  NAND2_X1 U603 ( .A1(G113), .A2(n897), .ZN(n533) );
  NAND2_X1 U604 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND2_X1 U605 ( .A1(n535), .A2(G101), .ZN(n537) );
  NAND2_X1 U606 ( .A1(n900), .A2(G125), .ZN(n538) );
  NAND2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U608 ( .A1(G91), .A2(n803), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n542), .B(KEYINPUT72), .ZN(n553) );
  NOR2_X1 U610 ( .A1(n584), .A2(n546), .ZN(n805) );
  NAND2_X1 U611 ( .A1(G78), .A2(n805), .ZN(n545) );
  NOR2_X1 U612 ( .A1(G651), .A2(n584), .ZN(n543) );
  NAND2_X1 U613 ( .A1(G53), .A2(n800), .ZN(n544) );
  NAND2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n551) );
  NOR2_X1 U615 ( .A1(G543), .A2(n546), .ZN(n547) );
  XOR2_X1 U616 ( .A(KEYINPUT1), .B(n547), .Z(n548) );
  NAND2_X1 U617 ( .A1(G65), .A2(n799), .ZN(n549) );
  XNOR2_X1 U618 ( .A(KEYINPUT73), .B(n549), .ZN(n550) );
  NOR2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(G299) );
  NAND2_X1 U621 ( .A1(G90), .A2(n803), .ZN(n555) );
  NAND2_X1 U622 ( .A1(G77), .A2(n805), .ZN(n554) );
  NAND2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT9), .ZN(n558) );
  NAND2_X1 U625 ( .A1(G64), .A2(n799), .ZN(n557) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U627 ( .A1(G52), .A2(n800), .ZN(n559) );
  XNOR2_X1 U628 ( .A(KEYINPUT71), .B(n559), .ZN(n560) );
  NOR2_X1 U629 ( .A1(n561), .A2(n560), .ZN(G171) );
  NAND2_X1 U630 ( .A1(n803), .A2(G89), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U632 ( .A1(G76), .A2(n805), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U634 ( .A(KEYINPUT5), .B(n565), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G63), .A2(n799), .ZN(n566) );
  XOR2_X1 U636 ( .A(KEYINPUT79), .B(n566), .Z(n568) );
  NAND2_X1 U637 ( .A1(G51), .A2(n800), .ZN(n567) );
  NAND2_X1 U638 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U639 ( .A(KEYINPUT6), .B(n569), .Z(n570) );
  NAND2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U641 ( .A(KEYINPUT7), .B(n572), .ZN(G168) );
  XOR2_X1 U642 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U643 ( .A1(G88), .A2(n803), .ZN(n574) );
  NAND2_X1 U644 ( .A1(G75), .A2(n805), .ZN(n573) );
  NAND2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G62), .A2(n799), .ZN(n576) );
  NAND2_X1 U647 ( .A1(G50), .A2(n800), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U649 ( .A1(n578), .A2(n577), .ZN(G166) );
  INV_X1 U650 ( .A(G166), .ZN(G303) );
  NAND2_X1 U651 ( .A1(n800), .A2(G49), .ZN(n579) );
  XNOR2_X1 U652 ( .A(n579), .B(KEYINPUT84), .ZN(n582) );
  NAND2_X1 U653 ( .A1(G74), .A2(G651), .ZN(n580) );
  XOR2_X1 U654 ( .A(KEYINPUT85), .B(n580), .Z(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U656 ( .A1(n799), .A2(n583), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n584), .A2(G87), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(G288) );
  NAND2_X1 U659 ( .A1(n803), .A2(G86), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G61), .A2(n799), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U662 ( .A(KEYINPUT86), .B(n589), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n805), .A2(G73), .ZN(n590) );
  XOR2_X1 U664 ( .A(KEYINPUT2), .B(n590), .Z(n591) );
  NOR2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G48), .A2(n800), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(G305) );
  NAND2_X1 U668 ( .A1(G85), .A2(n803), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G72), .A2(n805), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G60), .A2(n799), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G47), .A2(n800), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  OR2_X1 U674 ( .A1(n600), .A2(n599), .ZN(G290) );
  NAND2_X1 U675 ( .A1(n799), .A2(G56), .ZN(n601) );
  XOR2_X1 U676 ( .A(KEYINPUT14), .B(n601), .Z(n609) );
  NAND2_X1 U677 ( .A1(G81), .A2(n803), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G68), .A2(n805), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U680 ( .A(KEYINPUT13), .B(n607), .Z(n608) );
  NAND2_X1 U681 ( .A1(G43), .A2(n800), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G160), .A2(G40), .ZN(n741) );
  INV_X1 U683 ( .A(n741), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n612), .A2(n742), .ZN(n653) );
  INV_X1 U685 ( .A(G1996), .ZN(n985) );
  NOR2_X1 U686 ( .A1(n653), .A2(n985), .ZN(n614) );
  XOR2_X1 U687 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n613) );
  XNOR2_X1 U688 ( .A(n614), .B(n613), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n669), .A2(G1341), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n618), .B(KEYINPUT65), .ZN(n631) );
  NAND2_X1 U692 ( .A1(n803), .A2(G92), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G66), .A2(n799), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U695 ( .A1(G79), .A2(n805), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G54), .A2(n800), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n626) );
  XNOR2_X1 U699 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X2 U701 ( .A(KEYINPUT15), .B(n627), .ZN(n908) );
  INV_X1 U702 ( .A(G1348), .ZN(n1011) );
  NOR2_X1 U703 ( .A1(n648), .A2(n1011), .ZN(n629) );
  AND2_X1 U704 ( .A1(n648), .A2(G2067), .ZN(n628) );
  NOR2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n632) );
  NOR2_X1 U706 ( .A1(n908), .A2(n632), .ZN(n630) );
  NOR2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n634) );
  AND2_X1 U708 ( .A1(n908), .A2(n632), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n635), .B(KEYINPUT96), .ZN(n640) );
  NAND2_X1 U710 ( .A1(n648), .A2(G2072), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(KEYINPUT27), .ZN(n638) );
  INV_X1 U712 ( .A(G1956), .ZN(n958) );
  NOR2_X1 U713 ( .A1(n958), .A2(n648), .ZN(n637) );
  NOR2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n641) );
  INV_X1 U715 ( .A(G299), .ZN(n812) );
  NAND2_X1 U716 ( .A1(n641), .A2(n812), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n644) );
  NOR2_X1 U718 ( .A1(n641), .A2(n812), .ZN(n642) );
  XOR2_X1 U719 ( .A(n642), .B(KEYINPUT28), .Z(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X1 U721 ( .A(KEYINPUT29), .B(KEYINPUT97), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n646), .B(n645), .ZN(n652) );
  NOR2_X1 U723 ( .A1(n648), .A2(G1961), .ZN(n647) );
  XNOR2_X1 U724 ( .A(n647), .B(KEYINPUT95), .ZN(n650) );
  XNOR2_X1 U725 ( .A(G2078), .B(KEYINPUT25), .ZN(n984) );
  NAND2_X1 U726 ( .A1(n648), .A2(n984), .ZN(n649) );
  NAND2_X1 U727 ( .A1(n650), .A2(n649), .ZN(n659) );
  NAND2_X1 U728 ( .A1(n659), .A2(G171), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n665) );
  NAND2_X1 U730 ( .A1(G8), .A2(n653), .ZN(n715) );
  NOR2_X1 U731 ( .A1(G1966), .A2(n715), .ZN(n654) );
  XOR2_X1 U732 ( .A(KEYINPUT94), .B(n654), .Z(n681) );
  INV_X1 U733 ( .A(G8), .ZN(n674) );
  NOR2_X1 U734 ( .A1(G2084), .A2(n669), .ZN(n679) );
  NOR2_X1 U735 ( .A1(n674), .A2(n679), .ZN(n655) );
  AND2_X1 U736 ( .A1(n681), .A2(n655), .ZN(n657) );
  XOR2_X1 U737 ( .A(KEYINPUT98), .B(KEYINPUT30), .Z(n656) );
  XNOR2_X1 U738 ( .A(n657), .B(n656), .ZN(n658) );
  NOR2_X1 U739 ( .A1(G168), .A2(n658), .ZN(n661) );
  NOR2_X1 U740 ( .A1(G171), .A2(n659), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n665), .A2(n664), .ZN(n667) );
  AND2_X1 U742 ( .A1(G286), .A2(G8), .ZN(n668) );
  NAND2_X1 U743 ( .A1(n678), .A2(n668), .ZN(n676) );
  NOR2_X1 U744 ( .A1(G1971), .A2(n715), .ZN(n671) );
  NOR2_X1 U745 ( .A1(G2090), .A2(n669), .ZN(n670) );
  NOR2_X1 U746 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n672), .A2(G303), .ZN(n673) );
  OR2_X1 U748 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U749 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X2 U750 ( .A(n677), .B(KEYINPUT32), .ZN(n704) );
  XNOR2_X1 U751 ( .A(n678), .B(KEYINPUT100), .ZN(n683) );
  NAND2_X1 U752 ( .A1(G8), .A2(n679), .ZN(n680) );
  AND2_X1 U753 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U754 ( .A1(n683), .A2(n682), .ZN(n702) );
  NAND2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n1021) );
  INV_X1 U756 ( .A(n1021), .ZN(n684) );
  NOR2_X1 U757 ( .A1(KEYINPUT33), .A2(n521), .ZN(n689) );
  NOR2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n685) );
  XOR2_X1 U759 ( .A(KEYINPUT101), .B(n685), .Z(n693) );
  NAND2_X1 U760 ( .A1(n693), .A2(KEYINPUT33), .ZN(n686) );
  XOR2_X1 U761 ( .A(KEYINPUT103), .B(n686), .Z(n687) );
  NOR2_X1 U762 ( .A1(n715), .A2(n687), .ZN(n688) );
  NOR2_X1 U763 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U764 ( .A1(n704), .A2(n690), .ZN(n699) );
  INV_X1 U765 ( .A(n691), .ZN(n697) );
  NOR2_X1 U766 ( .A1(G1971), .A2(G303), .ZN(n692) );
  NOR2_X1 U767 ( .A1(n693), .A2(n692), .ZN(n1030) );
  XNOR2_X1 U768 ( .A(KEYINPUT102), .B(n1030), .ZN(n695) );
  INV_X1 U769 ( .A(KEYINPUT33), .ZN(n694) );
  AND2_X1 U770 ( .A1(n695), .A2(n694), .ZN(n696) );
  OR2_X1 U771 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U772 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U773 ( .A(n700), .B(KEYINPUT104), .ZN(n701) );
  XOR2_X1 U774 ( .A(G1981), .B(G305), .Z(n1027) );
  AND2_X1 U775 ( .A1(n701), .A2(n1027), .ZN(n720) );
  AND2_X1 U776 ( .A1(n702), .A2(n715), .ZN(n703) );
  NAND2_X1 U777 ( .A1(n704), .A2(n703), .ZN(n710) );
  INV_X1 U778 ( .A(n715), .ZN(n708) );
  NAND2_X1 U779 ( .A1(G8), .A2(G166), .ZN(n705) );
  NOR2_X1 U780 ( .A1(G2090), .A2(n705), .ZN(n706) );
  XNOR2_X1 U781 ( .A(n706), .B(KEYINPUT105), .ZN(n707) );
  OR2_X1 U782 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U783 ( .A1(n710), .A2(n709), .ZN(n712) );
  XNOR2_X1 U784 ( .A(n712), .B(n711), .ZN(n718) );
  NOR2_X1 U785 ( .A1(G1981), .A2(G305), .ZN(n713) );
  XNOR2_X1 U786 ( .A(n713), .B(KEYINPUT24), .ZN(n714) );
  XNOR2_X1 U787 ( .A(n714), .B(KEYINPUT93), .ZN(n716) );
  OR2_X1 U788 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U789 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n722) );
  XNOR2_X1 U791 ( .A(n722), .B(n721), .ZN(n756) );
  NAND2_X1 U792 ( .A1(G141), .A2(n892), .ZN(n724) );
  NAND2_X1 U793 ( .A1(G117), .A2(n897), .ZN(n723) );
  NAND2_X1 U794 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U795 ( .A1(n893), .A2(G105), .ZN(n725) );
  XOR2_X1 U796 ( .A(KEYINPUT38), .B(n725), .Z(n726) );
  NOR2_X1 U797 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n900), .A2(G129), .ZN(n728) );
  NAND2_X1 U799 ( .A1(n729), .A2(n728), .ZN(n876) );
  NAND2_X1 U800 ( .A1(G1996), .A2(n876), .ZN(n730) );
  XOR2_X1 U801 ( .A(KEYINPUT92), .B(n730), .Z(n740) );
  NAND2_X1 U802 ( .A1(G107), .A2(n897), .ZN(n737) );
  NAND2_X1 U803 ( .A1(n892), .A2(G131), .ZN(n732) );
  NAND2_X1 U804 ( .A1(G95), .A2(n893), .ZN(n731) );
  NAND2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n735) );
  NAND2_X1 U806 ( .A1(n900), .A2(G119), .ZN(n733) );
  XOR2_X1 U807 ( .A(KEYINPUT90), .B(n733), .Z(n734) );
  NOR2_X1 U808 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U810 ( .A(n738), .B(KEYINPUT91), .Z(n873) );
  AND2_X1 U811 ( .A1(n873), .A2(G1991), .ZN(n739) );
  NOR2_X1 U812 ( .A1(n740), .A2(n739), .ZN(n937) );
  XOR2_X1 U813 ( .A(G1986), .B(G290), .Z(n1017) );
  NAND2_X1 U814 ( .A1(n937), .A2(n1017), .ZN(n743) );
  NOR2_X1 U815 ( .A1(n742), .A2(n741), .ZN(n767) );
  NAND2_X1 U816 ( .A1(n743), .A2(n767), .ZN(n754) );
  NAND2_X1 U817 ( .A1(n892), .A2(G140), .ZN(n745) );
  NAND2_X1 U818 ( .A1(G104), .A2(n893), .ZN(n744) );
  NAND2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U820 ( .A(KEYINPUT34), .B(n746), .ZN(n752) );
  NAND2_X1 U821 ( .A1(n900), .A2(G128), .ZN(n747) );
  XOR2_X1 U822 ( .A(KEYINPUT89), .B(n747), .Z(n749) );
  NAND2_X1 U823 ( .A1(n897), .A2(G116), .ZN(n748) );
  NAND2_X1 U824 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U825 ( .A(KEYINPUT35), .B(n750), .Z(n751) );
  NOR2_X1 U826 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U827 ( .A(KEYINPUT36), .B(n753), .ZN(n872) );
  XNOR2_X1 U828 ( .A(KEYINPUT37), .B(G2067), .ZN(n765) );
  NOR2_X1 U829 ( .A1(n872), .A2(n765), .ZN(n932) );
  NAND2_X1 U830 ( .A1(n767), .A2(n932), .ZN(n763) );
  INV_X1 U831 ( .A(n937), .ZN(n759) );
  NOR2_X1 U832 ( .A1(G1991), .A2(n873), .ZN(n939) );
  NOR2_X1 U833 ( .A1(G1986), .A2(G290), .ZN(n757) );
  NOR2_X1 U834 ( .A1(n939), .A2(n757), .ZN(n758) );
  NOR2_X1 U835 ( .A1(n759), .A2(n758), .ZN(n761) );
  NOR2_X1 U836 ( .A1(n876), .A2(G1996), .ZN(n760) );
  XNOR2_X1 U837 ( .A(n760), .B(KEYINPUT108), .ZN(n947) );
  NOR2_X1 U838 ( .A1(n761), .A2(n947), .ZN(n762) );
  XNOR2_X1 U839 ( .A(KEYINPUT39), .B(n762), .ZN(n764) );
  NAND2_X1 U840 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U841 ( .A1(n872), .A2(n765), .ZN(n931) );
  NAND2_X1 U842 ( .A1(n766), .A2(n931), .ZN(n768) );
  NAND2_X1 U843 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U844 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U845 ( .A(n771), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U846 ( .A(G171), .ZN(G301) );
  AND2_X1 U847 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U848 ( .A(G132), .ZN(G219) );
  INV_X1 U849 ( .A(G82), .ZN(G220) );
  INV_X1 U850 ( .A(G57), .ZN(G237) );
  NAND2_X1 U851 ( .A1(G7), .A2(G661), .ZN(n772) );
  XNOR2_X1 U852 ( .A(n772), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U853 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n774) );
  INV_X1 U854 ( .A(G223), .ZN(n837) );
  NAND2_X1 U855 ( .A1(G567), .A2(n837), .ZN(n773) );
  XNOR2_X1 U856 ( .A(n774), .B(n773), .ZN(G234) );
  INV_X1 U857 ( .A(G860), .ZN(n798) );
  OR2_X1 U858 ( .A1(n1018), .A2(n798), .ZN(G153) );
  INV_X1 U859 ( .A(G868), .ZN(n778) );
  NOR2_X1 U860 ( .A1(G301), .A2(n778), .ZN(n776) );
  INV_X1 U861 ( .A(n908), .ZN(n1010) );
  NOR2_X1 U862 ( .A1(n1010), .A2(G868), .ZN(n775) );
  NOR2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U864 ( .A(KEYINPUT78), .B(n777), .ZN(G284) );
  NOR2_X1 U865 ( .A1(G286), .A2(n778), .ZN(n780) );
  NOR2_X1 U866 ( .A1(G868), .A2(G299), .ZN(n779) );
  NOR2_X1 U867 ( .A1(n780), .A2(n779), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n798), .A2(G559), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n781), .A2(n908), .ZN(n782) );
  XNOR2_X1 U870 ( .A(n782), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U871 ( .A1(G868), .A2(n1018), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n908), .A2(G868), .ZN(n783) );
  NOR2_X1 U873 ( .A1(G559), .A2(n783), .ZN(n784) );
  NOR2_X1 U874 ( .A1(n785), .A2(n784), .ZN(G282) );
  NAND2_X1 U875 ( .A1(n897), .A2(G111), .ZN(n786) );
  XNOR2_X1 U876 ( .A(n786), .B(KEYINPUT80), .ZN(n788) );
  NAND2_X1 U877 ( .A1(G99), .A2(n893), .ZN(n787) );
  NAND2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U879 ( .A(n789), .B(KEYINPUT81), .ZN(n791) );
  NAND2_X1 U880 ( .A1(G135), .A2(n892), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n900), .A2(G123), .ZN(n792) );
  XOR2_X1 U883 ( .A(KEYINPUT18), .B(n792), .Z(n793) );
  NOR2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n935) );
  XNOR2_X1 U885 ( .A(n935), .B(G2096), .ZN(n796) );
  INV_X1 U886 ( .A(G2100), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(G156) );
  NAND2_X1 U888 ( .A1(n908), .A2(G559), .ZN(n797) );
  XOR2_X1 U889 ( .A(n1018), .B(n797), .Z(n819) );
  NAND2_X1 U890 ( .A1(n798), .A2(n819), .ZN(n811) );
  NAND2_X1 U891 ( .A1(G67), .A2(n799), .ZN(n802) );
  NAND2_X1 U892 ( .A1(G55), .A2(n800), .ZN(n801) );
  NAND2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n810) );
  NAND2_X1 U894 ( .A1(n803), .A2(G93), .ZN(n804) );
  XNOR2_X1 U895 ( .A(n804), .B(KEYINPUT82), .ZN(n807) );
  NAND2_X1 U896 ( .A1(G80), .A2(n805), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U898 ( .A(KEYINPUT83), .B(n808), .Z(n809) );
  NOR2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n821) );
  XOR2_X1 U900 ( .A(n811), .B(n821), .Z(G145) );
  XNOR2_X1 U901 ( .A(n812), .B(G290), .ZN(n818) );
  XNOR2_X1 U902 ( .A(KEYINPUT87), .B(KEYINPUT19), .ZN(n814) );
  XNOR2_X1 U903 ( .A(G305), .B(G166), .ZN(n813) );
  XNOR2_X1 U904 ( .A(n814), .B(n813), .ZN(n815) );
  XNOR2_X1 U905 ( .A(n821), .B(n815), .ZN(n816) );
  XNOR2_X1 U906 ( .A(n816), .B(G288), .ZN(n817) );
  XNOR2_X1 U907 ( .A(n818), .B(n817), .ZN(n910) );
  XNOR2_X1 U908 ( .A(n819), .B(n910), .ZN(n820) );
  NAND2_X1 U909 ( .A1(n820), .A2(G868), .ZN(n823) );
  OR2_X1 U910 ( .A1(G868), .A2(n821), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n823), .A2(n822), .ZN(G295) );
  NAND2_X1 U912 ( .A1(G2084), .A2(G2078), .ZN(n824) );
  XOR2_X1 U913 ( .A(KEYINPUT20), .B(n824), .Z(n825) );
  NAND2_X1 U914 ( .A1(G2090), .A2(n825), .ZN(n826) );
  XNOR2_X1 U915 ( .A(KEYINPUT21), .B(n826), .ZN(n827) );
  NAND2_X1 U916 ( .A1(n827), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U917 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U918 ( .A1(G69), .A2(G120), .ZN(n828) );
  NOR2_X1 U919 ( .A1(G237), .A2(n828), .ZN(n829) );
  NAND2_X1 U920 ( .A1(G108), .A2(n829), .ZN(n843) );
  NAND2_X1 U921 ( .A1(n843), .A2(G567), .ZN(n835) );
  NOR2_X1 U922 ( .A1(G220), .A2(G219), .ZN(n830) );
  XOR2_X1 U923 ( .A(KEYINPUT22), .B(n830), .Z(n831) );
  NOR2_X1 U924 ( .A1(G218), .A2(n831), .ZN(n832) );
  NAND2_X1 U925 ( .A1(G96), .A2(n832), .ZN(n842) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n842), .ZN(n833) );
  XNOR2_X1 U927 ( .A(KEYINPUT88), .B(n833), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n844) );
  NAND2_X1 U929 ( .A1(G483), .A2(G661), .ZN(n836) );
  NOR2_X1 U930 ( .A1(n844), .A2(n836), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U934 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U937 ( .A(KEYINPUT111), .B(n841), .Z(G188) );
  XOR2_X1 U938 ( .A(G96), .B(KEYINPUT112), .Z(G221) );
  INV_X1 U940 ( .A(G120), .ZN(G236) );
  INV_X1 U941 ( .A(G69), .ZN(G235) );
  NOR2_X1 U942 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U943 ( .A(G325), .ZN(G261) );
  INV_X1 U944 ( .A(n844), .ZN(G319) );
  XOR2_X1 U945 ( .A(KEYINPUT42), .B(G2078), .Z(n846) );
  XNOR2_X1 U946 ( .A(G2084), .B(G2072), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U948 ( .A(n847), .B(G2100), .Z(n849) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2090), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(G2096), .B(KEYINPUT43), .Z(n851) );
  XNOR2_X1 U952 ( .A(KEYINPUT113), .B(G2678), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U954 ( .A(n853), .B(n852), .Z(G227) );
  XOR2_X1 U955 ( .A(G2474), .B(G1961), .Z(n855) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1956), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U958 ( .A(n856), .B(KEYINPUT114), .Z(n858) );
  XNOR2_X1 U959 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U961 ( .A(G1971), .B(G1966), .Z(n860) );
  XNOR2_X1 U962 ( .A(G1981), .B(G1976), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U964 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U965 ( .A(KEYINPUT115), .B(KEYINPUT41), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U967 ( .A1(G124), .A2(n900), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n897), .A2(G112), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n892), .A2(G136), .ZN(n869) );
  NAND2_X1 U972 ( .A1(G100), .A2(n893), .ZN(n868) );
  NAND2_X1 U973 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(G162) );
  XNOR2_X1 U975 ( .A(n935), .B(n872), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U977 ( .A(G160), .B(G162), .Z(n875) );
  XNOR2_X1 U978 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U979 ( .A(n878), .B(n877), .Z(n883) );
  XOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n880) );
  XNOR2_X1 U981 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U983 ( .A(G164), .B(n881), .ZN(n882) );
  XNOR2_X1 U984 ( .A(n883), .B(n882), .ZN(n906) );
  NAND2_X1 U985 ( .A1(n892), .A2(G139), .ZN(n885) );
  NAND2_X1 U986 ( .A1(G103), .A2(n893), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n890) );
  NAND2_X1 U988 ( .A1(G115), .A2(n897), .ZN(n887) );
  NAND2_X1 U989 ( .A1(G127), .A2(n900), .ZN(n886) );
  NAND2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U993 ( .A(KEYINPUT117), .B(n891), .Z(n942) );
  NAND2_X1 U994 ( .A1(n892), .A2(G142), .ZN(n895) );
  NAND2_X1 U995 ( .A1(G106), .A2(n893), .ZN(n894) );
  NAND2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n896), .B(KEYINPUT45), .ZN(n899) );
  NAND2_X1 U998 ( .A1(G118), .A2(n897), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n903) );
  NAND2_X1 U1000 ( .A1(n900), .A2(G130), .ZN(n901) );
  XOR2_X1 U1001 ( .A(KEYINPUT116), .B(n901), .Z(n902) );
  NOR2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n942), .B(n904), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n907), .ZN(G395) );
  XNOR2_X1 U1006 ( .A(G286), .B(n908), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n909), .B(n1018), .ZN(n912) );
  XOR2_X1 U1008 ( .A(G301), .B(n910), .Z(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n913), .ZN(G397) );
  XNOR2_X1 U1011 ( .A(G2451), .B(G2427), .ZN(n923) );
  XOR2_X1 U1012 ( .A(G2430), .B(G2443), .Z(n915) );
  XNOR2_X1 U1013 ( .A(KEYINPUT109), .B(G2438), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n915), .B(n914), .ZN(n919) );
  XOR2_X1 U1015 ( .A(G2435), .B(G2454), .Z(n917) );
  XNOR2_X1 U1016 ( .A(G1348), .B(G1341), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1018 ( .A(n919), .B(n918), .Z(n921) );
  XNOR2_X1 U1019 ( .A(G2446), .B(KEYINPUT110), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(n921), .B(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n923), .B(n922), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n924), .A2(G14), .ZN(n930) );
  NAND2_X1 U1023 ( .A1(G319), .A2(n930), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(KEYINPUT49), .B(n925), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(G395), .A2(G397), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  INV_X1 U1031 ( .A(n930), .ZN(G401) );
  INV_X1 U1032 ( .A(n931), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n941) );
  XOR2_X1 U1034 ( .A(G2084), .B(G160), .Z(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n952) );
  XOR2_X1 U1039 ( .A(G2072), .B(n942), .Z(n944) );
  XOR2_X1 U1040 ( .A(G164), .B(G2078), .Z(n943) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1042 ( .A(KEYINPUT50), .B(n945), .ZN(n950) );
  XOR2_X1 U1043 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1045 ( .A(KEYINPUT51), .B(n948), .Z(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n953), .ZN(n955) );
  INV_X1 U1049 ( .A(KEYINPUT55), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1051 ( .A1(n956), .A2(G29), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(KEYINPUT120), .B(n957), .ZN(n1009) );
  XOR2_X1 U1053 ( .A(G1961), .B(G5), .Z(n972) );
  XOR2_X1 U1054 ( .A(G1981), .B(G6), .Z(n960) );
  XNOR2_X1 U1055 ( .A(n958), .B(G20), .ZN(n959) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n966) );
  XOR2_X1 U1057 ( .A(G1341), .B(G19), .Z(n964) );
  XNOR2_X1 U1058 ( .A(G4), .B(KEYINPUT125), .ZN(n961) );
  XNOR2_X1 U1059 ( .A(n961), .B(n1011), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(n962), .B(KEYINPUT59), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1063 ( .A(KEYINPUT60), .B(n967), .Z(n969) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G21), .ZN(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(KEYINPUT126), .B(n970), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(G1986), .B(G24), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G22), .B(G1971), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(G1976), .B(KEYINPUT127), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(n975), .B(G23), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(KEYINPUT58), .B(n978), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1076 ( .A(KEYINPUT61), .B(n981), .Z(n982) );
  NOR2_X1 U1077 ( .A1(G16), .A2(n982), .ZN(n1007) );
  XOR2_X1 U1078 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n1002) );
  XNOR2_X1 U1079 ( .A(G2090), .B(G35), .ZN(n997) );
  XOR2_X1 U1080 ( .A(G2072), .B(G33), .Z(n983) );
  NAND2_X1 U1081 ( .A1(n983), .A2(G28), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(n984), .B(G27), .ZN(n987) );
  XNOR2_X1 U1083 ( .A(n985), .B(G32), .ZN(n986) );
  NAND2_X1 U1084 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1085 ( .A(KEYINPUT121), .B(n988), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(G2067), .B(G26), .ZN(n990) );
  XNOR2_X1 U1087 ( .A(G1991), .B(G25), .ZN(n989) );
  NOR2_X1 U1088 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1089 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1090 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1091 ( .A(KEYINPUT53), .B(n995), .ZN(n996) );
  NOR2_X1 U1092 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1093 ( .A(G2084), .B(G34), .Z(n998) );
  XNOR2_X1 U1094 ( .A(KEYINPUT54), .B(n998), .ZN(n999) );
  NAND2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1096 ( .A(n1002), .B(n1001), .ZN(n1004) );
  INV_X1 U1097 ( .A(G29), .ZN(n1003) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1099 ( .A1(G11), .A2(n1005), .ZN(n1006) );
  NOR2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1037) );
  XOR2_X1 U1102 ( .A(KEYINPUT56), .B(G16), .Z(n1035) );
  XNOR2_X1 U1103 ( .A(n1010), .B(KEYINPUT123), .ZN(n1012) );
  XNOR2_X1 U1104 ( .A(n1012), .B(n1011), .ZN(n1014) );
  XNOR2_X1 U1105 ( .A(G1961), .B(G301), .ZN(n1013) );
  NOR2_X1 U1106 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1107 ( .A(KEYINPUT124), .B(n1015), .ZN(n1026) );
  NAND2_X1 U1108 ( .A1(G1971), .A2(G303), .ZN(n1016) );
  NAND2_X1 U1109 ( .A1(n1017), .A2(n1016), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(G299), .B(G1956), .ZN(n1020) );
  XNOR2_X1 U1111 ( .A(n1018), .B(G1341), .ZN(n1019) );
  NOR2_X1 U1112 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  NAND2_X1 U1113 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(G1966), .B(G168), .ZN(n1028) );
  NAND2_X1 U1117 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1118 ( .A(n1029), .B(KEYINPUT57), .ZN(n1031) );
  NAND2_X1 U1119 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1120 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1122 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1123 ( .A(n1038), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

