//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(new_n202), .A2(new_n203), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G20), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  INV_X1    g0016(.A(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(G250), .B1(G257), .B2(G264), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n214), .B1(new_n220), .B2(KEYINPUT0), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  INV_X1    g0028(.A(G87), .ZN(new_n229));
  INV_X1    g0029(.A(G250), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n233));
  INV_X1    g0033(.A(KEYINPUT66), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G68), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(G238), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(KEYINPUT67), .ZN(new_n238));
  INV_X1    g0038(.A(KEYINPUT67), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G238), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g0041(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g0042(.A(new_n216), .B1(new_n232), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  AOI211_X1 g0045(.A(new_n221), .B(new_n245), .C1(KEYINPUT0), .C2(new_n220), .ZN(G361));
  XNOR2_X1  g0046(.A(G238), .B(G244), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G232), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT2), .B(G226), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G250), .B(G257), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G270), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT69), .B(G264), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n250), .B(new_n254), .ZN(G358));
  XOR2_X1   g0055(.A(G50), .B(G68), .Z(new_n256));
  XNOR2_X1  g0056(.A(G58), .B(G77), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(G87), .B(G116), .ZN(new_n259));
  XNOR2_X1  g0059(.A(G97), .B(G107), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n258), .B(new_n261), .Z(G351));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G222), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G223), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n270), .A3(G1698), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n265), .B1(new_n223), .B2(new_n263), .C1(new_n266), .C2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n211), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G41), .B2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(G1), .B(G13), .C1(new_n267), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n277), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n279), .B1(new_n283), .B2(G226), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n275), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g0085(.A(KEYINPUT72), .B(G200), .Z(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G190), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(new_n285), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n211), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n291), .A2(KEYINPUT70), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(KEYINPUT70), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n204), .A2(G20), .ZN(new_n295));
  INV_X1    g0095(.A(G150), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(KEYINPUT8), .A2(G58), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT8), .A2(G58), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n267), .A2(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n295), .B1(new_n296), .B2(new_n298), .C1(new_n301), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n276), .A2(G20), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n217), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n294), .A2(new_n304), .B1(new_n201), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n292), .A2(new_n293), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(G50), .A3(new_n305), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n307), .A2(KEYINPUT9), .A3(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n289), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT10), .B1(new_n289), .B2(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n285), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n310), .B1(new_n320), .B2(G169), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n285), .A2(G179), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G107), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n271), .A2(new_n241), .B1(new_n263), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n268), .A2(new_n270), .ZN(new_n327));
  INV_X1    g0127(.A(G232), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n327), .A2(new_n328), .A3(G1698), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n274), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n279), .B1(new_n283), .B2(G244), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n306), .A2(new_n223), .ZN(new_n335));
  INV_X1    g0135(.A(new_n291), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n305), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n335), .B1(new_n337), .B2(new_n223), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n299), .A2(new_n297), .A3(new_n300), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G20), .A2(G77), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n340), .A2(KEYINPUT71), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT71), .B1(new_n340), .B2(new_n341), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT15), .B(G87), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n303), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n339), .B1(new_n346), .B2(new_n336), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n334), .A2(new_n347), .A3(KEYINPUT73), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT73), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n340), .A2(new_n341), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT71), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n340), .A2(KEYINPUT71), .A3(new_n341), .ZN(new_n353));
  INV_X1    g0153(.A(new_n345), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n338), .B1(new_n355), .B2(new_n291), .ZN(new_n356));
  AOI21_X1  g0156(.A(G169), .B1(new_n330), .B2(new_n331), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n349), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n332), .A2(G179), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n348), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n332), .A2(new_n286), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n330), .A2(G190), .A3(new_n331), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(new_n356), .ZN(new_n364));
  AND4_X1   g0164(.A1(new_n319), .A2(new_n324), .A3(new_n361), .A4(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n302), .A2(G77), .B1(new_n297), .B2(G50), .ZN(new_n366));
  INV_X1    g0166(.A(new_n236), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(new_n212), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n294), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g0169(.A(new_n369), .B(KEYINPUT11), .Z(new_n370));
  INV_X1    g0170(.A(KEYINPUT12), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n306), .B2(new_n236), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT75), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n306), .A2(new_n371), .A3(new_n203), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n373), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n203), .B2(new_n337), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n279), .B1(new_n283), .B2(G238), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n263), .A2(G232), .A3(G1698), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n263), .A2(G226), .A3(new_n264), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n384), .A2(KEYINPUT74), .A3(new_n274), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT74), .B1(new_n384), .B2(new_n274), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n380), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT13), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT13), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n389), .B(new_n380), .C1(new_n385), .C2(new_n386), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(G179), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n333), .B1(new_n388), .B2(new_n390), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT14), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI211_X1 g0194(.A(KEYINPUT14), .B(new_n333), .C1(new_n388), .C2(new_n390), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n379), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n388), .A2(G190), .A3(new_n390), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n388), .A2(new_n390), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n378), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n279), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n282), .B2(new_n328), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n263), .A2(G226), .A3(G1698), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n263), .A2(G223), .A3(new_n264), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n404), .B(new_n405), .C1(new_n267), .C2(new_n229), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n403), .B1(new_n406), .B2(new_n274), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(new_n399), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(G190), .B2(new_n407), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n233), .A2(new_n235), .A3(G58), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT76), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT76), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n233), .A2(new_n235), .A3(new_n412), .A4(G58), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n208), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G20), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n297), .A2(G159), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n263), .A2(new_n417), .A3(G20), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT7), .B1(new_n327), .B2(new_n212), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n367), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n415), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT16), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(G68), .B1(new_n418), .B2(new_n419), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n415), .A2(KEYINPUT16), .A3(new_n424), .A4(new_n416), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n291), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n301), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(new_n306), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n308), .A2(new_n305), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(new_n427), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n409), .A2(new_n426), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT17), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n336), .B1(new_n421), .B2(new_n422), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n434), .B2(new_n425), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT17), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n409), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n426), .A2(new_n431), .ZN(new_n438));
  INV_X1    g0238(.A(G179), .ZN(new_n439));
  AOI211_X1 g0239(.A(new_n439), .B(new_n403), .C1(new_n274), .C2(new_n406), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n406), .A2(new_n274), .ZN(new_n441));
  INV_X1    g0241(.A(new_n403), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n333), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n438), .A2(KEYINPUT18), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT18), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n435), .B2(new_n444), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n433), .A2(new_n437), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n365), .A2(new_n401), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT77), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT6), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n260), .A2(new_n452), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n452), .A2(new_n225), .A3(G107), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(G20), .B1(G77), .B2(new_n297), .ZN(new_n457));
  OAI21_X1  g0257(.A(G107), .B1(new_n418), .B2(new_n419), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n336), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n212), .A2(G1), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G13), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G97), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(G1), .B2(new_n267), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n308), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n463), .B1(new_n466), .B2(new_n225), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n451), .B1(new_n459), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n454), .B1(new_n452), .B2(new_n260), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n469), .A2(new_n212), .B1(new_n223), .B2(new_n298), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n417), .B1(new_n263), .B2(G20), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n327), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n325), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n291), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n464), .B1(new_n293), .B2(new_n292), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n462), .B1(new_n475), .B2(G97), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n476), .A3(KEYINPUT77), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n468), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n276), .A2(G45), .ZN(new_n482));
  OAI211_X1 g0282(.A(G257), .B(new_n281), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n276), .A2(G45), .A3(G274), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n480), .B2(new_n479), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT79), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n483), .A2(KEYINPUT79), .A3(new_n486), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n268), .A2(new_n270), .A3(G244), .A4(new_n264), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .A4(new_n264), .ZN(new_n495));
  AND3_X1   g0295(.A1(KEYINPUT78), .A2(G33), .A3(G283), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT78), .B1(G33), .B2(G283), .ZN(new_n497));
  OR2_X1    g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n263), .A2(G250), .A3(G1698), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n494), .A2(new_n495), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n274), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n491), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n487), .B1(new_n500), .B2(new_n274), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n502), .A2(G200), .B1(G190), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n489), .A2(new_n490), .B1(new_n274), .B2(new_n500), .ZN(new_n505));
  INV_X1    g0305(.A(new_n487), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n505), .A2(new_n439), .B1(new_n507), .B2(new_n333), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n474), .A2(new_n476), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n478), .A2(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n482), .B1(new_n273), .B2(new_n211), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n484), .B1(new_n511), .B2(new_n230), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT80), .B1(new_n271), .B2(new_n224), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT80), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n263), .A2(new_n514), .A3(G244), .A4(G1698), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT81), .A2(G116), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(KEYINPUT81), .A2(G116), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G33), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n263), .A2(G238), .A3(new_n264), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n513), .A2(new_n515), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n512), .B1(new_n522), .B2(new_n274), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n439), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT19), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n303), .B2(new_n225), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n263), .A2(new_n212), .A3(G68), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n212), .B1(new_n383), .B2(new_n525), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n229), .A2(new_n225), .A3(new_n325), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n291), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n306), .A2(new_n344), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n532), .B(new_n533), .C1(new_n466), .C2(new_n344), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n524), .B(new_n534), .C1(G169), .C2(new_n523), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n523), .A2(G190), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n308), .A2(new_n465), .A3(G87), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n532), .A2(new_n537), .A3(new_n533), .ZN(new_n538));
  INV_X1    g0338(.A(new_n286), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n536), .B(new_n538), .C1(new_n539), .C2(new_n523), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n510), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(G116), .B1(new_n267), .B2(G1), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n306), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g0344(.A1(KEYINPUT81), .A2(G116), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n516), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n544), .A2(new_n336), .B1(new_n306), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n546), .A2(G20), .B1(new_n211), .B2(new_n290), .ZN(new_n548));
  AOI21_X1  g0348(.A(G20), .B1(new_n267), .B2(G97), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n496), .B2(new_n497), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT20), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(G20), .B1(new_n517), .B2(new_n518), .ZN(new_n552));
  AND4_X1   g0352(.A1(KEYINPUT20), .A2(new_n550), .A3(new_n291), .A4(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n547), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n268), .A2(new_n270), .A3(G264), .A4(G1698), .ZN(new_n555));
  INV_X1    g0355(.A(G303), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(new_n263), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n327), .A2(new_n226), .A3(G1698), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n274), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n481), .A2(new_n484), .ZN(new_n560));
  OR2_X1    g0360(.A1(KEYINPUT5), .A2(G41), .ZN(new_n561));
  NAND2_X1  g0361(.A1(KEYINPUT5), .A2(G41), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(new_n562), .C1(new_n273), .C2(new_n211), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n511), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n560), .B1(new_n564), .B2(G270), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n554), .A2(new_n566), .A3(KEYINPUT21), .A4(G169), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n554), .A2(G179), .A3(new_n559), .A4(new_n565), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n554), .A2(G169), .A3(new_n566), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n268), .A2(new_n270), .A3(G257), .A4(G1698), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT83), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n263), .A2(KEYINPUT83), .A3(G257), .A4(G1698), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G294), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n263), .A2(G250), .A3(new_n264), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n274), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n564), .A2(G264), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n486), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n333), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT25), .B1(new_n461), .B2(G107), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT25), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n306), .A2(new_n586), .A3(new_n325), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n475), .B2(G107), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n268), .A2(new_n270), .A3(new_n212), .A4(G87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT22), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT22), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n263), .A2(new_n592), .A3(new_n212), .A4(G87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n302), .A2(new_n545), .A3(new_n516), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT23), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n212), .B2(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n325), .A2(KEYINPUT23), .A3(G20), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  XOR2_X1   g0401(.A(KEYINPUT82), .B(KEYINPUT24), .Z(new_n602));
  NAND3_X1  g0402(.A1(new_n594), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n291), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n591), .B2(new_n593), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n602), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n589), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n580), .A2(new_n274), .B1(G264), .B2(new_n564), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n439), .A3(new_n486), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n584), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT84), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n584), .A2(new_n607), .A3(new_n609), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT84), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n573), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT85), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n336), .B1(new_n605), .B2(new_n602), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n594), .A2(new_n601), .ZN(new_n618));
  INV_X1    g0418(.A(new_n602), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n581), .A2(G190), .A3(new_n582), .A4(new_n486), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n622), .A3(new_n589), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n399), .B1(new_n608), .B2(new_n486), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n616), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n585), .B(new_n587), .C1(new_n466), .C2(new_n325), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n620), .B2(new_n617), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n583), .A2(G200), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT85), .A4(new_n622), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n554), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n566), .A2(G200), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n631), .B(new_n632), .C1(new_n288), .C2(new_n566), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n542), .A2(new_n615), .A3(new_n630), .A4(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n450), .A2(new_n634), .ZN(G372));
  INV_X1    g0435(.A(KEYINPUT87), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT18), .B1(new_n438), .B2(new_n445), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n435), .A2(new_n447), .A3(new_n444), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n446), .A2(new_n448), .A3(KEYINPUT87), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n334), .A2(new_n347), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n359), .B1(new_n643), .B2(new_n349), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n400), .A2(new_n348), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n396), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT88), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n646), .A2(new_n647), .B1(new_n433), .B2(new_n437), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(new_n396), .A3(KEYINPUT88), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n642), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n319), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n450), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n569), .A2(new_n613), .A3(new_n572), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n630), .A2(new_n541), .A3(new_n510), .A4(new_n654), .ZN(new_n655));
  OAI22_X1  g0455(.A1(new_n502), .A2(G179), .B1(G169), .B2(new_n503), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n478), .B1(KEYINPUT86), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT86), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n508), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n657), .A2(new_n541), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n535), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n535), .A2(new_n540), .A3(new_n508), .A4(new_n509), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(KEYINPUT26), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n655), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n653), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n652), .A2(new_n324), .A3(new_n666), .ZN(G369));
  NAND2_X1  g0467(.A1(new_n612), .A2(new_n614), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(new_n630), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n217), .A2(G20), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(new_n276), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n276), .A2(new_n212), .A3(G13), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(new_n674), .A3(G213), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT89), .ZN(new_n676));
  XOR2_X1   g0476(.A(KEYINPUT90), .B(G343), .Z(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n669), .B1(new_n627), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n613), .B2(new_n680), .ZN(new_n682));
  INV_X1    g0482(.A(new_n573), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n633), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n680), .A2(new_n631), .ZN(new_n685));
  MUX2_X1   g0485(.A(new_n684), .B(new_n683), .S(new_n685), .Z(new_n686));
  INV_X1    g0486(.A(G330), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n683), .A2(new_n679), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n669), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n613), .B2(new_n679), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n690), .A2(new_n693), .ZN(G399));
  NOR2_X1   g0494(.A1(new_n218), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n529), .A2(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n209), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g0499(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n700));
  XNOR2_X1  g0500(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n657), .A2(new_n541), .A3(new_n660), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT26), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n662), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n542), .A2(new_n630), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n704), .B(new_n706), .C1(new_n707), .C2(new_n615), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n702), .B1(new_n708), .B2(new_n680), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n665), .A2(new_n680), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(KEYINPUT29), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n523), .A2(new_n503), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n566), .A2(new_n439), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(KEYINPUT30), .A3(new_n608), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n522), .A2(new_n274), .ZN(new_n717));
  INV_X1    g0517(.A(new_n512), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(G179), .B1(new_n559), .B2(new_n565), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n502), .A2(new_n583), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n608), .A2(G179), .A3(new_n559), .A4(new_n565), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n713), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n716), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n679), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT31), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n634), .B2(new_n679), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n712), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(KEYINPUT92), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(KEYINPUT92), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n701), .B1(new_n734), .B2(G1), .ZN(G364));
  NAND2_X1  g0535(.A1(new_n670), .A2(G45), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT93), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n276), .B1(new_n736), .B2(KEYINPUT93), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n695), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n211), .B1(G20), .B2(new_n333), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n218), .A2(new_n263), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT94), .Z(new_n748));
  INV_X1    g0548(.A(G45), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n210), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n748), .B(new_n750), .C1(new_n749), .C2(new_n258), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n218), .A2(new_n327), .ZN(new_n752));
  INV_X1    g0552(.A(G116), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n752), .A2(G355), .B1(new_n753), .B2(new_n218), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(G20), .A2(G179), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT95), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G190), .A3(new_n399), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n757), .A2(new_n288), .A3(new_n399), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G58), .A2(new_n759), .B1(new_n761), .B2(G77), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n757), .A2(new_n288), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n399), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n762), .B1(new_n203), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n212), .A2(G179), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n286), .A2(G190), .A3(new_n767), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT97), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT97), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G87), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n212), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G159), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT32), .Z(new_n776));
  NAND3_X1  g0576(.A1(new_n286), .A2(new_n288), .A3(new_n767), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n325), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n288), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n212), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n327), .B(new_n778), .C1(G97), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n773), .A2(new_n776), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(KEYINPUT96), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(KEYINPUT96), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n766), .B(new_n783), .C1(G50), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G326), .ZN(new_n791));
  INV_X1    g0591(.A(G294), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n788), .A2(new_n791), .B1(new_n792), .B2(new_n780), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT98), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n263), .B1(new_n774), .B2(G329), .ZN(new_n796));
  INV_X1    g0596(.A(G283), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n777), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(new_n764), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G311), .A2(new_n761), .B1(new_n759), .B2(G322), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n800), .B(new_n801), .C1(new_n556), .C2(new_n771), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n794), .B2(new_n793), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n790), .B1(new_n795), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n744), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n740), .B1(new_n746), .B2(new_n755), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n686), .B2(new_n743), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n686), .A2(new_n687), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n688), .A2(new_n740), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  NAND2_X1  g0611(.A1(new_n679), .A2(new_n347), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n364), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n361), .A2(KEYINPUT99), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n812), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(new_n361), .B2(KEYINPUT99), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT100), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT100), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n361), .A2(KEYINPUT99), .A3(new_n813), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT99), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n644), .B2(new_n348), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n818), .B(new_n819), .C1(new_n821), .C2(new_n815), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n710), .B(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n634), .A2(new_n679), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n687), .B1(new_n825), .B2(new_n727), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n740), .B1(new_n824), .B2(new_n826), .ZN(new_n829));
  INV_X1    g0629(.A(new_n823), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n741), .ZN(new_n831));
  INV_X1    g0631(.A(new_n740), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G143), .A2(new_n759), .B1(new_n761), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n296), .B2(new_n765), .C1(new_n788), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT34), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  INV_X1    g0637(.A(new_n774), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n263), .B1(new_n780), .B2(new_n202), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n777), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(G68), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n836), .B(new_n841), .C1(new_n201), .C2(new_n771), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n765), .A2(new_n797), .B1(new_n792), .B2(new_n758), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n760), .A2(new_n546), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n777), .A2(new_n229), .ZN(new_n845));
  INV_X1    g0645(.A(G311), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n327), .B1(new_n780), .B2(new_n225), .C1(new_n846), .C2(new_n838), .ZN(new_n847));
  NOR4_X1   g0647(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n848), .B1(new_n325), .B2(new_n771), .C1(new_n556), .C2(new_n788), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n805), .B1(new_n842), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n744), .A2(new_n741), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n832), .B(new_n850), .C1(new_n223), .C2(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n828), .A2(new_n829), .B1(new_n831), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G384));
  OAI211_X1 g0654(.A(G116), .B(new_n213), .C1(new_n456), .C2(KEYINPUT35), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(KEYINPUT35), .B2(new_n456), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT36), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n411), .A2(G77), .A3(new_n210), .A4(new_n413), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(G50), .B2(new_n203), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n276), .A2(G13), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n642), .A2(new_n676), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n379), .A2(new_n679), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n396), .A2(new_n400), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n379), .B(new_n679), .C1(new_n394), .C2(new_n395), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n823), .A2(new_n665), .A3(new_n680), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n361), .A2(new_n679), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n867), .A2(KEYINPUT101), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT101), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n866), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n425), .A2(new_n294), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n414), .A2(G20), .B1(G159), .B2(new_n297), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT16), .B1(new_n875), .B2(new_n424), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n431), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n676), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n433), .A2(new_n437), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n446), .A2(new_n448), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n444), .A2(new_n676), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n877), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n885), .B2(new_n432), .ZN(new_n886));
  INV_X1    g0686(.A(new_n432), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n426), .A2(new_n431), .B1(new_n444), .B2(new_n676), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n886), .B1(new_n889), .B2(new_n883), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n873), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n886), .ZN(new_n892));
  INV_X1    g0692(.A(new_n888), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(new_n883), .A3(new_n432), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(KEYINPUT38), .C1(new_n449), .C2(new_n879), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n862), .B1(new_n872), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT37), .B1(new_n887), .B2(new_n888), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n901), .A2(new_n894), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n446), .A2(new_n448), .A3(KEYINPUT87), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT87), .B1(new_n446), .B2(new_n448), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n880), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n438), .A2(new_n878), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n902), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n900), .B(new_n896), .C1(new_n908), .C2(KEYINPUT38), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT102), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n897), .A2(KEYINPUT39), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n396), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n680), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n899), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n653), .B1(new_n709), .B2(new_n711), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n324), .B1(new_n650), .B2(new_n651), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n918), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n653), .A2(new_n728), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT104), .Z(new_n925));
  AND3_X1   g0725(.A1(new_n728), .A2(new_n823), .A3(new_n866), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT40), .B1(new_n926), .B2(new_n897), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n896), .B1(new_n908), .B2(KEYINPUT38), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT103), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT103), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(new_n896), .C1(new_n908), .C2(KEYINPUT38), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n728), .A2(new_n866), .A3(KEYINPUT40), .A4(new_n823), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n927), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n687), .B1(new_n925), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n935), .B2(new_n925), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n923), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n276), .B2(new_n670), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n923), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n861), .B1(new_n939), .B2(new_n940), .ZN(G367));
  INV_X1    g0741(.A(new_n748), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(new_n254), .ZN(new_n943));
  INV_X1    g0743(.A(new_n218), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n745), .B1(new_n944), .B2(new_n344), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n740), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(G159), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n765), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n777), .A2(new_n223), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n781), .A2(G68), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n263), .C1(new_n834), .C2(new_n838), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n201), .A2(new_n760), .B1(new_n758), .B2(new_n296), .ZN(new_n952));
  NOR4_X1   g0752(.A1(new_n948), .A2(new_n949), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(G143), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n953), .B1(new_n202), .B2(new_n771), .C1(new_n954), .C2(new_n788), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n777), .A2(new_n225), .ZN(new_n956));
  INV_X1    g0756(.A(G317), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n327), .B1(new_n780), .B2(new_n325), .C1(new_n957), .C2(new_n838), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n956), .B(new_n958), .C1(G303), .C2(new_n759), .ZN(new_n959));
  AOI22_X1  g0759(.A1(G294), .A2(new_n764), .B1(new_n761), .B2(G283), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(new_n846), .C2(new_n788), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n546), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n772), .A2(G116), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n962), .B1(KEYINPUT46), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n955), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT47), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n805), .B1(new_n965), .B2(new_n966), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n946), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n743), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n541), .B1(new_n538), .B2(new_n680), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n535), .A2(new_n538), .A3(new_n680), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n969), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT110), .Z(new_n975));
  NAND2_X1  g0775(.A1(new_n508), .A2(new_n509), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n657), .A2(new_n660), .A3(new_n679), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n510), .B1(new_n478), .B2(new_n680), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT105), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n976), .B1(new_n980), .B2(new_n668), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n680), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n692), .A2(new_n979), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT42), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n982), .A2(new_n984), .B1(KEYINPUT43), .B2(new_n973), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n987), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n689), .A2(new_n980), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT106), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n992), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n990), .A2(KEYINPUT106), .A3(new_n992), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n693), .A2(new_n979), .ZN(new_n998));
  XOR2_X1   g0798(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n693), .A2(new_n979), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(KEYINPUT108), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT108), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n693), .A2(new_n1003), .A3(new_n979), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(KEYINPUT44), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT44), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n690), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1007), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1009), .A2(new_n1000), .A3(new_n689), .A4(new_n1005), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n688), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1012), .A2(KEYINPUT109), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n682), .A2(new_n691), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n692), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n1012), .B2(KEYINPUT109), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1013), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n734), .B1(new_n1011), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n695), .B(KEYINPUT41), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n739), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n975), .B1(new_n997), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(G387));
  OR2_X1    g0826(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n734), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1019), .A2(new_n732), .A3(new_n733), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n695), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n682), .A2(new_n970), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n697), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n752), .A2(new_n1032), .B1(new_n325), .B2(new_n218), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n749), .B1(new_n203), .B2(new_n223), .C1(new_n1032), .C2(KEYINPUT111), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(KEYINPUT111), .ZN(new_n1035));
  OR3_X1    g0835(.A1(new_n301), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1036));
  OAI21_X1  g0836(.A(KEYINPUT50), .B1(new_n301), .B2(G50), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n748), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n250), .A2(new_n749), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1033), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n745), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n740), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n789), .A2(G159), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n772), .A2(G77), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n760), .A2(new_n203), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n263), .B1(new_n838), .B2(new_n296), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n780), .A2(new_n344), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1046), .A2(new_n956), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n427), .A2(new_n764), .B1(new_n759), .B2(G50), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1044), .A2(new_n1045), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n263), .B1(new_n774), .B2(G326), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n789), .A2(G322), .B1(G311), .B2(new_n764), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n556), .A2(new_n760), .B1(new_n758), .B2(new_n957), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT112), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT48), .Z(new_n1057));
  OAI22_X1  g0857(.A1(new_n771), .A2(new_n792), .B1(new_n797), .B2(new_n780), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1052), .B1(new_n546), .B2(new_n777), .C1(new_n1059), .C2(KEYINPUT49), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1059), .A2(KEYINPUT49), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1051), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1031), .B(new_n1043), .C1(new_n1062), .C2(new_n744), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n1027), .B2(new_n739), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1030), .A2(new_n1064), .ZN(G393));
  NAND3_X1  g0865(.A1(new_n1008), .A2(KEYINPUT113), .A3(new_n1010), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT113), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n690), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(new_n1028), .A3(new_n1068), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n695), .C1(new_n1028), .C2(new_n1011), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n263), .B1(new_n780), .B2(new_n223), .C1(new_n954), .C2(new_n838), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n845), .B(new_n1071), .C1(G50), .C2(new_n764), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n301), .B2(new_n760), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n788), .A2(new_n296), .B1(new_n947), .B2(new_n758), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT51), .Z(new_n1075));
  AOI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(new_n367), .C2(new_n772), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n788), .A2(new_n957), .B1(new_n846), .B2(new_n758), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT52), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n772), .A2(G283), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n765), .A2(new_n556), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n760), .A2(new_n792), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n263), .B1(new_n774), .B2(G322), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n546), .B2(new_n780), .ZN(new_n1084));
  NOR4_X1   g0884(.A1(new_n1081), .A2(new_n778), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1079), .A2(new_n1080), .A3(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n744), .B1(new_n1076), .B2(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n748), .A2(new_n261), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n745), .B1(new_n944), .B2(new_n225), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1089), .B(new_n740), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n980), .B2(new_n743), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n739), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1070), .A2(new_n1095), .ZN(G390));
  INV_X1    g0896(.A(new_n866), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n729), .A2(new_n830), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n909), .A2(new_n911), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT102), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n909), .A2(new_n911), .A3(new_n910), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1100), .A2(new_n1101), .B1(new_n916), .B2(new_n872), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n708), .A2(new_n680), .A3(new_n823), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n869), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n917), .B1(new_n1104), .B2(new_n866), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n932), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1098), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n872), .A2(new_n916), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n912), .B2(new_n913), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1098), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n932), .A2(new_n1105), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n914), .A2(new_n742), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n832), .B1(new_n301), .B2(new_n851), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n773), .A2(new_n327), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT117), .Z(new_n1117));
  OAI22_X1  g0917(.A1(new_n777), .A2(new_n203), .B1(new_n792), .B2(new_n838), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT118), .Z(new_n1119));
  AOI22_X1  g0919(.A1(new_n764), .A2(G107), .B1(G77), .B2(new_n781), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n225), .B2(new_n760), .C1(new_n753), .C2(new_n758), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1119), .B(new_n1121), .C1(G283), .C2(new_n789), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n765), .A2(new_n834), .B1(new_n837), .B2(new_n758), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n780), .A2(new_n947), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n327), .B(new_n1124), .C1(G125), .C2(new_n774), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT54), .B(G143), .Z(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1125), .B1(new_n201), .B2(new_n777), .C1(new_n760), .C2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1123), .B(new_n1128), .C1(G128), .C2(new_n789), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n771), .A2(new_n296), .ZN(new_n1130));
  XOR2_X1   g0930(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1131));
  XNOR2_X1  g0931(.A(new_n1130), .B(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1117), .A2(new_n1122), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1115), .B1(new_n1133), .B2(new_n805), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1113), .A2(new_n1023), .B1(new_n1114), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n653), .A2(G330), .A3(new_n728), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n652), .A2(new_n324), .A3(new_n919), .A4(new_n1137), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n870), .A2(new_n871), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n728), .A2(G330), .A3(new_n823), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1140), .A2(new_n1097), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1141), .B2(new_n1098), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n866), .B1(KEYINPUT114), .B2(new_n823), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1104), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1138), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1107), .A2(new_n1112), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT115), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n695), .B(new_n1149), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1148), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1113), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(KEYINPUT115), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1136), .B1(new_n1152), .B2(new_n1155), .ZN(G378));
  INV_X1    g0956(.A(KEYINPUT121), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n931), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n906), .B1(new_n641), .B2(new_n880), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n873), .B1(new_n1159), .B2(new_n902), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n930), .B1(new_n1160), .B2(new_n896), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n934), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n927), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1163), .A3(G330), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT120), .B1(new_n319), .B2(new_n324), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n310), .A2(new_n878), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n319), .A2(KEYINPUT120), .A3(new_n324), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT120), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1170), .B(new_n323), .C1(new_n317), .C2(new_n318), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n310), .B(new_n878), .C1(new_n1165), .C2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1169), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1164), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1176), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n935), .A2(G330), .A3(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1177), .A2(new_n918), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n918), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT57), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1110), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1138), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1157), .B1(new_n1182), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1138), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1149), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1100), .A2(new_n917), .A3(new_n1101), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1191), .B(new_n862), .C1(new_n898), .C2(new_n872), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1178), .B1(new_n935), .B2(G330), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n933), .B1(new_n929), .B2(new_n931), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1194), .A2(new_n1176), .A3(new_n927), .A4(new_n687), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1192), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1177), .A2(new_n918), .A3(new_n1179), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1190), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT57), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1200), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1202), .A2(KEYINPUT121), .A3(new_n1190), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1188), .A2(new_n1201), .A3(new_n695), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1176), .A2(new_n741), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n263), .A2(G41), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n838), .B2(new_n797), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n777), .A2(new_n202), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(G68), .C2(new_n781), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n760), .A2(new_n344), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G97), .A2(new_n764), .B1(new_n759), .B2(G107), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1212), .B(new_n1045), .C1(new_n753), .C2(new_n788), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT58), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1215), .B(new_n1216), .C1(new_n1206), .C2(new_n1217), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G132), .A2(new_n764), .B1(new_n761), .B2(G137), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n759), .A2(G128), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n771), .C2(new_n1127), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n789), .A2(G125), .B1(G150), .B2(new_n781), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(KEYINPUT119), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(KEYINPUT119), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1221), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G33), .B(G41), .C1(new_n774), .C2(G124), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n947), .B2(new_n777), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1228), .B2(KEYINPUT59), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1218), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(new_n805), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n832), .B(new_n1235), .C1(new_n201), .C2(new_n851), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1198), .A2(new_n739), .B1(new_n1205), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1204), .A2(new_n1237), .ZN(G375));
  NAND2_X1  g1038(.A1(new_n1097), .A2(new_n741), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n744), .A2(G68), .A3(new_n741), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n760), .A2(new_n296), .B1(new_n201), .B2(new_n780), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT122), .Z(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n837), .B2(new_n788), .ZN(new_n1243));
  INV_X1    g1043(.A(G128), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n263), .B1(new_n838), .B2(new_n1244), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1245), .B(new_n1208), .C1(new_n764), .C2(new_n1126), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1246), .B1(new_n834), .B2(new_n758), .C1(new_n947), .C2(new_n771), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n788), .A2(new_n792), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n772), .A2(G97), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n519), .A2(new_n764), .B1(new_n759), .B2(G283), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n761), .A2(G107), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n327), .B1(new_n838), .B2(new_n556), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n949), .A2(new_n1252), .A3(new_n1048), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .A4(new_n1253), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n1243), .A2(new_n1247), .B1(new_n1248), .B2(new_n1254), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n832), .B(new_n1240), .C1(new_n1255), .C2(new_n744), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1186), .A2(new_n739), .B1(new_n1239), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1153), .A2(new_n1021), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(G381));
  INV_X1    g1060(.A(new_n1237), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1202), .A2(KEYINPUT121), .A3(new_n1190), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT121), .B1(new_n1202), .B2(new_n1190), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n696), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1261), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G378), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1030), .A2(new_n810), .A3(new_n1064), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1266), .A2(new_n1025), .A3(new_n1267), .A4(new_n1269), .ZN(G407));
  NAND2_X1  g1070(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G407), .B(G213), .C1(new_n677), .C2(new_n1271), .ZN(G409));
  NAND2_X1  g1072(.A1(G393), .A2(G396), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1268), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n1070), .A3(new_n1095), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(G390), .A2(new_n1268), .A3(new_n1273), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1025), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(new_n1275), .A3(new_n1025), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1281), .A2(KEYINPUT123), .A3(KEYINPUT60), .A4(new_n1138), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1138), .A2(new_n1142), .A3(new_n1147), .A4(KEYINPUT60), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT123), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n696), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1282), .A2(new_n1285), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1289), .A2(G384), .A3(new_n1257), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G384), .B1(new_n1289), .B2(new_n1257), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT124), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT124), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n678), .A2(G213), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(G2897), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1295), .A2(new_n1299), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1294), .B(new_n1298), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1267), .B1(new_n1204), .B2(new_n1237), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1190), .A2(new_n1198), .A3(new_n1021), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1237), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1296), .B1(G378), .B2(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1293), .B(new_n1302), .C1(new_n1303), .C2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1292), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(new_n1303), .A2(new_n1309), .A3(new_n1306), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1307), .B(new_n1308), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1306), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1313), .B(new_n1292), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1314), .A2(KEYINPUT62), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1280), .B1(new_n1312), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT125), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1306), .B1(G375), .B2(G378), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1302), .A2(new_n1293), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1308), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT63), .B1(new_n1318), .B2(new_n1292), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1280), .B1(new_n1310), .B2(KEYINPUT63), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1317), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1307), .B(new_n1308), .C1(new_n1310), .C2(KEYINPUT63), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1279), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1326), .A2(new_n1277), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1327), .B1(new_n1314), .B2(new_n1328), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1325), .A2(new_n1329), .A3(KEYINPUT125), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1316), .B1(new_n1324), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT126), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1333), .B(new_n1316), .C1(new_n1324), .C2(new_n1330), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1332), .A2(new_n1334), .ZN(G405));
  INV_X1    g1135(.A(new_n1303), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1271), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1309), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1336), .A2(new_n1271), .A3(new_n1292), .ZN(new_n1339));
  AOI22_X1  g1139(.A1(new_n1338), .A2(new_n1339), .B1(KEYINPUT127), .B2(new_n1280), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1280), .A2(KEYINPUT127), .ZN(new_n1341));
  XOR2_X1   g1141(.A(new_n1340), .B(new_n1341), .Z(G402));
endmodule


