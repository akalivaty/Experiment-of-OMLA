

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596;

  XOR2_X1 U325 ( .A(KEYINPUT111), .B(n367), .Z(n293) );
  NOR2_X1 U326 ( .A1(n537), .A2(n526), .ZN(n472) );
  NOR2_X1 U327 ( .A1(n562), .A2(n371), .ZN(n372) );
  NOR2_X1 U328 ( .A1(n535), .A2(n526), .ZN(n400) );
  XOR2_X1 U329 ( .A(G176GAT), .B(G64GAT), .Z(n384) );
  INV_X1 U330 ( .A(KEYINPUT97), .ZN(n395) );
  XNOR2_X1 U331 ( .A(n566), .B(KEYINPUT55), .ZN(n567) );
  NOR2_X1 U332 ( .A1(n373), .A2(n482), .ZN(n483) );
  XNOR2_X1 U333 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U334 ( .A(n568), .B(n567), .ZN(n572) );
  XOR2_X1 U335 ( .A(n348), .B(n347), .Z(n353) );
  XNOR2_X1 U336 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U337 ( .A(KEYINPUT124), .B(n463), .Z(n595) );
  XOR2_X1 U338 ( .A(n353), .B(n352), .Z(n569) );
  XOR2_X1 U339 ( .A(n441), .B(n440), .Z(n573) );
  XNOR2_X1 U340 ( .A(n464), .B(G218GAT), .ZN(n465) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n485) );
  XNOR2_X1 U342 ( .A(n466), .B(n465), .ZN(G1355GAT) );
  XNOR2_X1 U343 ( .A(n486), .B(n485), .ZN(G1330GAT) );
  INV_X1 U344 ( .A(KEYINPUT74), .ZN(n318) );
  XOR2_X1 U345 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n295) );
  XNOR2_X1 U346 ( .A(G134GAT), .B(KEYINPUT72), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n309) );
  XNOR2_X1 U348 ( .A(G36GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n296), .B(G218GAT), .ZN(n394) );
  XOR2_X1 U350 ( .A(G50GAT), .B(G162GAT), .Z(n449) );
  XNOR2_X1 U351 ( .A(n394), .B(n449), .ZN(n297) );
  AND2_X1 U352 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  NAND2_X1 U353 ( .A1(n297), .A2(n298), .ZN(n302) );
  INV_X1 U354 ( .A(n297), .ZN(n300) );
  INV_X1 U355 ( .A(n298), .ZN(n299) );
  NAND2_X1 U356 ( .A1(n300), .A2(n299), .ZN(n301) );
  NAND2_X1 U357 ( .A1(n302), .A2(n301), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n303), .B(KEYINPUT9), .ZN(n307) );
  XOR2_X1 U359 ( .A(G92GAT), .B(G85GAT), .Z(n305) );
  XNOR2_X1 U360 ( .A(G99GAT), .B(G106GAT), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n305), .B(n304), .ZN(n354) );
  XOR2_X1 U362 ( .A(n354), .B(KEYINPUT10), .Z(n306) );
  XNOR2_X1 U363 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n317) );
  INV_X1 U365 ( .A(KEYINPUT7), .ZN(n310) );
  NAND2_X1 U366 ( .A1(KEYINPUT69), .A2(n310), .ZN(n313) );
  INV_X1 U367 ( .A(KEYINPUT69), .ZN(n311) );
  NAND2_X1 U368 ( .A1(n311), .A2(KEYINPUT7), .ZN(n312) );
  NAND2_X1 U369 ( .A1(n313), .A2(n312), .ZN(n315) );
  XNOR2_X1 U370 ( .A(G43GAT), .B(G29GAT), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U372 ( .A(KEYINPUT8), .B(n316), .Z(n339) );
  XOR2_X1 U373 ( .A(n317), .B(n339), .Z(n562) );
  XNOR2_X1 U374 ( .A(n318), .B(n562), .ZN(n487) );
  XNOR2_X1 U375 ( .A(n487), .B(KEYINPUT36), .ZN(n373) );
  XOR2_X1 U376 ( .A(KEYINPUT76), .B(KEYINPUT14), .Z(n320) );
  XNOR2_X1 U377 ( .A(KEYINPUT78), .B(KEYINPUT15), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U379 ( .A(KEYINPUT79), .B(KEYINPUT77), .Z(n322) );
  XNOR2_X1 U380 ( .A(G64GAT), .B(KEYINPUT75), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n337) );
  XOR2_X1 U383 ( .A(G71GAT), .B(G127GAT), .Z(n326) );
  XNOR2_X1 U384 ( .A(G22GAT), .B(G183GAT), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U386 ( .A(KEYINPUT12), .B(G155GAT), .Z(n328) );
  XNOR2_X1 U387 ( .A(G211GAT), .B(G78GAT), .ZN(n327) );
  XNOR2_X1 U388 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U389 ( .A(n330), .B(n329), .Z(n335) );
  XOR2_X1 U390 ( .A(G15GAT), .B(G1GAT), .Z(n338) );
  XOR2_X1 U391 ( .A(G57GAT), .B(KEYINPUT13), .Z(n356) );
  XOR2_X1 U392 ( .A(n356), .B(G8GAT), .Z(n332) );
  NAND2_X1 U393 ( .A1(G231GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n338), .B(n333), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U397 ( .A(n337), .B(n336), .Z(n480) );
  INV_X1 U398 ( .A(n480), .ZN(n594) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n344) );
  XOR2_X1 U400 ( .A(G197GAT), .B(G113GAT), .Z(n341) );
  XNOR2_X1 U401 ( .A(G50GAT), .B(G36GAT), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U403 ( .A(G169GAT), .B(G8GAT), .Z(n385) );
  XOR2_X1 U404 ( .A(n342), .B(n385), .Z(n343) );
  XNOR2_X1 U405 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U406 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n346) );
  NAND2_X1 U407 ( .A1(G229GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U409 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n350) );
  XNOR2_X1 U410 ( .A(KEYINPUT30), .B(KEYINPUT66), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U412 ( .A(G141GAT), .B(G22GAT), .Z(n455) );
  XNOR2_X1 U413 ( .A(n351), .B(n455), .ZN(n352) );
  XNOR2_X1 U414 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n366) );
  XOR2_X1 U415 ( .A(n354), .B(n384), .Z(n358) );
  XNOR2_X1 U416 ( .A(G78GAT), .B(G204GAT), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n355), .B(G148GAT), .ZN(n451) );
  XNOR2_X1 U418 ( .A(n451), .B(n356), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n365) );
  XOR2_X1 U420 ( .A(G120GAT), .B(G71GAT), .Z(n429) );
  XOR2_X1 U421 ( .A(KEYINPUT71), .B(KEYINPUT31), .Z(n360) );
  XNOR2_X1 U422 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U424 ( .A(n429), .B(n361), .Z(n363) );
  NAND2_X1 U425 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n591) );
  XOR2_X1 U428 ( .A(n366), .B(n591), .Z(n571) );
  NAND2_X1 U429 ( .A1(n569), .A2(n571), .ZN(n368) );
  XOR2_X1 U430 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n293), .ZN(n369) );
  NOR2_X1 U432 ( .A1(n594), .A2(n369), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n370), .B(KEYINPUT113), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(KEYINPUT47), .ZN(n378) );
  NOR2_X1 U435 ( .A1(n373), .A2(n480), .ZN(n374) );
  XOR2_X1 U436 ( .A(KEYINPUT45), .B(n374), .Z(n375) );
  NOR2_X1 U437 ( .A1(n591), .A2(n375), .ZN(n376) );
  INV_X1 U438 ( .A(n569), .ZN(n588) );
  NAND2_X1 U439 ( .A1(n376), .A2(n588), .ZN(n377) );
  NAND2_X1 U440 ( .A1(n378), .A2(n377), .ZN(n380) );
  INV_X1 U441 ( .A(KEYINPUT48), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n380), .B(n379), .ZN(n535) );
  XOR2_X1 U443 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n382) );
  XNOR2_X1 U444 ( .A(KEYINPUT84), .B(G183GAT), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U446 ( .A(KEYINPUT17), .B(n383), .Z(n441) );
  XOR2_X1 U447 ( .A(G92GAT), .B(n384), .Z(n387) );
  XNOR2_X1 U448 ( .A(n385), .B(G204GAT), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U450 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n389) );
  XNOR2_X1 U451 ( .A(KEYINPUT86), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U453 ( .A(G197GAT), .B(n390), .Z(n442) );
  XNOR2_X1 U454 ( .A(n391), .B(n442), .ZN(n393) );
  AND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n394), .B(KEYINPUT96), .ZN(n396) );
  XOR2_X1 U458 ( .A(n441), .B(n399), .Z(n505) );
  INV_X1 U459 ( .A(n505), .ZN(n526) );
  XNOR2_X1 U460 ( .A(n400), .B(KEYINPUT54), .ZN(n425) );
  XOR2_X1 U461 ( .A(KEYINPUT92), .B(KEYINPUT95), .Z(n402) );
  XNOR2_X1 U462 ( .A(G1GAT), .B(G57GAT), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n412) );
  XOR2_X1 U464 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n410) );
  XNOR2_X1 U465 ( .A(G127GAT), .B(KEYINPUT80), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n403), .B(KEYINPUT0), .ZN(n404) );
  XOR2_X1 U467 ( .A(n404), .B(KEYINPUT81), .Z(n406) );
  XNOR2_X1 U468 ( .A(G113GAT), .B(G134GAT), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n437) );
  XOR2_X1 U470 ( .A(G155GAT), .B(KEYINPUT3), .Z(n408) );
  XNOR2_X1 U471 ( .A(KEYINPUT88), .B(KEYINPUT2), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n408), .B(n407), .ZN(n450) );
  XNOR2_X1 U473 ( .A(n437), .B(n450), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n424) );
  NAND2_X1 U476 ( .A1(G225GAT), .A2(G233GAT), .ZN(n418) );
  XOR2_X1 U477 ( .A(G148GAT), .B(G120GAT), .Z(n414) );
  XNOR2_X1 U478 ( .A(G29GAT), .B(G141GAT), .ZN(n413) );
  XNOR2_X1 U479 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U480 ( .A(G162GAT), .B(G85GAT), .Z(n415) );
  XNOR2_X1 U481 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U483 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n420) );
  XNOR2_X1 U484 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n419) );
  XNOR2_X1 U485 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U487 ( .A(n424), .B(n423), .Z(n523) );
  NAND2_X1 U488 ( .A1(n425), .A2(n523), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n426), .B(KEYINPUT65), .ZN(n565) );
  XOR2_X1 U490 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n428) );
  XNOR2_X1 U491 ( .A(G99GAT), .B(G190GAT), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U493 ( .A(n430), .B(n429), .Z(n432) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(G15GAT), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U496 ( .A(KEYINPUT83), .B(G176GAT), .Z(n434) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U499 ( .A(n436), .B(n435), .Z(n439) );
  XNOR2_X1 U500 ( .A(G169GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U502 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n444) );
  XNOR2_X1 U503 ( .A(KEYINPUT22), .B(KEYINPUT91), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U505 ( .A(KEYINPUT85), .B(KEYINPUT90), .Z(n446) );
  XNOR2_X1 U506 ( .A(G218GAT), .B(G106GAT), .ZN(n445) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n459) );
  XOR2_X1 U509 ( .A(n450), .B(n449), .Z(n457) );
  XOR2_X1 U510 ( .A(n451), .B(KEYINPUT24), .Z(n453) );
  NAND2_X1 U511 ( .A1(G228GAT), .A2(G233GAT), .ZN(n452) );
  XNOR2_X1 U512 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n442), .B(n460), .ZN(n564) );
  NOR2_X1 U517 ( .A1(n573), .A2(n564), .ZN(n462) );
  XNOR2_X1 U518 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n461) );
  XOR2_X1 U519 ( .A(n462), .B(n461), .Z(n552) );
  INV_X1 U520 ( .A(n552), .ZN(n470) );
  NAND2_X1 U521 ( .A1(n565), .A2(n470), .ZN(n463) );
  INV_X1 U522 ( .A(n595), .ZN(n587) );
  NOR2_X1 U523 ( .A1(n373), .A2(n587), .ZN(n466) );
  XNOR2_X1 U524 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n464) );
  INV_X1 U525 ( .A(n523), .ZN(n502) );
  XNOR2_X1 U526 ( .A(KEYINPUT27), .B(n505), .ZN(n471) );
  NAND2_X1 U527 ( .A1(n502), .A2(n471), .ZN(n534) );
  XOR2_X1 U528 ( .A(KEYINPUT28), .B(n564), .Z(n517) );
  NOR2_X1 U529 ( .A1(n534), .A2(n517), .ZN(n467) );
  XOR2_X1 U530 ( .A(KEYINPUT98), .B(n467), .Z(n468) );
  NOR2_X1 U531 ( .A1(n573), .A2(n468), .ZN(n469) );
  XNOR2_X1 U532 ( .A(n469), .B(KEYINPUT99), .ZN(n479) );
  NAND2_X1 U533 ( .A1(n471), .A2(n470), .ZN(n476) );
  INV_X1 U534 ( .A(n573), .ZN(n537) );
  XNOR2_X1 U535 ( .A(n472), .B(KEYINPUT101), .ZN(n473) );
  NAND2_X1 U536 ( .A1(n473), .A2(n564), .ZN(n474) );
  XOR2_X1 U537 ( .A(KEYINPUT25), .B(n474), .Z(n475) );
  NAND2_X1 U538 ( .A1(n476), .A2(n475), .ZN(n477) );
  NAND2_X1 U539 ( .A1(n477), .A2(n523), .ZN(n478) );
  NAND2_X1 U540 ( .A1(n479), .A2(n478), .ZN(n490) );
  NAND2_X1 U541 ( .A1(n490), .A2(n480), .ZN(n481) );
  XOR2_X1 U542 ( .A(KEYINPUT105), .B(n481), .Z(n482) );
  XOR2_X1 U543 ( .A(KEYINPUT37), .B(n483), .Z(n522) );
  NOR2_X1 U544 ( .A1(n588), .A2(n591), .ZN(n491) );
  NAND2_X1 U545 ( .A1(n522), .A2(n491), .ZN(n484) );
  XOR2_X1 U546 ( .A(KEYINPUT38), .B(n484), .Z(n508) );
  NAND2_X1 U547 ( .A1(n508), .A2(n573), .ZN(n486) );
  XOR2_X1 U548 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n494) );
  NAND2_X1 U549 ( .A1(n594), .A2(n487), .ZN(n488) );
  XOR2_X1 U550 ( .A(KEYINPUT16), .B(n488), .Z(n489) );
  AND2_X1 U551 ( .A1(n490), .A2(n489), .ZN(n512) );
  NAND2_X1 U552 ( .A1(n491), .A2(n512), .ZN(n492) );
  XOR2_X1 U553 ( .A(KEYINPUT102), .B(n492), .Z(n500) );
  NAND2_X1 U554 ( .A1(n502), .A2(n500), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G1GAT), .B(n495), .ZN(G1324GAT) );
  NAND2_X1 U557 ( .A1(n500), .A2(n505), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT35), .B(KEYINPUT104), .Z(n498) );
  NAND2_X1 U560 ( .A1(n573), .A2(n500), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G15GAT), .B(n499), .ZN(G1326GAT) );
  NAND2_X1 U563 ( .A1(n500), .A2(n517), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n501), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  NAND2_X1 U566 ( .A1(n502), .A2(n508), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  XNOR2_X1 U568 ( .A(G36GAT), .B(KEYINPUT106), .ZN(n507) );
  NAND2_X1 U569 ( .A1(n505), .A2(n508), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1329GAT) );
  XOR2_X1 U571 ( .A(G50GAT), .B(KEYINPUT107), .Z(n510) );
  NAND2_X1 U572 ( .A1(n508), .A2(n517), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1331GAT) );
  INV_X1 U574 ( .A(n571), .ZN(n511) );
  NOR2_X1 U575 ( .A1(n569), .A2(n511), .ZN(n521) );
  NAND2_X1 U576 ( .A1(n521), .A2(n512), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n523), .A2(n518), .ZN(n513) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n513), .Z(n514) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n526), .A2(n518), .ZN(n515) );
  XOR2_X1 U581 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U582 ( .A1(n537), .A2(n518), .ZN(n516) );
  XOR2_X1 U583 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  INV_X1 U584 ( .A(n517), .ZN(n539) );
  NOR2_X1 U585 ( .A1(n539), .A2(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n530) );
  NOR2_X1 U589 ( .A1(n523), .A2(n530), .ZN(n524) );
  XOR2_X1 U590 ( .A(G85GAT), .B(n524), .Z(n525) );
  XNOR2_X1 U591 ( .A(KEYINPUT108), .B(n525), .ZN(G1336GAT) );
  NOR2_X1 U592 ( .A1(n526), .A2(n530), .ZN(n527) );
  XOR2_X1 U593 ( .A(G92GAT), .B(n527), .Z(G1337GAT) );
  NOR2_X1 U594 ( .A1(n537), .A2(n530), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(G1338GAT) );
  NOR2_X1 U597 ( .A1(n539), .A2(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U600 ( .A(G106GAT), .B(n533), .Z(G1339GAT) );
  NOR2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U602 ( .A(KEYINPUT114), .B(n536), .Z(n553) );
  NOR2_X1 U603 ( .A1(n537), .A2(n553), .ZN(n538) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(KEYINPUT115), .B(n540), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n569), .A2(n548), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n541), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U609 ( .A1(n548), .A2(n571), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n546) );
  NAND2_X1 U613 ( .A1(n548), .A2(n594), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n550) );
  INV_X1 U617 ( .A(n487), .ZN(n580) );
  NAND2_X1 U618 ( .A1(n548), .A2(n580), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U620 ( .A(G134GAT), .B(n551), .ZN(G1343GAT) );
  NOR2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n561) );
  NAND2_X1 U622 ( .A1(n561), .A2(n569), .ZN(n554) );
  XNOR2_X1 U623 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n556) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n555) );
  XNOR2_X1 U626 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U627 ( .A(KEYINPUT52), .B(n557), .Z(n559) );
  NAND2_X1 U628 ( .A1(n561), .A2(n571), .ZN(n558) );
  XNOR2_X1 U629 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n561), .A2(n594), .ZN(n560) );
  XNOR2_X1 U631 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U633 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n565), .A2(n564), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n566) );
  AND2_X1 U636 ( .A1(n572), .A2(n573), .ZN(n581) );
  NAND2_X1 U637 ( .A1(n569), .A2(n581), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n570), .B(G169GAT), .ZN(G1348GAT) );
  AND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n576) );
  XOR2_X1 U641 ( .A(G176GAT), .B(KEYINPUT57), .Z(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n578) );
  XOR2_X1 U643 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1349GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n594), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n579), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT58), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n583), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n585) );
  XNOR2_X1 U651 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n584) );
  XNOR2_X1 U652 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U653 ( .A(KEYINPUT60), .B(n586), .ZN(n590) );
  NOR2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1352GAT) );
  XOR2_X1 U656 ( .A(G204GAT), .B(KEYINPUT61), .Z(n593) );
  NAND2_X1 U657 ( .A1(n595), .A2(n591), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(G1353GAT) );
  NAND2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(n596), .B(G211GAT), .ZN(G1354GAT) );
endmodule

