

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(n667), .ZN(n639) );
  NOR2_X1 U555 ( .A1(n706), .A2(n693), .ZN(n521) );
  OR2_X1 U556 ( .A1(n708), .A2(n707), .ZN(n522) );
  AND2_X1 U557 ( .A1(n741), .A2(n739), .ZN(n523) );
  AND2_X1 U558 ( .A1(n748), .A2(n523), .ZN(n524) );
  INV_X1 U559 ( .A(n675), .ZN(n656) );
  OR2_X1 U560 ( .A1(n678), .A2(n657), .ZN(n658) );
  NAND2_X1 U561 ( .A1(n605), .A2(n710), .ZN(n667) );
  NAND2_X1 U562 ( .A1(G8), .A2(n667), .ZN(n706) );
  INV_X1 U563 ( .A(KEYINPUT87), .ZN(n603) );
  NOR2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XNOR2_X1 U565 ( .A(n604), .B(n603), .ZN(n709) );
  AND2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n877) );
  XNOR2_X1 U567 ( .A(n530), .B(KEYINPUT66), .ZN(n773) );
  INV_X1 U568 ( .A(G2105), .ZN(n531) );
  AND2_X1 U569 ( .A1(n531), .A2(G2104), .ZN(n883) );
  NAND2_X1 U570 ( .A1(G101), .A2(n883), .ZN(n525) );
  XOR2_X1 U571 ( .A(KEYINPUT23), .B(n525), .Z(n528) );
  NAND2_X1 U572 ( .A1(G113), .A2(n877), .ZN(n526) );
  XOR2_X1 U573 ( .A(KEYINPUT65), .B(n526), .Z(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n535) );
  XOR2_X1 U575 ( .A(KEYINPUT17), .B(n529), .Z(n530) );
  NAND2_X1 U576 ( .A1(G137), .A2(n773), .ZN(n533) );
  NOR2_X1 U577 ( .A1(G2104), .A2(n531), .ZN(n878) );
  NAND2_X1 U578 ( .A1(G125), .A2(n878), .ZN(n532) );
  NAND2_X1 U579 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X2 U580 ( .A1(n535), .A2(n534), .ZN(G160) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n581) );
  NOR2_X1 U582 ( .A1(G651), .A2(n581), .ZN(n784) );
  NAND2_X1 U583 ( .A1(G51), .A2(n784), .ZN(n539) );
  INV_X1 U584 ( .A(G651), .ZN(n541) );
  NOR2_X1 U585 ( .A1(G543), .A2(n541), .ZN(n537) );
  XNOR2_X1 U586 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n536) );
  XNOR2_X1 U587 ( .A(n537), .B(n536), .ZN(n785) );
  NAND2_X1 U588 ( .A1(G63), .A2(n785), .ZN(n538) );
  NAND2_X1 U589 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U590 ( .A(KEYINPUT6), .B(n540), .Z(n550) );
  NOR2_X1 U591 ( .A1(n581), .A2(n541), .ZN(n780) );
  NAND2_X1 U592 ( .A1(n780), .A2(G76), .ZN(n542) );
  XNOR2_X1 U593 ( .A(KEYINPUT73), .B(n542), .ZN(n546) );
  NOR2_X1 U594 ( .A1(G543), .A2(G651), .ZN(n543) );
  XNOR2_X1 U595 ( .A(n543), .B(KEYINPUT64), .ZN(n781) );
  NAND2_X1 U596 ( .A1(G89), .A2(n781), .ZN(n544) );
  XOR2_X1 U597 ( .A(n544), .B(KEYINPUT4), .Z(n545) );
  NOR2_X1 U598 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U599 ( .A(KEYINPUT74), .B(n547), .Z(n548) );
  XNOR2_X1 U600 ( .A(KEYINPUT5), .B(n548), .ZN(n549) );
  NAND2_X1 U601 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U602 ( .A(KEYINPUT7), .B(n551), .ZN(G168) );
  XNOR2_X1 U603 ( .A(G168), .B(KEYINPUT8), .ZN(n552) );
  XNOR2_X1 U604 ( .A(n552), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U605 ( .A1(n883), .A2(G102), .ZN(n553) );
  XNOR2_X1 U606 ( .A(n553), .B(KEYINPUT86), .ZN(n555) );
  NAND2_X1 U607 ( .A1(G126), .A2(n878), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U609 ( .A1(G114), .A2(n877), .ZN(n557) );
  NAND2_X1 U610 ( .A1(G138), .A2(n773), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U612 ( .A1(n559), .A2(n558), .ZN(G164) );
  NAND2_X1 U613 ( .A1(G52), .A2(n784), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G64), .A2(n785), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n566) );
  NAND2_X1 U616 ( .A1(n780), .A2(G77), .ZN(n563) );
  NAND2_X1 U617 ( .A1(G90), .A2(n781), .ZN(n562) );
  NAND2_X1 U618 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U619 ( .A(KEYINPUT9), .B(n564), .Z(n565) );
  NOR2_X1 U620 ( .A1(n566), .A2(n565), .ZN(G171) );
  NAND2_X1 U621 ( .A1(n780), .A2(G78), .ZN(n568) );
  NAND2_X1 U622 ( .A1(G91), .A2(n781), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U624 ( .A1(G53), .A2(n784), .ZN(n570) );
  NAND2_X1 U625 ( .A1(G65), .A2(n785), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U627 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U628 ( .A(KEYINPUT68), .B(n573), .Z(G299) );
  NAND2_X1 U629 ( .A1(n780), .A2(G75), .ZN(n575) );
  NAND2_X1 U630 ( .A1(G88), .A2(n781), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n575), .A2(n574), .ZN(n580) );
  NAND2_X1 U632 ( .A1(n784), .A2(G50), .ZN(n576) );
  XNOR2_X1 U633 ( .A(n576), .B(KEYINPUT82), .ZN(n578) );
  NAND2_X1 U634 ( .A1(G62), .A2(n785), .ZN(n577) );
  NAND2_X1 U635 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U636 ( .A1(n580), .A2(n579), .ZN(G166) );
  INV_X1 U637 ( .A(G166), .ZN(G303) );
  NAND2_X1 U638 ( .A1(n581), .A2(G87), .ZN(n586) );
  NAND2_X1 U639 ( .A1(G49), .A2(n784), .ZN(n583) );
  NAND2_X1 U640 ( .A1(G74), .A2(G651), .ZN(n582) );
  NAND2_X1 U641 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U642 ( .A1(n785), .A2(n584), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U644 ( .A(KEYINPUT79), .B(n587), .Z(G288) );
  NAND2_X1 U645 ( .A1(G73), .A2(n780), .ZN(n588) );
  XNOR2_X1 U646 ( .A(n588), .B(KEYINPUT2), .ZN(n596) );
  NAND2_X1 U647 ( .A1(G61), .A2(n785), .ZN(n589) );
  XNOR2_X1 U648 ( .A(n589), .B(KEYINPUT80), .ZN(n591) );
  NAND2_X1 U649 ( .A1(G86), .A2(n781), .ZN(n590) );
  NAND2_X1 U650 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U651 ( .A1(G48), .A2(n784), .ZN(n592) );
  XNOR2_X1 U652 ( .A(KEYINPUT81), .B(n592), .ZN(n593) );
  NOR2_X1 U653 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U654 ( .A1(n596), .A2(n595), .ZN(G305) );
  NAND2_X1 U655 ( .A1(n780), .A2(G72), .ZN(n598) );
  NAND2_X1 U656 ( .A1(G85), .A2(n781), .ZN(n597) );
  NAND2_X1 U657 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U658 ( .A1(G47), .A2(n784), .ZN(n600) );
  NAND2_X1 U659 ( .A1(G60), .A2(n785), .ZN(n599) );
  NAND2_X1 U660 ( .A1(n600), .A2(n599), .ZN(n601) );
  OR2_X1 U661 ( .A1(n602), .A2(n601), .ZN(G290) );
  NAND2_X1 U662 ( .A1(G160), .A2(G40), .ZN(n604) );
  INV_X1 U663 ( .A(n709), .ZN(n605) );
  NOR2_X1 U664 ( .A1(G164), .A2(G1384), .ZN(n710) );
  INV_X1 U665 ( .A(G1961), .ZN(n996) );
  NAND2_X1 U666 ( .A1(n667), .A2(n996), .ZN(n608) );
  XNOR2_X1 U667 ( .A(G2078), .B(KEYINPUT92), .ZN(n606) );
  XNOR2_X1 U668 ( .A(n606), .B(KEYINPUT25), .ZN(n947) );
  NAND2_X1 U669 ( .A1(n639), .A2(n947), .ZN(n607) );
  NAND2_X1 U670 ( .A1(n608), .A2(n607), .ZN(n660) );
  NAND2_X1 U671 ( .A1(n660), .A2(G171), .ZN(n655) );
  NAND2_X1 U672 ( .A1(n639), .A2(G2072), .ZN(n609) );
  XNOR2_X1 U673 ( .A(n609), .B(KEYINPUT27), .ZN(n611) );
  INV_X1 U674 ( .A(G1956), .ZN(n997) );
  NOR2_X1 U675 ( .A1(n997), .A2(n639), .ZN(n610) );
  NOR2_X1 U676 ( .A1(n611), .A2(n610), .ZN(n615) );
  INV_X1 U677 ( .A(G299), .ZN(n614) );
  NOR2_X1 U678 ( .A1(n615), .A2(n614), .ZN(n613) );
  XNOR2_X1 U679 ( .A(KEYINPUT28), .B(KEYINPUT93), .ZN(n612) );
  XNOR2_X1 U680 ( .A(n613), .B(n612), .ZN(n651) );
  NAND2_X1 U681 ( .A1(n615), .A2(n614), .ZN(n649) );
  AND2_X1 U682 ( .A1(n639), .A2(G1996), .ZN(n617) );
  XOR2_X1 U683 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n616) );
  XNOR2_X1 U684 ( .A(n617), .B(n616), .ZN(n619) );
  NAND2_X1 U685 ( .A1(n667), .A2(G1341), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n619), .A2(n618), .ZN(n644) );
  NAND2_X1 U687 ( .A1(G81), .A2(n781), .ZN(n620) );
  XNOR2_X1 U688 ( .A(n620), .B(KEYINPUT12), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G68), .A2(n780), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U691 ( .A(n623), .B(KEYINPUT13), .ZN(n625) );
  NAND2_X1 U692 ( .A1(G43), .A2(n784), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U694 ( .A1(G56), .A2(n785), .ZN(n626) );
  XNOR2_X1 U695 ( .A(n626), .B(KEYINPUT14), .ZN(n627) );
  XNOR2_X1 U696 ( .A(n627), .B(KEYINPUT69), .ZN(n628) );
  NOR2_X1 U697 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U698 ( .A(KEYINPUT70), .B(n630), .ZN(n981) );
  NAND2_X1 U699 ( .A1(n780), .A2(G79), .ZN(n632) );
  NAND2_X1 U700 ( .A1(G92), .A2(n781), .ZN(n631) );
  NAND2_X1 U701 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U702 ( .A1(G54), .A2(n784), .ZN(n634) );
  NAND2_X1 U703 ( .A1(G66), .A2(n785), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U706 ( .A(KEYINPUT15), .B(n637), .Z(n638) );
  XNOR2_X1 U707 ( .A(KEYINPUT71), .B(n638), .ZN(n973) );
  NAND2_X1 U708 ( .A1(G1348), .A2(n667), .ZN(n641) );
  NAND2_X1 U709 ( .A1(G2067), .A2(n639), .ZN(n640) );
  NAND2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U711 ( .A1(n973), .A2(n645), .ZN(n642) );
  NAND2_X1 U712 ( .A1(n981), .A2(n642), .ZN(n643) );
  NOR2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n647) );
  NOR2_X1 U714 ( .A1(n645), .A2(n973), .ZN(n646) );
  NOR2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U718 ( .A(n652), .B(KEYINPUT29), .ZN(n653) );
  INV_X1 U719 ( .A(n653), .ZN(n654) );
  NAND2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n665) );
  NOR2_X1 U721 ( .A1(G1966), .A2(n706), .ZN(n678) );
  NOR2_X1 U722 ( .A1(G2084), .A2(n667), .ZN(n675) );
  NAND2_X1 U723 ( .A1(n656), .A2(G8), .ZN(n657) );
  XNOR2_X1 U724 ( .A(KEYINPUT30), .B(n658), .ZN(n659) );
  NOR2_X1 U725 ( .A1(G168), .A2(n659), .ZN(n662) );
  NOR2_X1 U726 ( .A1(G171), .A2(n660), .ZN(n661) );
  NOR2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U728 ( .A(KEYINPUT31), .B(n663), .Z(n664) );
  NAND2_X1 U729 ( .A1(n665), .A2(n664), .ZN(n676) );
  NAND2_X1 U730 ( .A1(G286), .A2(n676), .ZN(n666) );
  XNOR2_X1 U731 ( .A(n666), .B(KEYINPUT96), .ZN(n672) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n706), .ZN(n669) );
  NOR2_X1 U733 ( .A1(G2090), .A2(n667), .ZN(n668) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U735 ( .A1(n670), .A2(G303), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U737 ( .A1(n673), .A2(G8), .ZN(n674) );
  XNOR2_X1 U738 ( .A(n674), .B(KEYINPUT32), .ZN(n683) );
  NAND2_X1 U739 ( .A1(G8), .A2(n675), .ZN(n681) );
  INV_X1 U740 ( .A(n676), .ZN(n677) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U742 ( .A(KEYINPUT95), .B(n679), .Z(n680) );
  NAND2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U744 ( .A1(n683), .A2(n682), .ZN(n692) );
  NOR2_X1 U745 ( .A1(G2090), .A2(G303), .ZN(n684) );
  XOR2_X1 U746 ( .A(KEYINPUT97), .B(n684), .Z(n685) );
  NAND2_X1 U747 ( .A1(G8), .A2(n685), .ZN(n686) );
  NAND2_X1 U748 ( .A1(n692), .A2(n686), .ZN(n687) );
  NAND2_X1 U749 ( .A1(n687), .A2(n706), .ZN(n701) );
  NOR2_X1 U750 ( .A1(G1976), .A2(G288), .ZN(n970) );
  NOR2_X1 U751 ( .A1(G1971), .A2(G303), .ZN(n688) );
  NOR2_X1 U752 ( .A1(n970), .A2(n688), .ZN(n690) );
  INV_X1 U753 ( .A(KEYINPUT33), .ZN(n689) );
  AND2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n699) );
  XOR2_X1 U756 ( .A(G1981), .B(G305), .Z(n987) );
  NAND2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n971) );
  INV_X1 U758 ( .A(n971), .ZN(n693) );
  NOR2_X1 U759 ( .A1(KEYINPUT33), .A2(n521), .ZN(n696) );
  NAND2_X1 U760 ( .A1(n970), .A2(KEYINPUT33), .ZN(n694) );
  NOR2_X1 U761 ( .A1(n706), .A2(n694), .ZN(n695) );
  NOR2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U763 ( .A1(n987), .A2(n697), .ZN(n698) );
  NAND2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U766 ( .A(n702), .B(KEYINPUT98), .ZN(n708) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n703) );
  XNOR2_X1 U768 ( .A(n703), .B(KEYINPUT24), .ZN(n704) );
  XNOR2_X1 U769 ( .A(n704), .B(KEYINPUT91), .ZN(n705) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U771 ( .A1(n710), .A2(n709), .ZN(n752) );
  XNOR2_X1 U772 ( .A(KEYINPUT37), .B(G2067), .ZN(n750) );
  NAND2_X1 U773 ( .A1(G104), .A2(n883), .ZN(n712) );
  NAND2_X1 U774 ( .A1(G140), .A2(n773), .ZN(n711) );
  NAND2_X1 U775 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U776 ( .A(KEYINPUT34), .B(n713), .ZN(n719) );
  NAND2_X1 U777 ( .A1(G116), .A2(n877), .ZN(n715) );
  NAND2_X1 U778 ( .A1(G128), .A2(n878), .ZN(n714) );
  NAND2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U780 ( .A(KEYINPUT88), .B(n716), .Z(n717) );
  XNOR2_X1 U781 ( .A(KEYINPUT35), .B(n717), .ZN(n718) );
  NOR2_X1 U782 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U783 ( .A(n720), .B(KEYINPUT36), .Z(n721) );
  XNOR2_X1 U784 ( .A(KEYINPUT89), .B(n721), .ZN(n891) );
  NOR2_X1 U785 ( .A1(n750), .A2(n891), .ZN(n926) );
  NAND2_X1 U786 ( .A1(n752), .A2(n926), .ZN(n748) );
  NAND2_X1 U787 ( .A1(G119), .A2(n878), .ZN(n723) );
  NAND2_X1 U788 ( .A1(G131), .A2(n773), .ZN(n722) );
  NAND2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n727) );
  NAND2_X1 U790 ( .A1(G107), .A2(n877), .ZN(n725) );
  NAND2_X1 U791 ( .A1(G95), .A2(n883), .ZN(n724) );
  NAND2_X1 U792 ( .A1(n725), .A2(n724), .ZN(n726) );
  OR2_X1 U793 ( .A1(n727), .A2(n726), .ZN(n865) );
  AND2_X1 U794 ( .A1(n865), .A2(G1991), .ZN(n737) );
  NAND2_X1 U795 ( .A1(G129), .A2(n878), .ZN(n729) );
  NAND2_X1 U796 ( .A1(G141), .A2(n773), .ZN(n728) );
  NAND2_X1 U797 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U798 ( .A1(n883), .A2(G105), .ZN(n730) );
  XOR2_X1 U799 ( .A(KEYINPUT38), .B(n730), .Z(n731) );
  NOR2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U801 ( .A1(n877), .A2(G117), .ZN(n733) );
  NAND2_X1 U802 ( .A1(n734), .A2(n733), .ZN(n861) );
  NAND2_X1 U803 ( .A1(G1996), .A2(n861), .ZN(n735) );
  XOR2_X1 U804 ( .A(KEYINPUT90), .B(n735), .Z(n736) );
  NOR2_X1 U805 ( .A1(n737), .A2(n736), .ZN(n928) );
  INV_X1 U806 ( .A(n928), .ZN(n738) );
  NAND2_X1 U807 ( .A1(n738), .A2(n752), .ZN(n741) );
  XNOR2_X1 U808 ( .A(G1986), .B(G290), .ZN(n978) );
  NAND2_X1 U809 ( .A1(n752), .A2(n978), .ZN(n739) );
  NAND2_X1 U810 ( .A1(n522), .A2(n524), .ZN(n740) );
  XOR2_X1 U811 ( .A(KEYINPUT99), .B(n740), .Z(n755) );
  NOR2_X1 U812 ( .A1(G1996), .A2(n861), .ZN(n931) );
  INV_X1 U813 ( .A(n741), .ZN(n744) );
  NOR2_X1 U814 ( .A1(G1991), .A2(n865), .ZN(n922) );
  NOR2_X1 U815 ( .A1(G1986), .A2(G290), .ZN(n742) );
  NOR2_X1 U816 ( .A1(n922), .A2(n742), .ZN(n743) );
  NOR2_X1 U817 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U818 ( .A(n745), .B(KEYINPUT100), .ZN(n746) );
  NOR2_X1 U819 ( .A1(n931), .A2(n746), .ZN(n747) );
  XNOR2_X1 U820 ( .A(n747), .B(KEYINPUT39), .ZN(n749) );
  NAND2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n751) );
  NAND2_X1 U822 ( .A1(n750), .A2(n891), .ZN(n934) );
  NAND2_X1 U823 ( .A1(n751), .A2(n934), .ZN(n753) );
  NAND2_X1 U824 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U825 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U826 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U827 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U828 ( .A(G57), .ZN(G237) );
  NAND2_X1 U829 ( .A1(G7), .A2(G661), .ZN(n757) );
  XNOR2_X1 U830 ( .A(n757), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U831 ( .A(G223), .ZN(n823) );
  NAND2_X1 U832 ( .A1(n823), .A2(G567), .ZN(n758) );
  XOR2_X1 U833 ( .A(KEYINPUT11), .B(n758), .Z(G234) );
  NAND2_X1 U834 ( .A1(G860), .A2(n981), .ZN(G153) );
  INV_X1 U835 ( .A(G171), .ZN(G301) );
  INV_X1 U836 ( .A(G868), .ZN(n804) );
  NAND2_X1 U837 ( .A1(n973), .A2(n804), .ZN(n759) );
  XNOR2_X1 U838 ( .A(n759), .B(KEYINPUT72), .ZN(n761) );
  NAND2_X1 U839 ( .A1(G868), .A2(G301), .ZN(n760) );
  NAND2_X1 U840 ( .A1(n761), .A2(n760), .ZN(G284) );
  NOR2_X1 U841 ( .A1(G286), .A2(n804), .ZN(n763) );
  NOR2_X1 U842 ( .A1(G299), .A2(G868), .ZN(n762) );
  NOR2_X1 U843 ( .A1(n763), .A2(n762), .ZN(G297) );
  INV_X1 U844 ( .A(G860), .ZN(n764) );
  NAND2_X1 U845 ( .A1(n764), .A2(G559), .ZN(n765) );
  INV_X1 U846 ( .A(n973), .ZN(n791) );
  NAND2_X1 U847 ( .A1(n765), .A2(n791), .ZN(n766) );
  XNOR2_X1 U848 ( .A(n766), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U849 ( .A1(n791), .A2(G868), .ZN(n767) );
  NOR2_X1 U850 ( .A1(G559), .A2(n767), .ZN(n769) );
  AND2_X1 U851 ( .A1(n981), .A2(n804), .ZN(n768) );
  NOR2_X1 U852 ( .A1(n769), .A2(n768), .ZN(G282) );
  NAND2_X1 U853 ( .A1(G123), .A2(n878), .ZN(n770) );
  XNOR2_X1 U854 ( .A(n770), .B(KEYINPUT18), .ZN(n772) );
  NAND2_X1 U855 ( .A1(n883), .A2(G99), .ZN(n771) );
  NAND2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n777) );
  NAND2_X1 U857 ( .A1(G111), .A2(n877), .ZN(n775) );
  BUF_X1 U858 ( .A(n773), .Z(n881) );
  NAND2_X1 U859 ( .A1(G135), .A2(n881), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n921) );
  XNOR2_X1 U862 ( .A(n921), .B(G2096), .ZN(n779) );
  INV_X1 U863 ( .A(G2100), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n779), .A2(n778), .ZN(G156) );
  NAND2_X1 U865 ( .A1(n780), .A2(G80), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G93), .A2(n781), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n790) );
  NAND2_X1 U868 ( .A1(G55), .A2(n784), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G67), .A2(n785), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U871 ( .A(KEYINPUT77), .B(n788), .Z(n789) );
  NOR2_X1 U872 ( .A1(n790), .A2(n789), .ZN(n803) );
  XNOR2_X1 U873 ( .A(KEYINPUT76), .B(KEYINPUT78), .ZN(n794) );
  NAND2_X1 U874 ( .A1(G559), .A2(n791), .ZN(n792) );
  XOR2_X1 U875 ( .A(n981), .B(n792), .Z(n801) );
  NOR2_X1 U876 ( .A1(n801), .A2(G860), .ZN(n793) );
  XNOR2_X1 U877 ( .A(n794), .B(n793), .ZN(n795) );
  XNOR2_X1 U878 ( .A(n803), .B(n795), .ZN(G145) );
  XNOR2_X1 U879 ( .A(G166), .B(G288), .ZN(n798) );
  XNOR2_X1 U880 ( .A(G299), .B(n803), .ZN(n796) );
  XNOR2_X1 U881 ( .A(n796), .B(G305), .ZN(n797) );
  XNOR2_X1 U882 ( .A(n798), .B(n797), .ZN(n799) );
  XNOR2_X1 U883 ( .A(KEYINPUT19), .B(n799), .ZN(n800) );
  XNOR2_X1 U884 ( .A(n800), .B(G290), .ZN(n894) );
  XNOR2_X1 U885 ( .A(n894), .B(n801), .ZN(n802) );
  NAND2_X1 U886 ( .A1(n802), .A2(G868), .ZN(n806) );
  NAND2_X1 U887 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U888 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U889 ( .A(KEYINPUT83), .B(n807), .ZN(G295) );
  NAND2_X1 U890 ( .A1(G2084), .A2(G2078), .ZN(n808) );
  XOR2_X1 U891 ( .A(KEYINPUT20), .B(n808), .Z(n809) );
  NAND2_X1 U892 ( .A1(G2090), .A2(n809), .ZN(n810) );
  XNOR2_X1 U893 ( .A(KEYINPUT21), .B(n810), .ZN(n811) );
  NAND2_X1 U894 ( .A1(n811), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U895 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U896 ( .A1(G132), .A2(G82), .ZN(n812) );
  XNOR2_X1 U897 ( .A(n812), .B(KEYINPUT22), .ZN(n813) );
  XNOR2_X1 U898 ( .A(n813), .B(KEYINPUT84), .ZN(n814) );
  NOR2_X1 U899 ( .A1(G218), .A2(n814), .ZN(n815) );
  NAND2_X1 U900 ( .A1(G96), .A2(n815), .ZN(n829) );
  NAND2_X1 U901 ( .A1(G2106), .A2(n829), .ZN(n819) );
  NAND2_X1 U902 ( .A1(G69), .A2(G120), .ZN(n816) );
  NOR2_X1 U903 ( .A1(G237), .A2(n816), .ZN(n817) );
  NAND2_X1 U904 ( .A1(G108), .A2(n817), .ZN(n830) );
  NAND2_X1 U905 ( .A1(G567), .A2(n830), .ZN(n818) );
  NAND2_X1 U906 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U907 ( .A(KEYINPUT85), .B(n820), .ZN(G319) );
  INV_X1 U908 ( .A(G319), .ZN(n822) );
  NAND2_X1 U909 ( .A1(G661), .A2(G483), .ZN(n821) );
  NOR2_X1 U910 ( .A1(n822), .A2(n821), .ZN(n828) );
  NAND2_X1 U911 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n823), .ZN(G217) );
  NAND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n824) );
  XOR2_X1 U914 ( .A(KEYINPUT102), .B(n824), .Z(n825) );
  NAND2_X1 U915 ( .A1(n825), .A2(G661), .ZN(n826) );
  XOR2_X1 U916 ( .A(KEYINPUT103), .B(n826), .Z(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n828), .A2(n827), .ZN(G188) );
  INV_X1 U920 ( .A(G132), .ZN(G219) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G82), .ZN(G220) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  XOR2_X1 U926 ( .A(G2096), .B(G2072), .Z(n832) );
  XNOR2_X1 U927 ( .A(G2067), .B(G2090), .ZN(n831) );
  XNOR2_X1 U928 ( .A(n832), .B(n831), .ZN(n842) );
  XOR2_X1 U929 ( .A(KEYINPUT105), .B(G2678), .Z(n834) );
  XNOR2_X1 U930 ( .A(G2100), .B(KEYINPUT107), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U932 ( .A(KEYINPUT104), .B(KEYINPUT106), .Z(n836) );
  XNOR2_X1 U933 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U935 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U936 ( .A(G2084), .B(G2078), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U938 ( .A(n842), .B(n841), .Z(G227) );
  XOR2_X1 U939 ( .A(G1956), .B(G1966), .Z(n844) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1981), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(n845), .B(G2474), .Z(n847) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U945 ( .A(KEYINPUT41), .B(G1976), .Z(n849) );
  XNOR2_X1 U946 ( .A(G1961), .B(G1971), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(G229) );
  NAND2_X1 U949 ( .A1(n878), .A2(G124), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n852), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G136), .A2(n881), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(KEYINPUT108), .B(n855), .Z(n857) );
  NAND2_X1 U954 ( .A1(n883), .A2(G100), .ZN(n856) );
  NAND2_X1 U955 ( .A1(n857), .A2(n856), .ZN(n860) );
  NAND2_X1 U956 ( .A1(G112), .A2(n877), .ZN(n858) );
  XNOR2_X1 U957 ( .A(KEYINPUT109), .B(n858), .ZN(n859) );
  NOR2_X1 U958 ( .A1(n860), .A2(n859), .ZN(G162) );
  XNOR2_X1 U959 ( .A(n861), .B(n921), .ZN(n863) );
  XNOR2_X1 U960 ( .A(G160), .B(G164), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U962 ( .A(n865), .B(n864), .Z(n876) );
  XOR2_X1 U963 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n874) );
  NAND2_X1 U964 ( .A1(G103), .A2(n883), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G139), .A2(n881), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U967 ( .A1(G115), .A2(n877), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G127), .A2(n878), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n870), .Z(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n917) );
  XNOR2_X1 U972 ( .A(G162), .B(n917), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n890) );
  NAND2_X1 U975 ( .A1(G118), .A2(n877), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G130), .A2(n878), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n888) );
  NAND2_X1 U978 ( .A1(G142), .A2(n881), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n882), .B(KEYINPUT110), .ZN(n885) );
  NAND2_X1 U980 ( .A1(G106), .A2(n883), .ZN(n884) );
  NAND2_X1 U981 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U982 ( .A(n886), .B(KEYINPUT45), .Z(n887) );
  NOR2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U984 ( .A(n890), .B(n889), .Z(n892) );
  XOR2_X1 U985 ( .A(n892), .B(n891), .Z(n893) );
  NOR2_X1 U986 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U987 ( .A(G171), .B(n973), .ZN(n895) );
  XNOR2_X1 U988 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U989 ( .A(G286), .B(n896), .ZN(n897) );
  XNOR2_X1 U990 ( .A(n897), .B(n981), .ZN(n898) );
  NOR2_X1 U991 ( .A1(G37), .A2(n898), .ZN(G397) );
  XOR2_X1 U992 ( .A(G2454), .B(G2435), .Z(n900) );
  XNOR2_X1 U993 ( .A(G2438), .B(G2427), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n907) );
  XOR2_X1 U995 ( .A(KEYINPUT101), .B(G2446), .Z(n902) );
  XNOR2_X1 U996 ( .A(G2443), .B(G2430), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U998 ( .A(n903), .B(G2451), .Z(n905) );
  XNOR2_X1 U999 ( .A(G1348), .B(G1341), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1002 ( .A1(n908), .A2(G14), .ZN(n915) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n915), .ZN(n912) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n909) );
  XOR2_X1 U1005 ( .A(KEYINPUT111), .B(n909), .Z(n910) );
  XNOR2_X1 U1006 ( .A(n910), .B(KEYINPUT49), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  INV_X1 U1012 ( .A(G96), .ZN(G221) );
  INV_X1 U1013 ( .A(n915), .ZN(G401) );
  XNOR2_X1 U1014 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(n916), .B(KEYINPUT52), .ZN(n942) );
  XOR2_X1 U1016 ( .A(G2072), .B(n917), .Z(n919) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1019 ( .A(KEYINPUT50), .B(n920), .Z(n940) );
  XNOR2_X1 U1020 ( .A(G160), .B(G2084), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1025 ( .A(KEYINPUT112), .B(n929), .ZN(n937) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(KEYINPUT113), .B(n932), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(n933), .B(KEYINPUT51), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1032 ( .A(KEYINPUT114), .B(n938), .Z(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n942), .B(n941), .ZN(n943) );
  NOR2_X1 U1035 ( .A1(KEYINPUT55), .A2(n943), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(KEYINPUT117), .B(n944), .ZN(n945) );
  NAND2_X1 U1037 ( .A1(n945), .A2(G29), .ZN(n1027) );
  XNOR2_X1 U1038 ( .A(G1996), .B(KEYINPUT119), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(n946), .B(G32), .ZN(n951) );
  XOR2_X1 U1040 ( .A(n947), .B(G27), .Z(n949) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n954) );
  XNOR2_X1 U1044 ( .A(KEYINPUT118), .B(G2067), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G26), .B(n952), .ZN(n953) );
  NOR2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1047 ( .A(KEYINPUT120), .B(n955), .Z(n957) );
  XNOR2_X1 U1048 ( .A(G1991), .B(G25), .ZN(n956) );
  NOR2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1050 ( .A1(G28), .A2(n958), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(n959), .B(KEYINPUT53), .ZN(n962) );
  XOR2_X1 U1052 ( .A(G2084), .B(G34), .Z(n960) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(n960), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(G35), .B(G2090), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1057 ( .A(KEYINPUT55), .B(n965), .Z(n966) );
  NOR2_X1 U1058 ( .A1(G29), .A2(n966), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT121), .B(n967), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(n968), .A2(G11), .ZN(n1025) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XNOR2_X1 U1062 ( .A(G299), .B(G1956), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(G1348), .B(n973), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n985) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G166), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(KEYINPUT124), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G1961), .B(G301), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n983) );
  XOR2_X1 U1072 ( .A(G1341), .B(n981), .Z(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(n986), .B(KEYINPUT125), .ZN(n993) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(n989), .B(KEYINPUT123), .ZN(n991) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n990) );
  XNOR2_X1 U1080 ( .A(n991), .B(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n1023) );
  INV_X1 U1083 ( .A(G16), .ZN(n1021) );
  XNOR2_X1 U1084 ( .A(G5), .B(n996), .ZN(n1016) );
  XOR2_X1 U1085 ( .A(G1981), .B(G6), .Z(n999) );
  XNOR2_X1 U1086 ( .A(n997), .B(G20), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(G19), .B(G1341), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(KEYINPUT126), .B(n1002), .ZN(n1006) );
  XOR2_X1 U1091 ( .A(G4), .B(KEYINPUT127), .Z(n1004) );
  XNOR2_X1 U1092 ( .A(G1348), .B(KEYINPUT59), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1004), .B(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1007), .B(KEYINPUT60), .ZN(n1014) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(G23), .B(G1976), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(G1986), .B(G24), .Z(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(G21), .B(G1966), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

