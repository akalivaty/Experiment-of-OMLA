//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT93), .Z(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT91), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT14), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT92), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(KEYINPUT90), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n211), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n215), .A2(KEYINPUT90), .ZN(new_n221));
  OAI211_X1 g020(.A(KEYINPUT15), .B(new_n209), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n208), .B(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225));
  XOR2_X1   g024(.A(new_n225), .B(KEYINPUT13), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n223), .A2(new_n228), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n208), .A2(new_n223), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n233), .A3(new_n225), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n227), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT94), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n235), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(new_n237), .B2(new_n238), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT89), .ZN(new_n242));
  XOR2_X1   g041(.A(G113gat), .B(G141gat), .Z(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G169gat), .B(G197gat), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n244), .B(new_n245), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT12), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n240), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT95), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n238), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT95), .B1(new_n234), .B2(new_n235), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n227), .B(new_n247), .C1(new_n234), .C2(new_n235), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT96), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT96), .ZN(new_n257));
  NOR4_X1   g056(.A1(new_n251), .A2(new_n254), .A3(new_n252), .A4(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n249), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT24), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(G183gat), .A3(G190gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(G183gat), .A2(G190gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n261), .B1(new_n263), .B2(new_n260), .ZN(new_n264));
  INV_X1    g063(.A(G183gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G183gat), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT67), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G190gat), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n269), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(new_n269), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n264), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT23), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n279), .B1(KEYINPUT23), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n278), .A2(KEYINPUT25), .A3(new_n280), .A4(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT25), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n282), .B1(new_n286), .B2(new_n280), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n279), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n265), .A2(new_n270), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n264), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT64), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n287), .B(new_n288), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n290), .A2(new_n291), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n285), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n284), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n297));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G183gat), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n271), .A2(new_n273), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT27), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n265), .A2(KEYINPUT27), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n271), .A2(new_n273), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n296), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT27), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n271), .A2(new_n273), .A3(new_n299), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n274), .A2(KEYINPUT28), .A3(new_n299), .A4(new_n303), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(KEYINPUT70), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n279), .A2(KEYINPUT26), .ZN(new_n316));
  INV_X1    g115(.A(new_n281), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n263), .B1(KEYINPUT26), .B2(new_n279), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT71), .B1(new_n315), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n323));
  AOI211_X1 g122(.A(new_n323), .B(new_n320), .C1(new_n308), .C2(new_n314), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n295), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT72), .B(G134gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G127gat), .ZN(new_n328));
  INV_X1    g127(.A(G113gat), .ZN(new_n329));
  INV_X1    g128(.A(G120gat), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT1), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n329), .B2(new_n330), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n328), .B(new_n332), .C1(G127gat), .C2(G134gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT73), .B(G120gat), .Z(new_n335));
  OAI211_X1 g134(.A(new_n331), .B(new_n334), .C1(new_n335), .C2(new_n329), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n325), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n337), .B(new_n295), .C1(new_n322), .C2(new_n324), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G227gat), .ZN(new_n342));
  INV_X1    g141(.A(G233gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(KEYINPUT77), .B(KEYINPUT34), .Z(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT32), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n342), .A2(new_n343), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n339), .A2(new_n349), .A3(new_n340), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT74), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n339), .A2(new_n352), .A3(new_n349), .A4(new_n340), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n348), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G15gat), .B(G43gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n361), .B1(new_n354), .B2(new_n355), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n351), .A2(new_n353), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT33), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI211_X1 g166(.A(KEYINPUT75), .B(KEYINPUT33), .C1(new_n351), .C2(new_n353), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n354), .B1(new_n366), .B2(new_n360), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n347), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n365), .A2(KEYINPUT32), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT76), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(new_n361), .A3(new_n356), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n367), .A2(new_n368), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n371), .B(new_n347), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379));
  XOR2_X1   g178(.A(G155gat), .B(G162gat), .Z(new_n380));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G155gat), .ZN(new_n383));
  INV_X1    g182(.A(G162gat), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT2), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G141gat), .B(G148gat), .Z(new_n386));
  NAND2_X1  g185(.A1(new_n380), .A2(new_n381), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(KEYINPUT81), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n386), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n385), .A2(KEYINPUT81), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n380), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G197gat), .B(G204gat), .ZN(new_n394));
  INV_X1    g193(.A(G211gat), .ZN(new_n395));
  INV_X1    g194(.A(G218gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n394), .B1(KEYINPUT22), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G211gat), .B(G218gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(KEYINPUT29), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n393), .B1(new_n401), .B2(KEYINPUT3), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n379), .B1(new_n403), .B2(KEYINPUT83), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n393), .A2(KEYINPUT3), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n400), .B1(new_n405), .B2(KEYINPUT29), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n402), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n408), .B(new_n379), .C1(KEYINPUT83), .C2(new_n403), .ZN(new_n409));
  INV_X1    g208(.A(G22gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT84), .ZN(new_n412));
  XOR2_X1   g211(.A(G78gat), .B(G106gat), .Z(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT31), .B(G50gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n407), .A2(new_n409), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G22gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n411), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n416), .B(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n372), .A2(new_n378), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT78), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n325), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n423), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n284), .A2(new_n294), .B1(new_n315), .B2(new_n321), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(KEYINPUT29), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT79), .B1(new_n428), .B2(new_n400), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n423), .B1(new_n325), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n426), .A2(new_n425), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n400), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT79), .ZN(new_n434));
  INV_X1    g233(.A(new_n400), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n424), .A2(new_n427), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G8gat), .B(G36gat), .Z(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT80), .ZN(new_n438));
  XNOR2_X1  g237(.A(G64gat), .B(G92gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n429), .A2(new_n433), .A3(new_n436), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n433), .A3(new_n436), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n440), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n442), .A2(new_n443), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n338), .A2(KEYINPUT4), .A3(new_n392), .A4(new_n388), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT4), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n393), .B2(new_n337), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G225gat), .A2(G233gat), .ZN(new_n457));
  INV_X1    g256(.A(new_n405), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n393), .A2(KEYINPUT3), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n337), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n456), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n393), .B(new_n337), .ZN(new_n462));
  INV_X1    g261(.A(new_n457), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n456), .A2(KEYINPUT5), .A3(new_n457), .A4(new_n460), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G1gat), .B(G29gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT0), .ZN(new_n470));
  XNOR2_X1  g269(.A(G57gat), .B(G85gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  AOI21_X1  g271(.A(KEYINPUT6), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n472), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n466), .A2(new_n474), .A3(new_n467), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT86), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n466), .A2(KEYINPUT86), .A3(new_n474), .A4(new_n467), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n466), .A2(KEYINPUT6), .A3(new_n474), .A4(new_n467), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n451), .A2(new_n482), .A3(KEYINPUT35), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n371), .B1(new_n375), .B2(new_n376), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n346), .ZN(new_n485));
  INV_X1    g284(.A(new_n420), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n473), .A2(new_n475), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n487), .A2(new_n480), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n488), .A2(new_n449), .A3(new_n447), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n485), .A2(new_n377), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n421), .A2(new_n483), .B1(new_n490), .B2(KEYINPUT35), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n477), .A2(new_n478), .ZN(new_n492));
  INV_X1    g291(.A(new_n460), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n463), .B1(new_n493), .B2(new_n455), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT39), .B1(new_n462), .B2(new_n463), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT85), .B(KEYINPUT39), .C1(new_n462), .C2(new_n463), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n457), .B1(new_n456), .B2(new_n460), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT39), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n474), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n499), .A2(new_n502), .A3(KEYINPUT40), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT40), .B1(new_n499), .B2(new_n502), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n492), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n449), .B2(new_n447), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n486), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n479), .A2(new_n480), .A3(new_n442), .ZN(new_n508));
  XOR2_X1   g307(.A(KEYINPUT87), .B(KEYINPUT38), .Z(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n445), .B2(KEYINPUT37), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n510), .B(new_n440), .C1(KEYINPUT37), .C2(new_n445), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n435), .B1(new_n431), .B2(new_n432), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n512), .B(KEYINPUT37), .C1(new_n435), .C2(new_n428), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n440), .B(new_n513), .C1(new_n445), .C2(KEYINPUT37), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n509), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n508), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  OAI22_X1  g315(.A1(new_n507), .A2(new_n516), .B1(new_n486), .B2(new_n489), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(new_n372), .B2(new_n378), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n485), .A2(KEYINPUT36), .A3(new_n377), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n259), .B1(new_n491), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT97), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n490), .A2(KEYINPUT35), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n483), .A2(new_n485), .A3(new_n377), .A4(new_n486), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n420), .B1(new_n451), .B2(new_n505), .ZN(new_n528));
  INV_X1    g327(.A(new_n516), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n487), .A2(new_n480), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n448), .A2(new_n530), .A3(new_n450), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n528), .A2(new_n529), .B1(new_n420), .B2(new_n531), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n485), .A2(KEYINPUT36), .A3(new_n377), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT36), .B1(new_n485), .B2(new_n377), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(KEYINPUT97), .A3(new_n259), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n524), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G71gat), .A2(G78gat), .ZN(new_n539));
  OR2_X1    g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT9), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G64gat), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT98), .B1(new_n543), .B2(G57gat), .ZN(new_n544));
  INV_X1    g343(.A(G57gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n545), .B2(G64gat), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n543), .A2(KEYINPUT98), .A3(G57gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G57gat), .B(G64gat), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n539), .B(new_n540), .C1(new_n549), .C2(new_n541), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT99), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT100), .B(KEYINPUT21), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G127gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n552), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n208), .B1(KEYINPUT21), .B2(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n557), .B(new_n559), .Z(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT101), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G155gat), .ZN(new_n563));
  XOR2_X1   g362(.A(G183gat), .B(G211gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n560), .B(new_n565), .Z(new_n566));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(KEYINPUT102), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(KEYINPUT102), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n568), .A2(new_n569), .A3(G85gat), .A4(G92gat), .ZN(new_n570));
  INV_X1    g369(.A(G85gat), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  OAI211_X1 g371(.A(KEYINPUT102), .B(new_n567), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G99gat), .A2(G106gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n574), .B1(new_n571), .B2(new_n572), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G99gat), .B(G106gat), .Z(new_n577));
  OR2_X1    g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n223), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n229), .A2(new_n580), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n231), .ZN(new_n585));
  XOR2_X1   g384(.A(G190gat), .B(G218gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G134gat), .B(G162gat), .Z(new_n588));
  AOI21_X1  g387(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT103), .Z(new_n591));
  OR2_X1    g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(KEYINPUT103), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n566), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n558), .A2(new_n581), .A3(KEYINPUT10), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n580), .B1(new_n548), .B2(new_n550), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n600), .B1(new_n558), .B2(new_n580), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n599), .B1(new_n601), .B2(KEYINPUT10), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT104), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n598), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(new_n603), .B2(new_n602), .ZN(new_n605));
  XNOR2_X1  g404(.A(G120gat), .B(G148gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT105), .ZN(new_n607));
  XNOR2_X1  g406(.A(G176gat), .B(G204gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n601), .A2(new_n598), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n602), .A2(new_n597), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n611), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n609), .B(KEYINPUT106), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n596), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n538), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n488), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g423(.A(new_n206), .B1(new_n622), .B2(new_n451), .ZN(new_n625));
  INV_X1    g424(.A(new_n451), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT16), .B(G8gat), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n621), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT42), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(KEYINPUT42), .B2(new_n628), .ZN(G1325gat));
  NAND2_X1  g429(.A1(new_n485), .A2(new_n377), .ZN(new_n631));
  OR3_X1    g430(.A1(new_n621), .A2(G15gat), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT107), .B1(new_n533), .B2(new_n534), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT107), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n519), .A2(new_n634), .A3(new_n520), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(G15gat), .B1(new_n621), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n632), .A2(new_n638), .ZN(G1326gat));
  NAND3_X1  g438(.A1(new_n622), .A2(KEYINPUT108), .A3(new_n420), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT108), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(new_n621), .B2(new_n486), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT43), .B(G22gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(G1327gat));
  NAND3_X1  g444(.A1(new_n566), .A2(new_n595), .A3(new_n618), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(KEYINPUT109), .Z(new_n647));
  NAND2_X1  g446(.A1(new_n538), .A2(new_n647), .ZN(new_n648));
  OR3_X1    g447(.A1(new_n648), .A2(G29gat), .A3(new_n530), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n595), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n633), .A2(new_n635), .A3(new_n532), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n653), .B1(new_n654), .B2(new_n527), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n652), .B1(new_n536), .B2(new_n595), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n566), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n238), .B(new_n250), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n257), .B1(new_n659), .B2(new_n254), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n253), .A2(KEYINPUT96), .A3(new_n255), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n660), .A2(new_n661), .B1(new_n240), .B2(new_n248), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n658), .A2(new_n662), .A3(new_n617), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G29gat), .B1(new_n664), .B2(new_n530), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n665), .A3(new_n666), .ZN(G1328gat));
  OR3_X1    g466(.A1(new_n648), .A2(G36gat), .A3(new_n626), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT46), .ZN(new_n669));
  OAI21_X1  g468(.A(G36gat), .B1(new_n664), .B2(new_n626), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(KEYINPUT46), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(G1329gat));
  OAI21_X1  g471(.A(G43gat), .B1(new_n664), .B2(new_n637), .ZN(new_n673));
  OR3_X1    g472(.A1(new_n648), .A2(G43gat), .A3(new_n631), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g475(.A(KEYINPUT48), .ZN(new_n677));
  INV_X1    g476(.A(new_n647), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n524), .B2(new_n537), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n486), .A2(G50gat), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n420), .B(new_n663), .C1(new_n655), .C2(new_n656), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(G50gat), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n681), .A2(new_n683), .A3(KEYINPUT112), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT112), .B1(new_n681), .B2(new_n683), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n680), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n687), .B(new_n678), .C1(new_n524), .C2(new_n537), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n683), .B2(KEYINPUT111), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT111), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n682), .A2(new_n690), .A3(G50gat), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT48), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT113), .B1(new_n686), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n683), .A2(KEYINPUT111), .ZN(new_n694));
  INV_X1    g493(.A(new_n688), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n677), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n683), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT112), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n681), .A2(new_n683), .A3(KEYINPUT112), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT113), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n697), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n693), .A2(new_n704), .ZN(G1331gat));
  NAND3_X1  g504(.A1(new_n596), .A2(new_n662), .A3(new_n617), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n654), .B2(new_n527), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n488), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g508(.A(new_n451), .B(KEYINPUT114), .Z(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT49), .B(G64gat), .Z(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT115), .ZN(G1333gat));
  NAND2_X1  g515(.A1(new_n707), .A2(new_n636), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n631), .A2(G71gat), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n717), .A2(G71gat), .B1(new_n707), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g519(.A1(new_n707), .A2(new_n420), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g521(.A1(new_n259), .A2(new_n658), .A3(new_n618), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n657), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(G85gat), .B1(new_n724), .B2(new_n530), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n654), .A2(new_n527), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n726), .A2(new_n662), .A3(new_n566), .A4(new_n595), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT51), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n488), .A2(new_n571), .A3(new_n617), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(G1336gat));
  INV_X1    g529(.A(new_n728), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n710), .A2(G92gat), .A3(new_n618), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT52), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G92gat), .B1(new_n724), .B2(new_n710), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n724), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n572), .B1(new_n736), .B2(new_n451), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT117), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n727), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n727), .A2(new_n738), .A3(KEYINPUT51), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n732), .B(KEYINPUT116), .Z(new_n743));
  AND3_X1   g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT52), .B1(new_n737), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n735), .A2(new_n745), .ZN(G1337gat));
  OAI21_X1  g545(.A(G99gat), .B1(new_n724), .B2(new_n637), .ZN(new_n747));
  OR3_X1    g546(.A1(new_n631), .A2(G99gat), .A3(new_n618), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n728), .B2(new_n748), .ZN(G1338gat));
  NOR3_X1   g548(.A1(new_n486), .A2(G106gat), .A3(new_n618), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT53), .B1(new_n731), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n657), .A2(new_n420), .A3(new_n723), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT119), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G106gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n752), .A2(KEYINPUT119), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n752), .A2(KEYINPUT118), .A3(G106gat), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n741), .A2(new_n742), .A3(new_n750), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT118), .B1(new_n752), .B2(G106gat), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n756), .B1(new_n760), .B2(new_n761), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n620), .A2(new_n662), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n602), .A2(new_n597), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(KEYINPUT54), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n765), .A2(new_n605), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n609), .B1(new_n613), .B2(KEYINPUT54), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT55), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n766), .B2(new_n767), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n769), .A2(new_n595), .A3(new_n612), .A4(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n246), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n232), .A2(new_n233), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(G229gat), .A3(G233gat), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n224), .A2(new_n226), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n773), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n256), .B2(new_n258), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n772), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n617), .B(new_n779), .C1(new_n256), .C2(new_n258), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n769), .A2(new_n612), .A3(new_n771), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n662), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n595), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n763), .B1(new_n786), .B2(new_n658), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n486), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n711), .A2(new_n530), .ZN(new_n789));
  INV_X1    g588(.A(new_n631), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n329), .B1(new_n792), .B2(new_n259), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT120), .Z(new_n794));
  INV_X1    g593(.A(new_n787), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(new_n530), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n796), .A2(new_n421), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n710), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n259), .A2(new_n329), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n798), .B2(new_n799), .ZN(G1340gat));
  INV_X1    g599(.A(new_n792), .ZN(new_n801));
  OAI21_X1  g600(.A(G120gat), .B1(new_n801), .B2(new_n618), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n617), .A2(new_n335), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n798), .B2(new_n803), .ZN(G1341gat));
  AND3_X1   g603(.A1(new_n792), .A2(G127gat), .A3(new_n658), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n798), .A2(KEYINPUT121), .A3(new_n566), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(G127gat), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT121), .B1(new_n798), .B2(new_n566), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(G1342gat));
  NAND4_X1  g608(.A1(new_n797), .A2(new_n326), .A3(new_n626), .A4(new_n595), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n810), .A2(KEYINPUT56), .ZN(new_n811));
  OAI21_X1  g610(.A(G134gat), .B1(new_n801), .B2(new_n785), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(KEYINPUT56), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(G1343gat));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n636), .A2(new_n486), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n796), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n711), .ZN(new_n818));
  INV_X1    g617(.A(G141gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n819), .A3(new_n259), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n815), .B1(new_n820), .B2(KEYINPUT123), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT57), .B1(new_n787), .B2(new_n420), .ZN(new_n822));
  INV_X1    g621(.A(new_n781), .ZN(new_n823));
  INV_X1    g622(.A(new_n783), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n259), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n595), .B1(new_n825), .B2(new_n782), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n784), .A2(new_n827), .A3(new_n785), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n566), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n763), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n420), .A2(KEYINPUT57), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n822), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n637), .A2(new_n789), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n833), .A2(new_n662), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n820), .B1(new_n835), .B2(new_n819), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n836), .ZN(new_n837));
  OAI221_X1 g636(.A(new_n820), .B1(KEYINPUT123), .B2(new_n815), .C1(new_n835), .C2(new_n819), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1344gat));
  INV_X1    g638(.A(G148gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n818), .A2(new_n840), .A3(new_n617), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n787), .A2(KEYINPUT57), .A3(new_n420), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n617), .B1(new_n843), .B2(new_n822), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n834), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n840), .B1(new_n845), .B2(KEYINPUT124), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n844), .B2(new_n834), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n842), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n833), .A2(new_n618), .A3(new_n834), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(KEYINPUT59), .A3(new_n840), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n841), .B1(new_n849), .B2(new_n851), .ZN(G1345gat));
  NAND3_X1  g651(.A1(new_n818), .A2(new_n383), .A3(new_n658), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n833), .A2(new_n566), .A3(new_n834), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n383), .ZN(G1346gat));
  NAND3_X1  g654(.A1(new_n626), .A2(new_n384), .A3(new_n595), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n817), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n833), .A2(new_n785), .A3(new_n834), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n384), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT125), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n861), .B(new_n857), .C1(new_n858), .C2(new_n384), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1347gat));
  NOR3_X1   g662(.A1(new_n795), .A2(new_n488), .A3(new_n710), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n421), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(G169gat), .B1(new_n866), .B2(new_n259), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n626), .A2(new_n488), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n790), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n788), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n259), .A2(G169gat), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(G1348gat));
  INV_X1    g671(.A(new_n870), .ZN(new_n873));
  OAI21_X1  g672(.A(G176gat), .B1(new_n873), .B2(new_n618), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n618), .A2(G176gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n865), .B2(new_n875), .ZN(G1349gat));
  OR3_X1    g675(.A1(new_n865), .A2(new_n304), .A3(new_n566), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n873), .A2(new_n566), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n269), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT60), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT60), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n877), .B(new_n881), .C1(new_n878), .C2(new_n269), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1350gat));
  AOI21_X1  g682(.A(new_n270), .B1(new_n870), .B2(new_n595), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT61), .Z(new_n885));
  NAND3_X1  g684(.A1(new_n866), .A2(new_n274), .A3(new_n595), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1351gat));
  NAND2_X1  g686(.A1(new_n864), .A2(new_n816), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(G197gat), .B1(new_n889), .B2(new_n259), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n843), .A2(new_n822), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n637), .A2(new_n868), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n892), .A2(KEYINPUT126), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(KEYINPUT126), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n259), .A2(G197gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(G1352gat));
  NOR3_X1   g696(.A1(new_n888), .A2(G204gat), .A3(new_n618), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT62), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n844), .B1(new_n893), .B2(new_n894), .ZN(new_n900));
  INV_X1    g699(.A(G204gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(G1353gat));
  NAND3_X1  g701(.A1(new_n889), .A2(new_n395), .A3(new_n658), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(KEYINPUT127), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n895), .A2(new_n658), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n395), .B1(KEYINPUT127), .B2(new_n904), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n905), .ZN(new_n909));
  INV_X1    g708(.A(new_n907), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n909), .B(new_n910), .C1(new_n895), .C2(new_n658), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n903), .B1(new_n908), .B2(new_n911), .ZN(G1354gat));
  NAND3_X1  g711(.A1(new_n889), .A2(new_n396), .A3(new_n595), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n895), .A2(new_n595), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n396), .ZN(G1355gat));
endmodule


