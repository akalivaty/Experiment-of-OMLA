

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U322 ( .A(n332), .B(KEYINPUT92), .ZN(n539) );
  AND2_X1 U323 ( .A1(n557), .A2(n553), .ZN(n330) );
  XOR2_X1 U324 ( .A(n295), .B(KEYINPUT81), .Z(n290) );
  XOR2_X1 U325 ( .A(n425), .B(n350), .Z(n291) );
  OR2_X1 U326 ( .A1(n539), .A2(n460), .ZN(n456) );
  XNOR2_X1 U327 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n416) );
  XNOR2_X1 U328 ( .A(n417), .B(n416), .ZN(n422) );
  XNOR2_X1 U329 ( .A(KEYINPUT80), .B(KEYINPUT18), .ZN(n294) );
  INV_X1 U330 ( .A(KEYINPUT77), .ZN(n352) );
  XNOR2_X1 U331 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U332 ( .A(n355), .B(n354), .ZN(n361) );
  INV_X1 U333 ( .A(KEYINPUT59), .ZN(n446) );
  XNOR2_X1 U334 ( .A(n488), .B(n487), .ZN(n495) );
  XNOR2_X1 U335 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U336 ( .A(n449), .B(n448), .ZN(G1352GAT) );
  XNOR2_X1 U337 ( .A(KEYINPUT93), .B(KEYINPUT26), .ZN(n331) );
  XOR2_X1 U338 ( .A(KEYINPUT79), .B(G176GAT), .Z(n293) );
  XNOR2_X1 U339 ( .A(G71GAT), .B(G183GAT), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n309) );
  XNOR2_X1 U341 ( .A(n294), .B(G169GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n290), .B(n296), .ZN(n345) );
  XNOR2_X1 U344 ( .A(G127GAT), .B(n345), .ZN(n307) );
  XOR2_X1 U345 ( .A(G15GAT), .B(G190GAT), .Z(n298) );
  XNOR2_X1 U346 ( .A(G120GAT), .B(G99GAT), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U348 ( .A(n299), .B(G43GAT), .Z(n301) );
  XOR2_X1 U349 ( .A(KEYINPUT0), .B(G113GAT), .Z(n428) );
  XNOR2_X1 U350 ( .A(G134GAT), .B(n428), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U352 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n303) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XOR2_X1 U354 ( .A(n303), .B(n302), .Z(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X2 U357 ( .A(n309), .B(n308), .Z(n557) );
  XOR2_X1 U358 ( .A(KEYINPUT85), .B(G197GAT), .Z(n311) );
  XNOR2_X1 U359 ( .A(G218GAT), .B(KEYINPUT84), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U361 ( .A(KEYINPUT21), .B(n312), .Z(n341) );
  XOR2_X1 U362 ( .A(KEYINPUT23), .B(KEYINPUT83), .Z(n314) );
  XNOR2_X1 U363 ( .A(G106GAT), .B(G211GAT), .ZN(n313) );
  XNOR2_X1 U364 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U365 ( .A(G204GAT), .B(G22GAT), .Z(n316) );
  XNOR2_X1 U366 ( .A(G155GAT), .B(G148GAT), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U368 ( .A(n318), .B(n317), .Z(n328) );
  XOR2_X1 U369 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n320) );
  XNOR2_X1 U370 ( .A(G78GAT), .B(KEYINPUT22), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n326) );
  XOR2_X1 U372 ( .A(G162GAT), .B(G50GAT), .Z(n371) );
  XOR2_X1 U373 ( .A(G141GAT), .B(KEYINPUT2), .Z(n322) );
  XNOR2_X1 U374 ( .A(KEYINPUT3), .B(KEYINPUT86), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n426) );
  XOR2_X1 U376 ( .A(n371), .B(n426), .Z(n324) );
  NAND2_X1 U377 ( .A1(G228GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n341), .B(n329), .ZN(n553) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U383 ( .A(G190GAT), .B(G36GAT), .Z(n376) );
  XOR2_X1 U384 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n334) );
  XNOR2_X1 U385 ( .A(G92GAT), .B(G64GAT), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U387 ( .A(n376), .B(n335), .Z(n337) );
  NAND2_X1 U388 ( .A1(G226GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n339) );
  XNOR2_X1 U390 ( .A(G176GAT), .B(G204GAT), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n338), .B(KEYINPUT74), .ZN(n401) );
  XOR2_X1 U392 ( .A(n339), .B(n401), .Z(n343) );
  XNOR2_X1 U393 ( .A(G211GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U394 ( .A(n340), .B(G8GAT), .ZN(n350) );
  XNOR2_X1 U395 ( .A(n350), .B(n341), .ZN(n342) );
  XOR2_X1 U396 ( .A(n343), .B(n342), .Z(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n514) );
  XOR2_X1 U398 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n347) );
  NAND2_X1 U399 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U401 ( .A(n348), .B(KEYINPUT14), .Z(n351) );
  XNOR2_X1 U402 ( .A(G155GAT), .B(G127GAT), .ZN(n349) );
  XOR2_X1 U403 ( .A(n349), .B(G1GAT), .Z(n425) );
  XNOR2_X1 U404 ( .A(n351), .B(n291), .ZN(n355) );
  XOR2_X1 U405 ( .A(G22GAT), .B(G15GAT), .Z(n384) );
  XNOR2_X1 U406 ( .A(n384), .B(KEYINPUT78), .ZN(n353) );
  XNOR2_X1 U407 ( .A(KEYINPUT71), .B(G78GAT), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n356), .B(G71GAT), .ZN(n357) );
  XOR2_X1 U409 ( .A(n357), .B(G64GAT), .Z(n359) );
  XNOR2_X1 U410 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n359), .B(n358), .ZN(n408) );
  INV_X1 U412 ( .A(n408), .ZN(n360) );
  XOR2_X1 U413 ( .A(n361), .B(n360), .Z(n578) );
  INV_X1 U414 ( .A(n578), .ZN(n479) );
  XOR2_X1 U415 ( .A(n479), .B(KEYINPUT111), .Z(n567) );
  XNOR2_X1 U416 ( .A(G99GAT), .B(G106GAT), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n362), .B(KEYINPUT73), .ZN(n363) );
  XOR2_X1 U418 ( .A(n363), .B(KEYINPUT72), .Z(n365) );
  XNOR2_X1 U419 ( .A(G85GAT), .B(G92GAT), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n409) );
  XOR2_X1 U421 ( .A(KEYINPUT10), .B(KEYINPUT64), .Z(n367) );
  XNOR2_X1 U422 ( .A(KEYINPUT11), .B(KEYINPUT76), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n409), .B(n368), .ZN(n381) );
  XOR2_X1 U425 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n370) );
  XNOR2_X1 U426 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n372) );
  XOR2_X1 U428 ( .A(n372), .B(n371), .Z(n379) );
  XNOR2_X1 U429 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n373), .B(KEYINPUT7), .ZN(n388) );
  XOR2_X1 U431 ( .A(G29GAT), .B(G134GAT), .Z(n431) );
  XOR2_X1 U432 ( .A(n388), .B(n431), .Z(n375) );
  NAND2_X1 U433 ( .A1(G232GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n569) );
  XOR2_X1 U438 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n413) );
  XOR2_X1 U439 ( .A(G197GAT), .B(G50GAT), .Z(n383) );
  XNOR2_X1 U440 ( .A(G141GAT), .B(G113GAT), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U442 ( .A(n385), .B(n384), .Z(n387) );
  XNOR2_X1 U443 ( .A(G29GAT), .B(G36GAT), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n392) );
  XOR2_X1 U445 ( .A(n388), .B(KEYINPUT67), .Z(n390) );
  NAND2_X1 U446 ( .A1(G229GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U448 ( .A(n392), .B(n391), .Z(n400) );
  XOR2_X1 U449 ( .A(KEYINPUT70), .B(G169GAT), .Z(n394) );
  XNOR2_X1 U450 ( .A(G1GAT), .B(G8GAT), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U452 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n396) );
  XNOR2_X1 U453 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n558) );
  XOR2_X1 U457 ( .A(G148GAT), .B(G120GAT), .Z(n427) );
  XOR2_X1 U458 ( .A(n401), .B(n427), .Z(n403) );
  NAND2_X1 U459 ( .A1(G230GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U461 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n405) );
  XNOR2_X1 U462 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U464 ( .A(n407), .B(n406), .Z(n411) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n574) );
  XNOR2_X1 U467 ( .A(n574), .B(KEYINPUT41), .ZN(n542) );
  NAND2_X1 U468 ( .A1(n558), .A2(n542), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n414) );
  NOR2_X1 U470 ( .A1(n569), .A2(n414), .ZN(n415) );
  NAND2_X1 U471 ( .A1(n567), .A2(n415), .ZN(n417) );
  XNOR2_X1 U472 ( .A(KEYINPUT36), .B(n569), .ZN(n582) );
  NAND2_X1 U473 ( .A1(n582), .A2(n578), .ZN(n418) );
  XOR2_X1 U474 ( .A(KEYINPUT45), .B(n418), .Z(n419) );
  NAND2_X1 U475 ( .A1(n574), .A2(n419), .ZN(n420) );
  OR2_X1 U476 ( .A1(n558), .A2(n420), .ZN(n421) );
  AND2_X1 U477 ( .A1(n422), .A2(n421), .ZN(n423) );
  XNOR2_X1 U478 ( .A(KEYINPUT48), .B(n423), .ZN(n520) );
  NOR2_X1 U479 ( .A1(n514), .A2(n520), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n424), .B(KEYINPUT54), .ZN(n443) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n442) );
  XOR2_X1 U482 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U485 ( .A(n432), .B(n431), .Z(n440) );
  XOR2_X1 U486 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n434) );
  XNOR2_X1 U487 ( .A(G162GAT), .B(G85GAT), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U489 ( .A(KEYINPUT6), .B(KEYINPUT88), .Z(n436) );
  XNOR2_X1 U490 ( .A(KEYINPUT4), .B(G57GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n457) );
  XOR2_X1 U495 ( .A(KEYINPUT89), .B(n457), .Z(n512) );
  NAND2_X1 U496 ( .A1(n443), .A2(n512), .ZN(n552) );
  NOR2_X1 U497 ( .A1(n539), .A2(n552), .ZN(n444) );
  XOR2_X1 U498 ( .A(KEYINPUT125), .B(n444), .Z(n581) );
  NAND2_X1 U499 ( .A1(n581), .A2(n558), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n445), .B(KEYINPUT60), .ZN(n449) );
  XNOR2_X1 U501 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n447) );
  XNOR2_X1 U502 ( .A(KEYINPUT27), .B(n514), .ZN(n460) );
  XNOR2_X1 U503 ( .A(KEYINPUT25), .B(KEYINPUT95), .ZN(n454) );
  OR2_X1 U504 ( .A1(n557), .A2(n514), .ZN(n450) );
  XNOR2_X1 U505 ( .A(KEYINPUT94), .B(n450), .ZN(n452) );
  INV_X1 U506 ( .A(n553), .ZN(n451) );
  NAND2_X1 U507 ( .A1(n452), .A2(n451), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n456), .A2(n455), .ZN(n458) );
  NAND2_X1 U510 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n459), .B(KEYINPUT96), .ZN(n463) );
  NOR2_X1 U512 ( .A1(n512), .A2(n460), .ZN(n522) );
  XOR2_X1 U513 ( .A(KEYINPUT28), .B(n553), .Z(n523) );
  AND2_X1 U514 ( .A1(n557), .A2(n523), .ZN(n461) );
  NAND2_X1 U515 ( .A1(n522), .A2(n461), .ZN(n462) );
  NAND2_X1 U516 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U517 ( .A(KEYINPUT97), .B(n464), .ZN(n481) );
  NOR2_X1 U518 ( .A1(n569), .A2(n479), .ZN(n465) );
  XOR2_X1 U519 ( .A(KEYINPUT16), .B(n465), .Z(n466) );
  NOR2_X1 U520 ( .A1(n481), .A2(n466), .ZN(n467) );
  XOR2_X1 U521 ( .A(KEYINPUT98), .B(n467), .Z(n499) );
  NAND2_X1 U522 ( .A1(n574), .A2(n558), .ZN(n486) );
  OR2_X1 U523 ( .A1(n499), .A2(n486), .ZN(n476) );
  NOR2_X1 U524 ( .A1(n512), .A2(n476), .ZN(n469) );
  XNOR2_X1 U525 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U527 ( .A(G1GAT), .B(n470), .ZN(G1324GAT) );
  NOR2_X1 U528 ( .A1(n514), .A2(n476), .ZN(n471) );
  XOR2_X1 U529 ( .A(KEYINPUT100), .B(n471), .Z(n472) );
  XNOR2_X1 U530 ( .A(G8GAT), .B(n472), .ZN(G1325GAT) );
  NOR2_X1 U531 ( .A1(n557), .A2(n476), .ZN(n474) );
  XNOR2_X1 U532 ( .A(KEYINPUT35), .B(KEYINPUT101), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U534 ( .A(G15GAT), .B(n475), .Z(G1326GAT) );
  NOR2_X1 U535 ( .A1(n523), .A2(n476), .ZN(n477) );
  XOR2_X1 U536 ( .A(KEYINPUT102), .B(n477), .Z(n478) );
  XNOR2_X1 U537 ( .A(G22GAT), .B(n478), .ZN(G1327GAT) );
  INV_X1 U538 ( .A(KEYINPUT38), .ZN(n488) );
  INV_X1 U539 ( .A(KEYINPUT103), .ZN(n485) );
  NAND2_X1 U540 ( .A1(n479), .A2(n582), .ZN(n480) );
  NOR2_X1 U541 ( .A1(n481), .A2(n480), .ZN(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n511) );
  NOR2_X1 U545 ( .A1(n511), .A2(n486), .ZN(n487) );
  NOR2_X1 U546 ( .A1(n512), .A2(n495), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n489), .B(KEYINPUT39), .ZN(n491) );
  XOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT105), .Z(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NOR2_X1 U550 ( .A1(n514), .A2(n495), .ZN(n492) );
  XOR2_X1 U551 ( .A(G36GAT), .B(n492), .Z(G1329GAT) );
  NOR2_X1 U552 ( .A1(n557), .A2(n495), .ZN(n493) );
  XOR2_X1 U553 ( .A(n493), .B(KEYINPUT40), .Z(n494) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NOR2_X1 U555 ( .A1(n495), .A2(n523), .ZN(n496) );
  XOR2_X1 U556 ( .A(G50GAT), .B(n496), .Z(n497) );
  XNOR2_X1 U557 ( .A(KEYINPUT106), .B(n497), .ZN(G1331GAT) );
  INV_X1 U558 ( .A(n558), .ZN(n498) );
  XOR2_X1 U559 ( .A(KEYINPUT107), .B(n542), .Z(n561) );
  NAND2_X1 U560 ( .A1(n498), .A2(n561), .ZN(n510) );
  OR2_X1 U561 ( .A1(n499), .A2(n510), .ZN(n506) );
  NOR2_X1 U562 ( .A1(n512), .A2(n506), .ZN(n501) );
  XNOR2_X1 U563 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U565 ( .A(G57GAT), .B(n502), .Z(G1332GAT) );
  NOR2_X1 U566 ( .A1(n514), .A2(n506), .ZN(n503) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n503), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n557), .A2(n506), .ZN(n505) );
  XNOR2_X1 U569 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(G1334GAT) );
  NOR2_X1 U571 ( .A1(n523), .A2(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(n509), .ZN(G1335GAT) );
  OR2_X1 U575 ( .A1(n511), .A2(n510), .ZN(n517) );
  NOR2_X1 U576 ( .A1(n512), .A2(n517), .ZN(n513) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U578 ( .A1(n514), .A2(n517), .ZN(n515) );
  XOR2_X1 U579 ( .A(G92GAT), .B(n515), .Z(G1337GAT) );
  NOR2_X1 U580 ( .A1(n557), .A2(n517), .ZN(n516) );
  XOR2_X1 U581 ( .A(G99GAT), .B(n516), .Z(G1338GAT) );
  NOR2_X1 U582 ( .A1(n523), .A2(n517), .ZN(n518) );
  XOR2_X1 U583 ( .A(KEYINPUT44), .B(n518), .Z(n519) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  INV_X1 U585 ( .A(n520), .ZN(n521) );
  NAND2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n538) );
  INV_X1 U587 ( .A(n538), .ZN(n524) );
  NAND2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U589 ( .A1(n557), .A2(n525), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n558), .A2(n534), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U593 ( .A1(n534), .A2(n561), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(n529), .ZN(G1341GAT) );
  INV_X1 U596 ( .A(n534), .ZN(n530) );
  NOR2_X1 U597 ( .A1(n567), .A2(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U602 ( .A1(n534), .A2(n569), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n549) );
  AND2_X1 U606 ( .A1(n558), .A2(n549), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1344GAT) );
  NAND2_X1 U609 ( .A1(n542), .A2(n549), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n543), .B(KEYINPUT52), .ZN(n544) );
  XOR2_X1 U611 ( .A(n544), .B(KEYINPUT53), .Z(n546) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  XOR2_X1 U614 ( .A(G155GAT), .B(KEYINPUT119), .Z(n548) );
  NAND2_X1 U615 ( .A1(n549), .A2(n578), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n549), .A2(n569), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(KEYINPUT120), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n551), .ZN(G1347GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n555) );
  NOR2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n570) );
  NAND2_X1 U624 ( .A1(n570), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT122), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n560), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT123), .Z(n563) );
  NAND2_X1 U628 ( .A1(n570), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  INV_X1 U632 ( .A(n570), .ZN(n566) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n572) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G190GAT), .B(n573), .Z(G1351GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U640 ( .A(n574), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U643 ( .A(G211GAT), .B(KEYINPUT127), .Z(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1354GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

