//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969;
  XNOR2_X1  g000(.A(G169gat), .B(G197gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT86), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G113gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT87), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(G141gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n204), .B(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT12), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(G1gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G1gat), .B2(new_n211), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n214), .B(G8gat), .Z(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G29gat), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n217), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT14), .B(G29gat), .ZN(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G50gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(G43gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(G43gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT15), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT88), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n221), .A2(new_n225), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n223), .B(KEYINPUT90), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n224), .B(KEYINPUT89), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n228), .B1(new_n231), .B2(KEYINPUT15), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n216), .B(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT13), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT17), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n227), .A2(new_n238), .A3(new_n232), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n227), .B2(new_n232), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n215), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT91), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n242), .B1(new_n216), .B2(new_n233), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n242), .B(new_n215), .C1(new_n239), .C2(new_n240), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n244), .A2(new_n245), .B1(G229gat), .B2(G233gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n237), .B1(new_n246), .B2(KEYINPUT18), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n233), .A2(KEYINPUT17), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n232), .A3(new_n238), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n216), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n233), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT91), .B1(new_n251), .B2(new_n215), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n245), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(KEYINPUT18), .A3(new_n235), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n210), .B1(new_n247), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n235), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT18), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n259), .A2(new_n209), .A3(new_n254), .A4(new_n237), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT36), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(KEYINPUT68), .A2(KEYINPUT36), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT27), .B(G183gat), .ZN(new_n267));
  INV_X1    g066(.A(G190gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT28), .ZN(new_n270));
  NOR2_X1   g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT26), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n271), .A2(KEYINPUT26), .ZN(new_n274));
  AND2_X1   g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n272), .B(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n275), .B1(KEYINPUT23), .B2(new_n271), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n280), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT64), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n271), .B2(KEYINPUT23), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n279), .A2(KEYINPUT65), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n279), .A2(new_n273), .A3(new_n281), .A4(new_n283), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT25), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(KEYINPUT25), .B2(new_n284), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n279), .A2(new_n281), .A3(new_n283), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n286), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n279), .A2(new_n281), .A3(new_n283), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT25), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n293), .B(new_n273), .C1(KEYINPUT65), .C2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT25), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n278), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299));
  INV_X1    g098(.A(G120gat), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n300), .A2(G113gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(G113gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OR2_X1    g102(.A1(G127gat), .A2(G134gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G127gat), .A2(G134gat), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n304), .A2(new_n305), .B1(KEYINPUT66), .B2(new_n299), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n303), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n298), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G227gat), .ZN(new_n309));
  INV_X1    g108(.A(G233gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n290), .B1(new_n286), .B2(new_n287), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n292), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n277), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n303), .A2(new_n306), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n303), .A2(new_n306), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n308), .A2(new_n311), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT33), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT67), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G15gat), .B(G43gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(G71gat), .B(G99gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(new_n319), .B2(KEYINPUT32), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n319), .A2(KEYINPUT67), .A3(new_n320), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n323), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n311), .B1(new_n308), .B2(new_n318), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT34), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI211_X1 g131(.A(KEYINPUT34), .B(new_n311), .C1(new_n308), .C2(new_n318), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n319), .B(KEYINPUT32), .C1(new_n320), .C2(new_n326), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n329), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n334), .B1(new_n329), .B2(new_n335), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n265), .B(new_n266), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n329), .A2(new_n335), .ZN(new_n339));
  INV_X1    g138(.A(new_n334), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n329), .A2(new_n334), .A3(new_n335), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n341), .A2(new_n263), .A3(new_n264), .A4(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G78gat), .B(G106gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(G22gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT80), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT69), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT22), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n349), .A2(new_n350), .B1(G211gat), .B2(G218gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(new_n349), .B2(new_n350), .ZN(new_n352));
  XNOR2_X1  g151(.A(G197gat), .B(G204gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT70), .ZN(new_n354));
  XNOR2_X1  g153(.A(G211gat), .B(G218gat), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n352), .B(new_n353), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n354), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT3), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G148gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(G141gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT74), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(G141gat), .ZN(new_n364));
  INV_X1    g163(.A(G141gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G148gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370));
  INV_X1    g169(.A(G155gat), .ZN(new_n371));
  INV_X1    g170(.A(G162gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(new_n373), .B2(KEYINPUT2), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT73), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT2), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n365), .A2(G148gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n377), .B1(new_n362), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n373), .A2(new_n370), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n376), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT2), .B1(new_n366), .B2(new_n364), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n373), .A2(new_n370), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n382), .A2(KEYINPUT73), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n375), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT76), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n379), .A2(new_n376), .A3(new_n380), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT73), .B1(new_n382), .B2(new_n383), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n387), .A2(new_n388), .B1(new_n374), .B2(new_n369), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT76), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n348), .B1(new_n360), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G228gat), .A2(G233gat), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n356), .A2(new_n354), .A3(new_n355), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n355), .A2(new_n354), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n397), .A2(new_n357), .A3(new_n352), .A4(new_n353), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n395), .B1(new_n399), .B2(KEYINPUT29), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n386), .A2(new_n391), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(KEYINPUT80), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n389), .A2(new_n395), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n359), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n399), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n393), .A2(new_n394), .A3(new_n402), .A4(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n405), .B1(new_n360), .B2(new_n389), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(G228gat), .A3(G233gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT31), .B(G50gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n406), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(new_n406), .B2(new_n408), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n347), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n406), .A2(new_n408), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n409), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n406), .A2(new_n408), .A3(new_n410), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n346), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  XOR2_X1   g218(.A(G57gat), .B(G85gat), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT78), .ZN(new_n421));
  XOR2_X1   g220(.A(G1gat), .B(G29gat), .Z(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT5), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n385), .A2(new_n317), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n389), .A2(new_n307), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n426), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n386), .A2(new_n391), .A3(new_n307), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436));
  INV_X1    g235(.A(new_n428), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n433), .A2(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n307), .B1(new_n385), .B2(KEYINPUT3), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n403), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n430), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n432), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n386), .A2(new_n391), .A3(new_n307), .A4(new_n434), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT4), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n443), .A2(new_n444), .B1(new_n403), .B2(new_n439), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n431), .A2(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI211_X1 g246(.A(new_n419), .B(new_n425), .C1(new_n442), .C2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT83), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n425), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n429), .A2(new_n431), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n435), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n436), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n431), .B1(new_n439), .B2(new_n403), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n444), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n459), .A2(new_n440), .A3(new_n446), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n451), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n442), .A2(new_n425), .A3(new_n447), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n419), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n425), .B1(new_n442), .B2(new_n447), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT6), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n450), .B1(new_n466), .B2(new_n449), .ZN(new_n467));
  NAND2_X1  g266(.A1(G226gat), .A2(G233gat), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n468), .B(KEYINPUT71), .Z(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n470), .B1(new_n298), .B2(new_n359), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n314), .A2(new_n469), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n358), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n469), .B1(new_n314), .B2(KEYINPUT29), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n298), .A2(new_n470), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n399), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G8gat), .B(G36gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(G64gat), .B(G92gat), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n478), .B(new_n479), .Z(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n480), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n474), .A2(new_n399), .A3(new_n475), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n399), .B1(new_n474), .B2(new_n475), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT37), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n473), .B2(new_n476), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n482), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT38), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT38), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(new_n482), .C1(new_n485), .C2(new_n487), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n467), .A2(new_n481), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n482), .A3(new_n476), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT72), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT72), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n473), .A2(new_n495), .A3(new_n482), .A4(new_n476), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n477), .B2(new_n480), .ZN(new_n499));
  AOI211_X1 g298(.A(KEYINPUT30), .B(new_n482), .C1(new_n473), .C2(new_n476), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n502));
  OAI211_X1 g301(.A(KEYINPUT39), .B(new_n502), .C1(new_n445), .C2(new_n430), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n459), .A2(new_n440), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT39), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n431), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n506), .A3(new_n425), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(new_n464), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(KEYINPUT81), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT81), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n503), .A2(new_n506), .A3(new_n512), .A4(new_n425), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT82), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n511), .A2(new_n516), .A3(new_n508), .A4(new_n513), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n501), .A2(new_n510), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n418), .B1(new_n492), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT84), .B1(new_n467), .B2(new_n501), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n336), .A2(new_n337), .A3(new_n418), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n465), .A2(KEYINPUT83), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n442), .A2(new_n447), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT6), .B1(new_n523), .B2(new_n451), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n448), .B1(new_n524), .B2(new_n462), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n522), .B1(new_n525), .B2(KEYINPUT83), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT84), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n483), .A2(new_n484), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT30), .B1(new_n528), .B2(new_n482), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n477), .A2(new_n498), .A3(new_n480), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n529), .A2(new_n530), .B1(new_n494), .B2(new_n496), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n526), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n520), .A2(new_n521), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT35), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n344), .A2(new_n519), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n338), .A2(new_n343), .A3(new_n418), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT79), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(new_n501), .B2(new_n525), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n531), .A2(KEYINPUT79), .A3(new_n466), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n262), .B1(new_n535), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n546));
  INV_X1    g345(.A(G57gat), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n546), .B(G64gat), .C1(new_n547), .C2(KEYINPUT93), .ZN(new_n548));
  INV_X1    g347(.A(G64gat), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT92), .B1(new_n549), .B2(G57gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(new_n549), .A3(G57gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  OR2_X1    g353(.A1(G71gat), .A2(G78gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT9), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n554), .B(new_n555), .C1(new_n559), .C2(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT94), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT94), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n215), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(KEYINPUT97), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(KEYINPUT97), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G127gat), .B(G155gat), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT96), .ZN(new_n572));
  NAND2_X1  g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n573), .B(KEYINPUT95), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n572), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n568), .A2(new_n569), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n565), .A2(KEYINPUT21), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n581));
  AND2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  XOR2_X1   g382(.A(G183gat), .B(G211gat), .Z(new_n584));
  OR3_X1    g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n582), .B2(new_n583), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n579), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n576), .A2(new_n585), .A3(new_n586), .A4(new_n578), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT99), .ZN(new_n593));
  NAND2_X1  g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n596), .A2(KEYINPUT100), .A3(KEYINPUT7), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT100), .B1(new_n596), .B2(KEYINPUT7), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n592), .A2(KEYINPUT99), .B1(G85gat), .B2(G92gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(new_n592), .B2(KEYINPUT99), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n596), .A2(KEYINPUT100), .A3(KEYINPUT7), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G99gat), .A2(G106gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT8), .ZN(new_n606));
  OR2_X1    g405(.A1(G85gat), .A2(G92gat), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n606), .A2(KEYINPUT101), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT101), .B1(new_n606), .B2(new_n607), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n599), .B(new_n604), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(G99gat), .A2(G106gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT102), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n605), .ZN(new_n614));
  INV_X1    g413(.A(new_n605), .ZN(new_n615));
  OAI21_X1  g414(.A(KEYINPUT102), .B1(new_n615), .B2(new_n611), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n614), .A2(new_n616), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n602), .A2(new_n603), .B1(new_n593), .B2(new_n594), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT101), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n619), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  OAI22_X1  g427(.A1(new_n239), .A2(new_n240), .B1(new_n618), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT98), .Z(new_n631));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n628), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n233), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G190gat), .B(G218gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT103), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n629), .A2(new_n640), .A3(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n631), .A2(new_n632), .ZN(new_n643));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n639), .A2(new_n645), .A3(new_n641), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n591), .A2(KEYINPUT104), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n647), .A2(new_n648), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n651), .B1(new_n652), .B2(new_n590), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n563), .B1(new_n558), .B2(new_n560), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n558), .A2(new_n563), .A3(new_n560), .ZN(new_n655));
  OAI22_X1  g454(.A1(new_n618), .A2(new_n628), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G230gat), .A2(G233gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n610), .A2(new_n617), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n622), .A2(new_n619), .A3(new_n627), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n561), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n656), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n634), .A2(KEYINPUT10), .A3(new_n565), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT10), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n660), .A2(new_n659), .B1(new_n562), .B2(new_n564), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n659), .A2(new_n660), .A3(new_n561), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n656), .A2(new_n661), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(KEYINPUT105), .A3(new_n665), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n664), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n662), .B1(new_n673), .B2(new_n658), .ZN(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n677), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT105), .B1(new_n671), .B2(new_n665), .ZN(new_n681));
  AOI211_X1 g480(.A(new_n669), .B(KEYINPUT10), .C1(new_n656), .C2(new_n661), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n663), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n658), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n673), .A2(KEYINPUT106), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n680), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n650), .A2(new_n653), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n545), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n466), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT107), .B(G1gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1324gat));
  INV_X1    g493(.A(new_n691), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT16), .B(G8gat), .Z(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n501), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G8gat), .B1(new_n691), .B2(new_n531), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  MUX2_X1   g498(.A(new_n697), .B(new_n699), .S(KEYINPUT42), .Z(G1325gat));
  NOR2_X1   g499(.A1(new_n336), .A2(new_n337), .ZN(new_n701));
  AOI21_X1  g500(.A(G15gat), .B1(new_n695), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n344), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G15gat), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT108), .Z(new_n705));
  AOI21_X1  g504(.A(new_n702), .B1(new_n695), .B2(new_n705), .ZN(G1326gat));
  INV_X1    g505(.A(new_n418), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  AOI21_X1  g509(.A(new_n649), .B1(new_n535), .B2(new_n544), .ZN(new_n711));
  INV_X1    g510(.A(new_n688), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n262), .A2(new_n591), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(G29gat), .A3(new_n466), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n492), .A2(new_n518), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n718), .A2(new_n707), .A3(new_n343), .A4(new_n338), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n521), .A2(new_n532), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n527), .B1(new_n526), .B2(new_n531), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n534), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n542), .B1(new_n536), .B2(new_n537), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n652), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n535), .A2(new_n544), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(KEYINPUT44), .A3(new_n652), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n727), .A2(new_n713), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT110), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n727), .A2(new_n732), .A3(new_n729), .A4(new_n713), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n731), .A2(new_n525), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n717), .B1(new_n734), .B2(new_n217), .ZN(G1328gat));
  NOR3_X1   g534(.A1(new_n714), .A2(G36gat), .A3(new_n531), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT46), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n731), .A2(new_n501), .A3(new_n733), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(new_n220), .ZN(G1329gat));
  INV_X1    g538(.A(new_n701), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n714), .A2(G43gat), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n727), .A2(new_n703), .A3(new_n729), .A4(new_n713), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G43gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n743), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n731), .A2(new_n703), .A3(new_n733), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n741), .B1(new_n750), .B2(G43gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n751), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g551(.A(G50gat), .B1(new_n730), .B2(new_n707), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n712), .A2(new_n591), .A3(new_n649), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n418), .A2(new_n222), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT112), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n545), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n731), .A2(new_n418), .A3(new_n733), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n757), .B1(new_n761), .B2(G50gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n762), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g562(.A1(new_n650), .A2(new_n653), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n764), .A2(new_n262), .A3(new_n712), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n728), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n466), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(new_n547), .ZN(G1332gat));
  NOR2_X1   g567(.A1(new_n766), .A2(new_n531), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  AND2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(G1333gat));
  NOR3_X1   g572(.A1(new_n766), .A2(G71gat), .A3(new_n740), .ZN(new_n774));
  INV_X1    g573(.A(new_n766), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n703), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n774), .B1(G71gat), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n418), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g579(.A1(new_n261), .A2(new_n591), .A3(new_n688), .ZN(new_n781));
  AND4_X1   g580(.A1(new_n525), .A2(new_n727), .A3(new_n729), .A4(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(G85gat), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n261), .A2(new_n591), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n728), .A2(new_n652), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT51), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n711), .A2(new_n787), .A3(new_n784), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n712), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n525), .A2(new_n783), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n782), .A2(new_n783), .B1(new_n789), .B2(new_n790), .ZN(G1336gat));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n531), .A2(G92gat), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n786), .A2(new_n712), .A3(new_n788), .A4(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n727), .A2(new_n501), .A3(new_n729), .A4(new_n781), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n795), .A2(KEYINPUT114), .ZN(new_n796));
  OAI21_X1  g595(.A(G92gat), .B1(new_n795), .B2(KEYINPUT114), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n792), .B(new_n794), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n795), .A2(G92gat), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n688), .B1(new_n785), .B2(KEYINPUT51), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n802), .A2(KEYINPUT113), .A3(new_n788), .A4(new_n793), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n798), .B1(new_n804), .B2(new_n792), .ZN(G1337gat));
  NAND4_X1  g604(.A1(new_n727), .A2(new_n703), .A3(new_n729), .A4(new_n781), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g607(.A(KEYINPUT116), .B(G99gat), .Z(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n806), .A2(new_n807), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n740), .A2(new_n809), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n810), .A2(new_n811), .B1(new_n789), .B2(new_n812), .ZN(G1338gat));
  INV_X1    g612(.A(G106gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n789), .B2(new_n707), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n707), .A2(new_n814), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n727), .A2(new_n729), .A3(new_n781), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(KEYINPUT53), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1339gat));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n683), .A2(new_n823), .A3(new_n657), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n678), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n685), .A2(new_n686), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n823), .B1(new_n673), .B2(new_n658), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n687), .B1(new_n828), .B2(KEYINPUT55), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n658), .B(new_n663), .C1(new_n681), .C2(new_n682), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT54), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n685), .B2(new_n686), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n830), .B1(new_n833), .B2(new_n825), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n829), .A2(new_n261), .A3(new_n834), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n253), .A2(new_n235), .B1(new_n234), .B2(new_n236), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n208), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n260), .A2(new_n837), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n838), .A2(new_n688), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n652), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n260), .A2(new_n842), .A3(new_n837), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n652), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n834), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n590), .B1(new_n840), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n764), .A2(new_n262), .A3(KEYINPUT117), .A4(new_n688), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n689), .B2(new_n261), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n521), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n466), .A3(new_n501), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n261), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n712), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g657(.A1(new_n854), .A2(new_n591), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(G127gat), .ZN(G1342gat));
  INV_X1    g659(.A(new_n853), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n525), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n531), .A2(new_n652), .ZN(new_n863));
  OAI21_X1  g662(.A(G134gat), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(G134gat), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n861), .A2(new_n525), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(KEYINPUT119), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(KEYINPUT119), .ZN(new_n869));
  OAI221_X1 g668(.A(new_n864), .B1(KEYINPUT56), .B2(new_n866), .C1(new_n868), .C2(new_n869), .ZN(G1343gat));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n852), .A2(new_n871), .A3(new_n418), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n703), .A2(new_n466), .A3(new_n501), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT120), .B1(new_n833), .B2(new_n825), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n657), .B1(new_n673), .B2(KEYINPUT106), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n683), .A2(new_n684), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n827), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n824), .A2(new_n678), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n875), .A2(new_n830), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(KEYINPUT121), .A3(new_n829), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n261), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT121), .B1(new_n882), .B2(new_n829), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n839), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n846), .B1(new_n886), .B2(new_n649), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n851), .B1(new_n887), .B2(new_n591), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n418), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n874), .B1(new_n889), .B2(KEYINPUT57), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n365), .B1(new_n890), .B2(new_n261), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n852), .A2(new_n525), .A3(new_n418), .A4(new_n344), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n501), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n365), .A3(new_n261), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT58), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n871), .B1(new_n888), .B2(new_n418), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(new_n262), .A3(new_n874), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n897), .B(new_n894), .C1(new_n899), .C2(new_n365), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n896), .A2(new_n900), .ZN(G1344gat));
  NAND3_X1  g700(.A1(new_n893), .A2(new_n361), .A3(new_n712), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT122), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT59), .B(new_n361), .C1(new_n890), .C2(new_n712), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n707), .A2(KEYINPUT57), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n887), .A2(new_n591), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n689), .A2(new_n261), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n852), .A2(new_n418), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT57), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n909), .A2(new_n712), .A3(new_n873), .A4(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n905), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n903), .B1(new_n904), .B2(new_n913), .ZN(G1345gat));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n915), .B1(new_n893), .B2(new_n591), .ZN(new_n916));
  NOR4_X1   g715(.A1(new_n892), .A2(KEYINPUT123), .A3(new_n501), .A4(new_n590), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n916), .A2(G155gat), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n590), .A2(new_n371), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n890), .B2(new_n919), .ZN(G1346gat));
  OR3_X1    g719(.A1(new_n892), .A2(G162gat), .A3(new_n863), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n898), .A2(new_n649), .A3(new_n874), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n372), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n531), .A2(new_n525), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n853), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n261), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n712), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n591), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n931), .A2(G183gat), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n932));
  OR2_X1    g731(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n926), .A2(new_n267), .A3(new_n591), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(G1350gat));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n926), .A2(new_n652), .B1(new_n938), .B2(new_n268), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(new_n268), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(G1351gat));
  AOI211_X1 g740(.A(new_n536), .B(new_n925), .C1(new_n847), .C2(new_n851), .ZN(new_n942));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n261), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n703), .A2(new_n925), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n909), .A2(new_n911), .A3(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n261), .A2(G197gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  OAI21_X1  g747(.A(G204gat), .B1(new_n945), .B2(new_n688), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n688), .A2(G204gat), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n942), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n949), .A2(new_n953), .A3(new_n954), .ZN(G1353gat));
  INV_X1    g754(.A(G211gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n942), .A2(new_n956), .A3(new_n591), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n909), .A2(new_n591), .A3(new_n911), .A4(new_n944), .ZN(new_n958));
  AND4_X1   g757(.A1(KEYINPUT125), .A2(new_n958), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI22_X1  g760(.A1(new_n958), .A2(new_n961), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n957), .B1(new_n959), .B2(new_n962), .ZN(G1354gat));
  AOI21_X1  g762(.A(G218gat), .B1(new_n942), .B2(new_n652), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n652), .A2(G218gat), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n946), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(G1355gat));
endmodule


