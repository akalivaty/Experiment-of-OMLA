//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1198, new_n1199, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1253, new_n1254, new_n1255;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n203), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT65), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n214), .A2(G1), .A3(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n211), .A2(G20), .A3(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(KEYINPUT66), .B(G238), .Z(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G107), .A2(G264), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n209), .B(new_n217), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT67), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n232), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  XNOR2_X1  g0045(.A(KEYINPUT8), .B(G58), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G20), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT68), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT68), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(new_n248), .A3(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n247), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n253), .B(new_n254), .C1(new_n255), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n213), .A2(new_n215), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n258), .A2(new_n260), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n213), .A2(new_n215), .A3(new_n263), .A4(new_n259), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT69), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT69), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n266), .A2(new_n269), .B1(new_n262), .B2(G20), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n270), .A3(G50), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(G222), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(G223), .A3(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n275), .B(new_n276), .C1(new_n277), .C2(new_n273), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n213), .A2(new_n215), .B1(G33), .B2(G41), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G1), .A3(G13), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n285), .A3(G274), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n287), .B1(G226), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n280), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n280), .A2(new_n294), .A3(new_n290), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n272), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n272), .B(KEYINPUT9), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(G200), .B2(new_n291), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n297), .A2(new_n303), .A3(new_n300), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n296), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT16), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT7), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n273), .A2(new_n307), .A3(G20), .ZN(new_n308));
  INV_X1    g0108(.A(G33), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT3), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT7), .B1(new_n313), .B2(new_n248), .ZN(new_n314));
  OAI21_X1  g0114(.A(G68), .B1(new_n308), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G58), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(new_n219), .ZN(new_n317));
  OAI21_X1  g0117(.A(G20), .B1(new_n317), .B2(new_n202), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n256), .A2(G159), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n306), .B1(new_n315), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n307), .B1(new_n273), .B2(G20), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n311), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n309), .A2(KEYINPUT3), .ZN(new_n325));
  OAI211_X1 g0125(.A(KEYINPUT7), .B(new_n248), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n219), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n327), .A2(KEYINPUT16), .A3(new_n320), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n260), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n268), .A2(new_n270), .A3(new_n247), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n246), .A2(new_n264), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n310), .A2(new_n312), .A3(G226), .A4(G1698), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n310), .A2(new_n312), .A3(G223), .A4(new_n274), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G87), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n279), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n285), .A2(G232), .A3(new_n288), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n286), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT72), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n286), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n292), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(KEYINPUT73), .C1(G179), .C2(new_n345), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT73), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n286), .A2(new_n340), .A3(new_n343), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n343), .B1(new_n286), .B2(new_n340), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(G169), .B1(new_n351), .B2(new_n339), .ZN(new_n352));
  AND4_X1   g0152(.A1(new_n294), .A2(new_n339), .A3(new_n342), .A4(new_n344), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n334), .A2(new_n347), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT18), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT18), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n334), .A2(new_n347), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n315), .A2(new_n306), .A3(new_n321), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT16), .B1(new_n327), .B2(new_n320), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n332), .B1(new_n361), .B2(new_n260), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n339), .A2(new_n342), .A3(new_n298), .A4(new_n344), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT74), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT74), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n351), .A2(new_n365), .A3(new_n298), .A4(new_n339), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n345), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT17), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n362), .A2(new_n369), .A3(KEYINPUT17), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n356), .A2(new_n358), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n250), .A2(G77), .A3(new_n252), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n260), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT11), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n378), .A2(KEYINPUT11), .A3(new_n260), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n219), .B1(new_n262), .B2(G20), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n263), .A2(KEYINPUT12), .A3(G68), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT12), .B1(new_n263), .B2(G68), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n267), .A2(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT14), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G97), .ZN(new_n389));
  OR2_X1    g0189(.A1(G226), .A2(G1698), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n234), .A2(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n389), .B1(new_n392), .B2(new_n313), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n279), .ZN(new_n394));
  INV_X1    g0194(.A(G274), .ZN(new_n395));
  INV_X1    g0195(.A(new_n212), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(new_n284), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n289), .A2(G238), .B1(new_n283), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT13), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n394), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n394), .B2(new_n398), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n388), .B(G169), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n394), .A2(new_n398), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT13), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n394), .A2(new_n398), .A3(new_n399), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(G179), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n405), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n388), .B1(new_n408), .B2(G169), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n387), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(G200), .ZN(new_n411));
  INV_X1    g0211(.A(new_n387), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(new_n412), .C1(new_n298), .C2(new_n408), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n218), .A2(G1698), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n234), .A2(new_n274), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n313), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n279), .B1(G107), .B2(new_n273), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n289), .A2(G244), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n286), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n292), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n420), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n422), .B(new_n294), .C1(new_n416), .C2(new_n417), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n267), .B(G77), .C1(G1), .C2(new_n248), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n246), .A2(new_n257), .B1(new_n248), .B2(new_n277), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT15), .B(G87), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n249), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n260), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n263), .A2(G77), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT70), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n424), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n421), .A2(new_n423), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(G200), .B1(new_n418), .B2(new_n420), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT71), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n422), .B(G190), .C1(new_n416), .C2(new_n417), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n424), .A2(KEYINPUT71), .A3(new_n428), .A4(new_n430), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n433), .A2(new_n435), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  AND4_X1   g0238(.A1(new_n410), .A2(new_n413), .A3(new_n432), .A4(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n305), .A2(new_n375), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT75), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n273), .A2(G250), .A3(G1698), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G283), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT4), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n310), .A2(new_n312), .A3(G244), .A4(new_n274), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n442), .B(new_n443), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n444), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n279), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n262), .B(G45), .C1(new_n281), .C2(KEYINPUT5), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT5), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G41), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n285), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G257), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT79), .B1(new_n451), .B2(G41), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(new_n281), .A3(KEYINPUT5), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n451), .A2(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n282), .A2(G1), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n455), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n285), .A2(G274), .ZN(new_n461));
  OAI22_X1  g0261(.A1(new_n453), .A2(new_n454), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n449), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G179), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n445), .A2(new_n444), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n466), .A2(new_n447), .A3(new_n443), .A4(new_n442), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n462), .B1(new_n467), .B2(new_n279), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G169), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n263), .A2(G97), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n471), .B(KEYINPUT78), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n266), .B1(new_n262), .B2(G33), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n472), .B1(G97), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT6), .ZN(new_n475));
  INV_X1    g0275(.A(G97), .ZN(new_n476));
  INV_X1    g0276(.A(G107), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(KEYINPUT6), .A2(G97), .ZN(new_n481));
  OR3_X1    g0281(.A1(new_n481), .A2(KEYINPUT76), .A3(G107), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT76), .B1(new_n481), .B2(G107), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n485));
  OAI21_X1  g0285(.A(G107), .B1(new_n308), .B2(new_n314), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT77), .B1(new_n487), .B2(new_n260), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT77), .ZN(new_n489));
  INV_X1    g0289(.A(new_n260), .ZN(new_n490));
  AOI211_X1 g0290(.A(new_n489), .B(new_n490), .C1(new_n485), .C2(new_n486), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n474), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n470), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n459), .A2(new_n395), .ZN(new_n494));
  INV_X1    g0294(.A(G250), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n282), .B2(G1), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n285), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n273), .A2(G244), .A3(G1698), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n273), .A2(G238), .A3(new_n274), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G116), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n498), .B1(new_n502), .B2(new_n279), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(G169), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n294), .B2(new_n503), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n273), .A2(new_n248), .A3(G68), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT19), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n248), .B1(new_n389), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n479), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n507), .B1(new_n249), .B2(new_n476), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n490), .B1(new_n513), .B2(KEYINPUT80), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT80), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n506), .A2(new_n515), .A3(new_n511), .A4(new_n512), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n426), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n473), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n426), .A2(new_n264), .ZN(new_n520));
  AND4_X1   g0320(.A1(KEYINPUT81), .A2(new_n517), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n514), .A2(new_n516), .B1(new_n264), .B2(new_n426), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT81), .B1(new_n522), .B2(new_n519), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n505), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n449), .A2(new_n298), .A3(new_n463), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n468), .B2(G200), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(new_n474), .C1(new_n488), .C2(new_n491), .ZN(new_n527));
  INV_X1    g0327(.A(new_n503), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G200), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n473), .A2(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n503), .A2(G190), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n529), .A2(new_n522), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n493), .A2(new_n524), .A3(new_n527), .A4(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n473), .A2(G116), .ZN(new_n535));
  INV_X1    g0335(.A(G116), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n264), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n443), .B(new_n248), .C1(G33), .C2(new_n476), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT83), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(G20), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n260), .A2(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n540), .A2(KEYINPUT20), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT20), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n535), .B(new_n537), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G270), .B(new_n285), .C1(new_n450), .C2(new_n452), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n461), .B2(new_n460), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n310), .A2(new_n312), .A3(G264), .A4(G1698), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n310), .A2(new_n312), .A3(G257), .A4(new_n274), .ZN(new_n549));
  XNOR2_X1  g0349(.A(KEYINPUT82), .B(G303), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n548), .B(new_n549), .C1(new_n273), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n547), .B1(new_n279), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(new_n292), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n545), .A2(KEYINPUT21), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n552), .A2(G179), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n545), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT21), .B1(new_n545), .B2(new_n553), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n264), .A2(new_n477), .ZN(new_n560));
  NOR2_X1   g0360(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n560), .B2(new_n561), .ZN(new_n564));
  AOI22_X1  g0364(.A1(G107), .A2(new_n473), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n273), .A2(new_n248), .A3(G87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT22), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT22), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n273), .A2(new_n569), .A3(new_n248), .A4(G87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n501), .A2(G20), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT23), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n248), .B2(G107), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n477), .A2(KEYINPUT23), .A3(G20), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT24), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT24), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n571), .A2(new_n579), .A3(new_n576), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n566), .B1(new_n581), .B2(new_n260), .ZN(new_n582));
  OAI211_X1 g0382(.A(G264), .B(new_n285), .C1(new_n450), .C2(new_n452), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n310), .A2(new_n312), .A3(G250), .A4(new_n274), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT85), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT85), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n273), .A2(new_n587), .A3(G250), .A4(new_n274), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G294), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n273), .A2(G257), .A3(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n586), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n584), .B1(new_n591), .B2(new_n279), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n460), .A2(new_n461), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n298), .A3(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n595), .B2(G200), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n552), .A2(new_n367), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n545), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n552), .A2(G190), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n582), .A2(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n581), .A2(new_n260), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n565), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n592), .A2(new_n593), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n292), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n595), .A2(new_n294), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n559), .A2(new_n600), .A3(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n441), .A2(new_n534), .A3(new_n607), .ZN(G372));
  NAND2_X1  g0408(.A1(new_n524), .A2(new_n532), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n493), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(KEYINPUT26), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT26), .B1(new_n610), .B2(new_n611), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n524), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n606), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n559), .A2(KEYINPUT86), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n559), .A2(KEYINPUT86), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n582), .A2(new_n596), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n534), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n441), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n356), .A2(new_n358), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n432), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n413), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n628), .A2(new_n410), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n372), .A2(new_n373), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n302), .A2(new_n304), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n296), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n624), .A2(new_n633), .ZN(G369));
  NAND3_X1  g0434(.A1(new_n262), .A2(new_n248), .A3(G13), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n636), .B(KEYINPUT87), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(G213), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(G343), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n602), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n616), .B1(new_n620), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n606), .A2(new_n642), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n545), .A2(new_n642), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n617), .B2(new_n618), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n598), .A2(new_n599), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n559), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT88), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n649), .B1(new_n652), .B2(new_n648), .ZN(new_n653));
  XOR2_X1   g0453(.A(new_n653), .B(KEYINPUT89), .Z(new_n654));
  XNOR2_X1  g0454(.A(KEYINPUT90), .B(G330), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT91), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT91), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n647), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n559), .A2(new_n642), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n646), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n606), .B2(new_n642), .ZN(new_n664));
  XOR2_X1   g0464(.A(new_n664), .B(KEYINPUT92), .Z(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n661), .A2(new_n666), .ZN(G399));
  INV_X1    g0467(.A(KEYINPUT93), .ZN(new_n668));
  INV_X1    g0468(.A(new_n207), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(G41), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n207), .A2(KEYINPUT93), .A3(new_n281), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n510), .A2(G116), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n673), .A2(new_n262), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n211), .B2(new_n673), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT28), .Z(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  INV_X1    g0479(.A(new_n642), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n679), .B(new_n680), .C1(new_n615), .C2(new_n622), .ZN(new_n681));
  INV_X1    g0481(.A(new_n615), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n559), .A2(new_n606), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n534), .A2(new_n683), .A3(new_n620), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n642), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n681), .B1(new_n685), .B2(new_n679), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n592), .A2(new_n552), .A3(G179), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n449), .A2(new_n463), .A3(new_n503), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT94), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g0492(.A(KEYINPUT94), .B(new_n687), .C1(new_n688), .C2(new_n689), .ZN(new_n693));
  INV_X1    g0493(.A(new_n689), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(KEYINPUT30), .A3(new_n555), .A4(new_n592), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n552), .A2(new_n503), .A3(G179), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n464), .A3(new_n603), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n692), .A2(new_n693), .A3(new_n695), .A4(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT31), .B1(new_n698), .B2(new_n642), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n695), .A2(new_n690), .A3(new_n697), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(KEYINPUT31), .A3(new_n642), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n607), .A2(new_n534), .A3(new_n680), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n655), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n686), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n678), .B1(new_n706), .B2(G1), .ZN(G364));
  NAND2_X1  g0507(.A1(new_n658), .A2(new_n659), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n248), .A2(G13), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n262), .B1(new_n709), .B2(G45), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n673), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n654), .B2(new_n656), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT95), .ZN(new_n716));
  INV_X1    g0516(.A(new_n216), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(G20), .B2(new_n292), .ZN(new_n718));
  NOR2_X1   g0518(.A1(G13), .A2(G33), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G20), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n273), .A2(new_n207), .ZN(new_n724));
  INV_X1    g0524(.A(G355), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n724), .A2(new_n725), .B1(G116), .B2(new_n207), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n241), .A2(G45), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n313), .A2(new_n207), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n282), .B2(new_n211), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n248), .A2(new_n294), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G200), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n298), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT96), .Z(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT97), .B(G326), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G190), .A2(G200), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n248), .A2(G179), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n737), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(G311), .A2(new_n739), .B1(new_n742), .B2(G329), .ZN(new_n743));
  INV_X1    g0543(.A(G322), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n731), .A2(G190), .A3(new_n367), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n732), .A2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(G317), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT33), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n748), .A2(KEYINPUT33), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G283), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n740), .A2(new_n298), .A3(G200), .ZN(new_n753));
  INV_X1    g0553(.A(G294), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n298), .A2(G179), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n248), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n751), .B1(new_n752), .B2(new_n753), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n736), .A2(new_n746), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n273), .B1(new_n760), .B2(G303), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT98), .Z(new_n762));
  INV_X1    g0562(.A(new_n733), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT32), .ZN(new_n764));
  INV_X1    g0564(.A(G159), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n741), .A2(new_n765), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n763), .A2(new_n261), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n764), .B2(new_n766), .ZN(new_n768));
  INV_X1    g0568(.A(new_n747), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n769), .A2(new_n219), .B1(new_n753), .B2(new_n477), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n273), .B1(new_n738), .B2(new_n277), .C1(new_n316), .C2(new_n745), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n756), .A2(new_n476), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n759), .A2(new_n509), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n758), .A2(new_n762), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n718), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n712), .B1(new_n723), .B2(new_n730), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT99), .ZN(new_n778));
  INV_X1    g0578(.A(new_n721), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n778), .B1(new_n654), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n716), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  NAND2_X1  g0583(.A1(new_n623), .A2(new_n680), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n642), .A2(new_n431), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n627), .B1(new_n438), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n432), .A2(new_n642), .ZN(new_n787));
  OAI21_X1  g0587(.A(KEYINPUT103), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT103), .ZN(new_n789));
  INV_X1    g0589(.A(new_n787), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n438), .A2(new_n785), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n789), .B(new_n790), .C1(new_n791), .C2(new_n627), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n784), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n793), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n680), .B(new_n795), .C1(new_n615), .C2(new_n622), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n705), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n712), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n794), .A2(new_n705), .A3(new_n796), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n718), .A2(new_n719), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n713), .B1(new_n801), .B2(new_n277), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n753), .A2(new_n509), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n759), .A2(new_n477), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT100), .B(G283), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n803), .B(new_n804), .C1(new_n747), .C2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n273), .B1(new_n739), .B2(G116), .ZN(new_n807));
  INV_X1    g0607(.A(new_n745), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n808), .A2(G294), .B1(new_n742), .B2(G311), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n772), .B1(G303), .B2(new_n733), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n806), .A2(new_n807), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT101), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n273), .B1(new_n741), .B2(new_n813), .C1(new_n261), .C2(new_n759), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n756), .A2(new_n316), .B1(new_n753), .B2(new_n219), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n808), .A2(G143), .B1(new_n739), .B2(G159), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n763), .B2(new_n817), .C1(new_n255), .C2(new_n769), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT34), .Z(new_n819));
  INV_X1    g0619(.A(KEYINPUT102), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n814), .B(new_n815), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n812), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n802), .B1(new_n823), .B2(new_n776), .C1(new_n795), .C2(new_n720), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n800), .A2(new_n824), .ZN(G384));
  NOR3_X1   g0625(.A1(new_n717), .A2(new_n248), .A3(new_n536), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n484), .B(KEYINPUT104), .Z(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT35), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n829), .B2(new_n828), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT36), .ZN(new_n832));
  OR3_X1    g0632(.A1(new_n210), .A2(new_n277), .A3(new_n317), .ZN(new_n833));
  INV_X1    g0633(.A(new_n201), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G68), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n262), .B(G13), .C1(new_n833), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT111), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n686), .A2(new_n441), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n686), .B2(new_n441), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n633), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n640), .B(KEYINPUT107), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n490), .B1(new_n359), .B2(new_n360), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n845), .B2(new_n332), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n370), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n355), .A2(KEYINPUT106), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT106), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n334), .A2(new_n347), .A3(new_n354), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n640), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n334), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n355), .A2(new_n370), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n853), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n374), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT39), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n856), .B2(new_n858), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n851), .A2(new_n855), .B1(new_n374), .B2(new_n857), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT110), .B1(new_n865), .B2(KEYINPUT38), .ZN(new_n866));
  AND4_X1   g0666(.A1(KEYINPUT110), .A2(new_n856), .A3(new_n858), .A4(KEYINPUT38), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n355), .A2(new_n370), .A3(new_n846), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n870));
  INV_X1    g0670(.A(new_n846), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n851), .A2(new_n870), .B1(new_n374), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT109), .B1(new_n872), .B2(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n851), .A2(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n374), .A2(new_n871), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT109), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n860), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n868), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n864), .B1(new_n880), .B2(new_n862), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n410), .A2(new_n642), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n626), .A2(new_n844), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT105), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n387), .A2(new_n886), .A3(new_n642), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n387), .B2(new_n642), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n410), .A2(new_n890), .A3(new_n413), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n410), .B2(new_n413), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n796), .B2(new_n790), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT108), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n861), .B2(new_n863), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n859), .A2(new_n860), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n865), .A2(KEYINPUT38), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT108), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n885), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n884), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n842), .B(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n788), .B(new_n792), .C1(new_n891), .C2(new_n892), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n642), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n699), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n907), .B2(new_n704), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n861), .A2(new_n895), .A3(new_n863), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT108), .B1(new_n897), .B2(new_n898), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(KEYINPUT112), .B(KEYINPUT40), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT113), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n559), .A2(new_n600), .A3(new_n606), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n915), .A2(new_n533), .A3(new_n642), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n916), .A2(new_n699), .A3(new_n906), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n914), .B1(new_n917), .B2(new_n905), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n908), .B2(KEYINPUT113), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n918), .B(new_n920), .C1(new_n868), .C2(new_n879), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n907), .A2(new_n704), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n441), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n655), .B1(new_n922), .B2(new_n924), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n904), .A2(new_n927), .B1(new_n262), .B2(new_n709), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n904), .A2(new_n927), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n837), .B1(new_n928), .B2(new_n929), .ZN(G367));
  INV_X1    g0730(.A(new_n706), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n611), .A2(new_n642), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n492), .A2(new_n642), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n493), .A2(new_n933), .A3(new_n527), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n936));
  NAND3_X1  g0736(.A1(new_n666), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n936), .ZN(new_n938));
  INV_X1    g0738(.A(new_n935), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n938), .B1(new_n665), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n665), .A2(KEYINPUT44), .A3(new_n939), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT44), .B1(new_n665), .B2(new_n939), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n937), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n661), .B(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n658), .A2(new_n659), .A3(new_n647), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n662), .B1(new_n946), .B2(new_n660), .ZN(new_n947));
  INV_X1    g0747(.A(new_n662), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n661), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n931), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n672), .B(KEYINPUT41), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n710), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n935), .B(KEYINPUT114), .Z(new_n954));
  NAND2_X1  g0754(.A1(new_n660), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n663), .A2(new_n939), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT42), .Z(new_n957));
  NAND2_X1  g0757(.A1(new_n954), .A2(new_n616), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n642), .B1(new_n958), .B2(new_n493), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT43), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n680), .B1(new_n522), .B2(new_n530), .ZN(new_n961));
  MUX2_X1   g0761(.A(new_n609), .B(new_n524), .S(new_n961), .Z(new_n962));
  OAI22_X1  g0762(.A1(new_n957), .A2(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n960), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n955), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n962), .A2(new_n721), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n722), .B1(new_n207), .B2(new_n426), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n231), .A2(new_n207), .A3(new_n313), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n712), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n756), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G107), .A2(new_n971), .B1(new_n747), .B2(G294), .ZN(new_n972));
  INV_X1    g0772(.A(G311), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n972), .B1(new_n476), .B2(new_n753), .C1(new_n734), .C2(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n739), .A2(new_n805), .B1(new_n742), .B2(G317), .ZN(new_n975));
  INV_X1    g0775(.A(new_n550), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n273), .B1(new_n808), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n760), .A2(KEYINPUT46), .A3(G116), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT46), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n759), .B2(new_n536), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n975), .A2(new_n977), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n756), .A2(new_n219), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G58), .B2(new_n760), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n313), .B1(new_n808), .B2(G150), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n201), .A2(new_n739), .B1(new_n742), .B2(G137), .ZN(new_n985));
  INV_X1    g0785(.A(new_n753), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n747), .A2(G159), .B1(new_n986), .B2(G77), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n983), .A2(new_n984), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(G143), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n734), .A2(new_n989), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n974), .A2(new_n981), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(KEYINPUT116), .B(KEYINPUT47), .Z(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n970), .B1(new_n993), .B2(new_n718), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n953), .A2(new_n966), .B1(new_n967), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(G387));
  NAND2_X1  g0796(.A1(new_n950), .A2(new_n706), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n947), .A2(new_n949), .A3(new_n931), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n673), .A3(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n724), .A2(new_n674), .B1(G107), .B2(new_n207), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n237), .A2(new_n282), .ZN(new_n1001));
  AOI211_X1 g0801(.A(G45), .B(new_n675), .C1(G68), .C2(G77), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n246), .A2(G50), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT50), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n728), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1000), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n756), .A2(new_n426), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n247), .B2(new_n747), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n277), .B2(new_n759), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G68), .A2(new_n739), .B1(new_n742), .B2(G150), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1010), .B(new_n273), .C1(new_n261), .C2(new_n745), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n763), .A2(new_n765), .B1(new_n753), .B2(new_n476), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n313), .B1(new_n741), .B2(new_n735), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n808), .A2(G317), .B1(new_n739), .B2(new_n976), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n973), .B2(new_n769), .C1(new_n734), .C2(new_n744), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT48), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n971), .A2(new_n805), .B1(new_n760), .B2(G294), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT49), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1014), .B(new_n1023), .C1(G116), .C2(new_n986), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1013), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n712), .B1(new_n723), .B2(new_n1006), .C1(new_n1026), .C2(new_n776), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n647), .B2(new_n721), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT117), .Z(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n950), .B2(new_n711), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n999), .A2(new_n1030), .ZN(G393));
  NAND3_X1  g0831(.A1(new_n944), .A2(new_n950), .A3(new_n706), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n944), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n997), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n673), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n944), .A2(new_n711), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n722), .B1(new_n476), .B2(new_n207), .C1(new_n244), .C2(new_n728), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT118), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(KEYINPUT118), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n712), .A3(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n769), .A2(new_n834), .B1(new_n759), .B2(new_n219), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n273), .B1(new_n741), .B2(new_n989), .C1(new_n246), .C2(new_n738), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n756), .A2(new_n277), .ZN(new_n1043));
  OR4_X1    g0843(.A1(new_n803), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G150), .A2(new_n733), .B1(new_n808), .B2(G159), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G317), .A2(new_n733), .B1(new_n808), .B2(G311), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT52), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n313), .B1(new_n741), .B2(new_n744), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G294), .B2(new_n739), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n971), .A2(G116), .B1(new_n760), .B2(new_n805), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n747), .A2(new_n976), .B1(new_n986), .B2(G107), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1044), .A2(new_n1046), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1040), .B1(new_n718), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n954), .B2(new_n779), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1035), .A2(new_n1036), .A3(new_n1056), .ZN(G390));
  AOI21_X1  g0857(.A(new_n787), .B1(new_n685), .B2(new_n795), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n880), .B(new_n882), .C1(new_n1058), .C2(new_n893), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n894), .A2(new_n883), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n881), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n923), .A2(G330), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1062), .A2(new_n905), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n893), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n705), .A2(new_n795), .A3(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1059), .B(new_n1066), .C1(new_n881), .C2(new_n1060), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n441), .A2(G330), .A3(new_n923), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n633), .B(new_n1069), .C1(new_n839), .C2(new_n840), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n893), .B1(new_n1062), .B2(new_n793), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1058), .A2(new_n1066), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n796), .A2(new_n790), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1065), .B1(new_n705), .B2(new_n795), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1073), .B1(new_n1074), .B2(new_n1063), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1070), .A2(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1068), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1068), .A2(new_n1078), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n673), .A3(new_n1080), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n881), .A2(new_n720), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n801), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n769), .A2(new_n477), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1043), .B(new_n1084), .C1(G283), .C2(new_n733), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G97), .A2(new_n739), .B1(new_n742), .B2(G294), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1086), .B(new_n313), .C1(new_n536), .C2(new_n745), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n773), .B(new_n1087), .C1(G68), .C2(new_n986), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G159), .A2(new_n971), .B1(new_n733), .B2(G128), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n817), .B2(new_n769), .C1(new_n834), .C2(new_n753), .ZN(new_n1090));
  INV_X1    g0890(.A(G125), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n273), .B1(new_n741), .B2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(KEYINPUT54), .B(G143), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n745), .A2(new_n813), .B1(new_n738), .B2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1090), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n759), .A2(new_n255), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT53), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1085), .A2(new_n1088), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n712), .B1(new_n247), .B2(new_n1083), .C1(new_n1098), .C2(new_n776), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT119), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1068), .A2(new_n711), .B1(new_n1082), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1081), .A2(new_n1101), .ZN(G378));
  NAND2_X1  g0902(.A1(new_n272), .A2(new_n852), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n305), .B(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n719), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n712), .B1(new_n1083), .B2(new_n201), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n753), .A2(new_n316), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n763), .A2(new_n536), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(G97), .C2(new_n747), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n273), .A2(G41), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n752), .B2(new_n741), .C1(new_n426), .C2(new_n738), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n982), .B(new_n1113), .C1(G77), .C2(new_n760), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n745), .A2(new_n477), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT120), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1111), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT58), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1112), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1120), .B(new_n261), .C1(G33), .C2(G41), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1091), .A2(new_n763), .B1(new_n769), .B2(new_n813), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n808), .A2(G128), .B1(new_n739), .B2(G137), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n759), .B2(new_n1093), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(G150), .C2(new_n971), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(KEYINPUT59), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n986), .A2(G159), .ZN(new_n1129));
  AOI211_X1 g0929(.A(G33), .B(G41), .C1(new_n742), .C2(G124), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1127), .A2(KEYINPUT59), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1122), .B1(new_n1118), .B2(new_n1117), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1108), .B1(new_n1133), .B2(new_n718), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1107), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n908), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n896), .B2(new_n899), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n912), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n921), .B(G330), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  OR2_X1    g0940(.A1(new_n1140), .A2(new_n1106), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1106), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n1140), .B2(KEYINPUT121), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT121), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n913), .A2(new_n1144), .A3(G330), .A4(new_n921), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1143), .A2(KEYINPUT122), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT122), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1141), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n902), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n884), .B(new_n901), .C1(new_n1140), .C2(new_n1106), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1136), .B1(new_n1153), .B2(new_n711), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1070), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1149), .A2(new_n1152), .B1(new_n1155), .B2(new_n1080), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n673), .B1(new_n1156), .B2(KEYINPUT57), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1152), .A2(KEYINPUT123), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1140), .A2(KEYINPUT121), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n1145), .A3(new_n1106), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT122), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1143), .A2(KEYINPUT122), .A3(new_n1145), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT123), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n1165), .A3(new_n1151), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1158), .A2(new_n1166), .B1(new_n902), .B2(new_n1148), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1080), .A2(new_n1155), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT57), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1154), .B1(new_n1157), .B2(new_n1170), .ZN(G375));
  INV_X1    g0971(.A(new_n1078), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n952), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1070), .A2(new_n1077), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n273), .B1(new_n742), .B2(G303), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n477), .B2(new_n738), .C1(new_n752), .C2(new_n745), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1007), .B(new_n1177), .C1(G77), .C2(new_n986), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n536), .A2(new_n769), .B1(new_n763), .B2(new_n754), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G97), .B2(new_n760), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n756), .A2(new_n261), .B1(new_n759), .B2(new_n765), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G132), .B2(new_n733), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n313), .B1(new_n742), .B2(G128), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n817), .B2(new_n745), .C1(new_n255), .C2(new_n738), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n769), .A2(new_n1093), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1184), .A2(new_n1109), .A3(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1178), .A2(new_n1180), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n712), .B1(G68), .B2(new_n1083), .C1(new_n1187), .C2(new_n776), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n893), .B2(new_n719), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n1076), .B2(new_n711), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1175), .A2(new_n1190), .ZN(G381));
  NOR2_X1   g0991(.A1(G390), .A2(G384), .ZN(new_n1192));
  INV_X1    g0992(.A(G378), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n999), .A2(new_n782), .A3(new_n1030), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(G381), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n995), .A3(new_n1193), .A4(new_n1195), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(G375), .ZN(G407));
  NAND2_X1  g0997(.A1(new_n641), .A2(G213), .ZN(new_n1198));
  OR3_X1    g0998(.A1(G375), .A2(G378), .A3(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(G407), .A2(G213), .A3(new_n1199), .ZN(G409));
  INV_X1    g1000(.A(KEYINPUT125), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1156), .A2(new_n1173), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1165), .B1(new_n1164), .B2(new_n1151), .ZN(new_n1203));
  AOI211_X1 g1003(.A(KEYINPUT123), .B(new_n1150), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1149), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1136), .B1(new_n1205), .B2(new_n711), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT124), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1202), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  AOI211_X1 g1008(.A(KEYINPUT124), .B(new_n1136), .C1(new_n1205), .C2(new_n711), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1201), .B(new_n1193), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1153), .A2(new_n1173), .A3(new_n1168), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1135), .B1(new_n1167), .B2(new_n710), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(KEYINPUT124), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G378), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(G378), .B(new_n1154), .C1(new_n1157), .C2(new_n1170), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT125), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1210), .B(new_n1198), .C1(new_n1215), .C2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT60), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1174), .B1(new_n1078), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n1077), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(new_n673), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1190), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(new_n824), .A3(new_n800), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(G384), .A3(new_n1190), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(KEYINPUT62), .B1(new_n1218), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n641), .A2(G213), .A3(G2897), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1226), .B(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT61), .B1(new_n1218), .B2(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1210), .A2(new_n1198), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT62), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1226), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1193), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(KEYINPUT125), .A3(new_n1216), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .A4(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1227), .A2(new_n1230), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G393), .A2(G396), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G387), .A2(new_n1194), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1194), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n995), .B2(KEYINPUT127), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G390), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1239), .A2(G390), .A3(new_n1241), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1237), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1218), .B2(new_n1226), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1231), .A2(KEYINPUT63), .A3(new_n1233), .A4(new_n1235), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1247), .A2(new_n1249), .A3(new_n1230), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1246), .A2(new_n1251), .ZN(G405));
  NAND2_X1  g1052(.A1(G375), .A2(new_n1193), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1216), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(new_n1226), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1247), .B(new_n1255), .ZN(G402));
endmodule


