//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G113gat), .B(G120gat), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206));
  XNOR2_X1  g005(.A(G127gat), .B(G134gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n205), .B(new_n206), .C1(KEYINPUT70), .C2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G127gat), .B(G134gat), .Z(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(KEYINPUT70), .ZN(new_n210));
  XNOR2_X1  g009(.A(G113gat), .B(G120gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n209), .B(new_n210), .C1(new_n211), .C2(KEYINPUT1), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n215));
  AND2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  OR2_X1    g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(G176gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221));
  INV_X1    g020(.A(G169gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n226), .B1(KEYINPUT65), .B2(new_n235), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n229), .A2(new_n230), .B1(new_n233), .B2(new_n232), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT25), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n234), .A2(new_n227), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n242), .B1(new_n217), .B2(new_n218), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n217), .B2(new_n218), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n246), .A2(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(KEYINPUT67), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n215), .B1(new_n240), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n225), .B(new_n219), .C1(new_n237), .C2(new_n238), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n231), .A2(new_n238), .A3(new_n234), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n242), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n246), .A2(KEYINPUT67), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n246), .A2(KEYINPUT67), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n241), .B(new_n243), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(KEYINPUT68), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT27), .B(G183gat), .Z(new_n259));
  OR2_X1    g058(.A1(new_n259), .A2(G190gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT28), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT69), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n217), .A2(KEYINPUT26), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n245), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n217), .A2(KEYINPUT26), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n261), .A2(KEYINPUT69), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n260), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n263), .A2(new_n267), .A3(new_n233), .A4(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n214), .B1(new_n258), .B2(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n260), .A2(new_n262), .A3(new_n268), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n233), .B1(new_n265), .B2(new_n266), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n260), .A2(new_n262), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AOI211_X1 g074(.A(new_n213), .B(new_n275), .C1(new_n250), .C2(new_n257), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n204), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n253), .A2(KEYINPUT68), .A3(new_n256), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT68), .B1(new_n253), .B2(new_n256), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n270), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n213), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n258), .A2(new_n214), .A3(new_n270), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT71), .A3(new_n204), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G15gat), .B(G43gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(G71gat), .B(G99gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT33), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT71), .B1(new_n285), .B2(new_n204), .ZN(new_n295));
  INV_X1    g094(.A(new_n204), .ZN(new_n296));
  AOI211_X1 g095(.A(new_n278), .B(new_n296), .C1(new_n283), .C2(new_n284), .ZN(new_n297));
  OAI211_X1 g096(.A(KEYINPUT72), .B(new_n294), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT32), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n291), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT72), .B1(new_n287), .B2(new_n294), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n293), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n296), .A3(new_n284), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT34), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(G211gat), .B(G218gat), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n308));
  OR2_X1    g107(.A1(G197gat), .A2(G204gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(G197gat), .A2(G204gat), .ZN(new_n310));
  AOI211_X1 g109(.A(KEYINPUT74), .B(new_n308), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n310), .ZN(new_n313));
  INV_X1    g112(.A(new_n308), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n307), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n312), .A3(new_n314), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n306), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT29), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  OR2_X1    g118(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(G141gat), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G141gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G148gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n322), .A2(new_n324), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n326), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n325), .ZN(new_n331));
  AND2_X1   g130(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n332));
  NOR2_X1   g131(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n325), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n323), .A2(G148gat), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n334), .A2(new_n335), .B1(new_n324), .B2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(KEYINPUT78), .B(new_n325), .C1(new_n332), .C2(new_n333), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n331), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI22_X1  g138(.A1(new_n319), .A2(KEYINPUT3), .B1(new_n329), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n313), .A2(new_n314), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT74), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n306), .B1(new_n342), .B2(new_n317), .ZN(new_n343));
  INV_X1    g142(.A(new_n318), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT75), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n316), .A2(new_n346), .A3(new_n318), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n334), .A2(new_n335), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n336), .A2(new_n324), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n338), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n331), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n329), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT29), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n340), .B1(new_n348), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(new_n348), .B2(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  OAI221_X1 g160(.A(new_n340), .B1(new_n357), .B2(new_n359), .C1(new_n348), .C2(new_n355), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G22gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(G22gat), .A3(new_n362), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT31), .B(G50gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT81), .ZN(new_n368));
  XOR2_X1   g167(.A(G78gat), .B(G106gat), .Z(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  AND4_X1   g169(.A1(KEYINPUT83), .A2(new_n365), .A3(new_n366), .A4(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n373), .A2(new_n370), .B1(new_n365), .B2(new_n366), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT72), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n290), .B1(new_n287), .B2(KEYINPUT32), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n379), .A3(new_n298), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT32), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n279), .B2(new_n286), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n304), .B1(new_n382), .B2(new_n292), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n375), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n305), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT86), .ZN(new_n386));
  XNOR2_X1  g185(.A(G8gat), .B(G36gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT76), .ZN(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  NAND2_X1  g189(.A1(new_n253), .A2(new_n256), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n391), .A2(new_n270), .ZN(new_n392));
  INV_X1    g191(.A(G226gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n203), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n348), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n275), .B1(new_n250), .B2(new_n257), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n394), .A2(KEYINPUT29), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n395), .B(new_n396), .C1(new_n397), .C2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n258), .A2(new_n270), .A3(new_n394), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n391), .A2(new_n270), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n398), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n396), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n390), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n394), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n404), .B1(new_n282), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n348), .ZN(new_n409));
  INV_X1    g208(.A(new_n390), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n400), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n406), .A2(KEYINPUT30), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n409), .A2(new_n413), .A3(new_n400), .A4(new_n410), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n416), .B(KEYINPUT80), .Z(new_n417));
  NOR2_X1   g216(.A1(new_n353), .A2(new_n214), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n339), .A2(new_n213), .A3(new_n329), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT5), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n353), .A2(new_n354), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT3), .B1(new_n339), .B2(new_n329), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n423), .A3(new_n213), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n353), .A2(new_n214), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n417), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n353), .A2(new_n214), .A3(KEYINPUT4), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n424), .A2(new_n427), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n421), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G1gat), .B(G29gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT0), .ZN(new_n433));
  XNOR2_X1  g232(.A(G57gat), .B(G85gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NOR4_X1   g235(.A1(new_n339), .A2(new_n213), .A3(new_n426), .A4(new_n329), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT4), .B1(new_n353), .B2(new_n214), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n439), .A2(KEYINPUT5), .A3(new_n428), .A4(new_n424), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n431), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n436), .B1(new_n431), .B2(new_n440), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT84), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n441), .A2(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n440), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n435), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT84), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n442), .A4(new_n441), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n445), .A2(new_n446), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n386), .B1(new_n415), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n412), .A2(new_n414), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n445), .A2(new_n446), .A3(new_n450), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT86), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT35), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n448), .A2(new_n442), .A3(new_n441), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n446), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n305), .A2(new_n384), .A3(new_n460), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n385), .A2(new_n456), .B1(new_n461), .B2(KEYINPUT35), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n213), .B1(new_n339), .B2(new_n329), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n425), .A2(new_n463), .A3(new_n428), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT39), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n424), .A2(new_n427), .A3(new_n429), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(new_n417), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT39), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(new_n469), .A3(new_n417), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n468), .A2(KEYINPUT40), .A3(new_n435), .A4(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT40), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n435), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(new_n467), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n471), .A2(new_n474), .A3(new_n441), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(new_n412), .A3(new_n414), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n371), .A2(new_n374), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n395), .B(new_n348), .C1(new_n397), .C2(new_n399), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT37), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n397), .A2(new_n394), .B1(new_n398), .B2(new_n403), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(new_n348), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n408), .A2(new_n396), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n485), .A2(KEYINPUT85), .A3(KEYINPUT37), .A4(new_n480), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n400), .B(new_n488), .C1(new_n482), .C2(new_n396), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT38), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n489), .A2(new_n490), .A3(new_n390), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n390), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n488), .B1(new_n409), .B2(new_n400), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT38), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n451), .A2(new_n492), .A3(new_n411), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n459), .A2(new_n375), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g298(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n500));
  INV_X1    g299(.A(new_n304), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(new_n380), .B2(new_n293), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n293), .A2(new_n501), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n298), .A2(new_n299), .A3(new_n291), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(new_n378), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n500), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n380), .A2(new_n383), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n305), .A2(KEYINPUT36), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n499), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n462), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(G57gat), .B(G64gat), .Z(new_n511));
  INV_X1    g310(.A(KEYINPUT9), .ZN(new_n512));
  INV_X1    g311(.A(G71gat), .ZN(new_n513));
  INV_X1    g312(.A(G78gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n511), .A2(KEYINPUT92), .A3(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G71gat), .B(G78gat), .Z(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT93), .ZN(new_n521));
  XOR2_X1   g320(.A(G127gat), .B(G155gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT20), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n521), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G183gat), .B(G211gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT16), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(G1gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(G1gat), .B2(new_n527), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(G8gat), .Z(new_n531));
  INV_X1    g330(.A(KEYINPUT95), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n518), .B(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n533), .B2(new_n519), .ZN(new_n534));
  XOR2_X1   g333(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n535));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n535), .B(new_n536), .Z(new_n537));
  XNOR2_X1  g336(.A(new_n534), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n526), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT87), .B(G29gat), .ZN(new_n540));
  INV_X1    g339(.A(G36gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(G29gat), .A2(G36gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT14), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G43gat), .B(G50gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n545), .B1(KEYINPUT88), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT15), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n546), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n542), .B2(new_n544), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n548), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT7), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT7), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT96), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n557), .A2(new_n559), .A3(G85gat), .A4(G92gat), .ZN(new_n560));
  INV_X1    g359(.A(G85gat), .ZN(new_n561));
  INV_X1    g360(.A(G92gat), .ZN(new_n562));
  OAI211_X1 g361(.A(KEYINPUT96), .B(new_n558), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(KEYINPUT8), .A2(new_n564), .B1(new_n561), .B2(new_n562), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G99gat), .B(G106gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT17), .B1(new_n549), .B2(new_n552), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n572), .B1(new_n553), .B2(new_n568), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G190gat), .B(G218gat), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n577), .A3(new_n573), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n583), .A2(KEYINPUT97), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(KEYINPUT97), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n579), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(new_n579), .B2(new_n585), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n539), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n568), .A2(KEYINPUT10), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT101), .B1(new_n533), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n518), .B(KEYINPUT95), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n591), .A2(new_n592), .A3(KEYINPUT10), .A4(new_n568), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n567), .B1(new_n566), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n595), .B2(new_n566), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n567), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n566), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n518), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n569), .A2(new_n518), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n594), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n603), .A2(new_n604), .ZN(new_n610));
  INV_X1    g409(.A(new_n608), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G120gat), .B(G148gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT102), .ZN(new_n614));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  NAND3_X1  g415(.A1(new_n609), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n611), .B1(new_n594), .B2(new_n606), .ZN(new_n619));
  INV_X1    g418(.A(new_n612), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n588), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G197gat), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT11), .B(G169gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  NAND3_X1  g428(.A1(new_n555), .A2(new_n531), .A3(new_n570), .ZN(new_n630));
  NAND2_X1  g429(.A1(G229gat), .A2(G233gat), .ZN(new_n631));
  OR3_X1    g430(.A1(new_n531), .A2(new_n549), .A3(new_n552), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n553), .B(new_n531), .Z(new_n634));
  XOR2_X1   g433(.A(new_n631), .B(KEYINPUT13), .Z(new_n635));
  AOI22_X1  g434(.A1(new_n633), .A2(KEYINPUT18), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT90), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n639), .A2(KEYINPUT90), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n629), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(KEYINPUT91), .ZN(new_n644));
  INV_X1    g443(.A(new_n629), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT91), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n637), .A2(new_n646), .A3(new_n638), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n636), .A2(new_n644), .A3(new_n645), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n510), .A2(new_n624), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n458), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT103), .B(G1gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n415), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT16), .B(G8gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT42), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(G8gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT104), .Z(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(G1325gat));
  INV_X1    g461(.A(G15gat), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n502), .A2(new_n505), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n651), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT36), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n502), .A2(new_n505), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n500), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n305), .B2(new_n507), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n651), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n665), .B1(new_n671), .B2(new_n663), .ZN(G1326gat));
  NAND2_X1  g471(.A1(new_n651), .A2(new_n375), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  INV_X1    g474(.A(new_n587), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n649), .A2(new_n539), .A3(new_n623), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n510), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n652), .A3(new_n540), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT45), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT105), .B1(new_n462), .B2(new_n509), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n461), .A2(KEYINPUT35), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n456), .A2(new_n305), .A3(new_n384), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n497), .A2(new_n498), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n667), .B2(new_n669), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n676), .A2(KEYINPUT44), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n681), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT44), .B1(new_n510), .B2(new_n676), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n677), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n692), .A2(KEYINPUT106), .A3(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(new_n458), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n680), .B1(new_n699), .B2(new_n540), .ZN(G1328gat));
  OAI21_X1  g499(.A(G36gat), .B1(new_n698), .B2(new_n453), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n678), .A2(new_n541), .A3(new_n415), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT46), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(G1329gat));
  INV_X1    g503(.A(new_n678), .ZN(new_n705));
  NOR4_X1   g504(.A1(new_n705), .A2(G43gat), .A3(new_n505), .A4(new_n502), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n670), .ZN(new_n709));
  OAI21_X1  g508(.A(G43gat), .B1(new_n694), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n670), .A3(new_n697), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n706), .B1(new_n712), .B2(G43gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n713), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g513(.A(G50gat), .B1(new_n694), .B2(new_n477), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n678), .A2(KEYINPUT107), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n477), .A2(G50gat), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n705), .B2(new_n718), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n715), .B(KEYINPUT48), .C1(new_n716), .C2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n716), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n696), .A2(new_n375), .A3(new_n697), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(G50gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n720), .B1(new_n723), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g523(.A1(new_n681), .A2(new_n688), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n649), .A2(new_n539), .A3(new_n587), .A4(new_n623), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n458), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT108), .B(G57gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1332gat));
  AOI21_X1  g529(.A(new_n453), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OR3_X1    g531(.A1(new_n727), .A2(KEYINPUT109), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT109), .B1(new_n727), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1333gat));
  OAI21_X1  g536(.A(G71gat), .B1(new_n727), .B2(new_n709), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n664), .A2(new_n513), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n727), .B2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g540(.A1(new_n727), .A2(new_n477), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(new_n514), .ZN(G1335gat));
  INV_X1    g542(.A(new_n539), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n744), .A2(new_n649), .A3(new_n623), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n692), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n746), .A2(new_n652), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n744), .A2(new_n649), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n587), .B(new_n748), .C1(new_n462), .C2(new_n509), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n684), .A2(new_n686), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n752), .A2(KEYINPUT51), .A3(new_n587), .A4(new_n748), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n622), .A2(new_n561), .A3(new_n652), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n747), .A2(new_n561), .B1(new_n755), .B2(new_n756), .ZN(G1336gat));
  NOR4_X1   g556(.A1(new_n755), .A2(G92gat), .A3(new_n453), .A4(new_n623), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n746), .A2(new_n415), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n759), .B(new_n760), .C1(new_n761), .C2(new_n562), .ZN(new_n762));
  INV_X1    g561(.A(new_n760), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n562), .B1(new_n746), .B2(new_n415), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n758), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(new_n765), .ZN(G1337gat));
  AND2_X1   g565(.A1(new_n746), .A2(new_n670), .ZN(new_n767));
  INV_X1    g566(.A(G99gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n664), .A2(new_n768), .A3(new_n622), .ZN(new_n769));
  OAI22_X1  g568(.A1(new_n767), .A2(new_n768), .B1(new_n755), .B2(new_n769), .ZN(G1338gat));
  NAND3_X1  g569(.A1(new_n692), .A2(new_n375), .A3(new_n745), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n623), .A2(new_n477), .A3(G106gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n751), .B2(new_n753), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT111), .B1(new_n754), .B2(new_n773), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780));
  AOI211_X1 g579(.A(new_n780), .B(new_n774), .C1(new_n751), .C2(new_n753), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n779), .A2(new_n781), .A3(KEYINPUT53), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT112), .B1(new_n782), .B2(new_n772), .ZN(new_n783));
  INV_X1    g582(.A(new_n779), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT53), .B1(new_n775), .B2(KEYINPUT111), .ZN(new_n785));
  AND4_X1   g584(.A1(KEYINPUT112), .A2(new_n772), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n778), .B1(new_n783), .B2(new_n786), .ZN(G1339gat));
  NAND2_X1  g586(.A1(new_n305), .A2(new_n384), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n594), .A2(new_n611), .A3(new_n606), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n609), .A2(KEYINPUT54), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n616), .B1(new_n619), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(KEYINPUT55), .A3(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(new_n617), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n792), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n649), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n634), .A2(new_n635), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n631), .B1(new_n630), .B2(new_n632), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n628), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n648), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n622), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n587), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n587), .A2(new_n797), .A3(new_n617), .A4(new_n793), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n802), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n539), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n624), .A2(new_n649), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n788), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n811), .A2(new_n652), .A3(new_n453), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n649), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n622), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n744), .ZN(new_n817));
  INV_X1    g616(.A(G127gat), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT113), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n817), .B(new_n819), .ZN(G1342gat));
  AOI21_X1  g619(.A(new_n458), .B1(new_n808), .B2(new_n810), .ZN(new_n821));
  INV_X1    g620(.A(G134gat), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n587), .A2(new_n453), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT114), .Z(new_n824));
  NAND4_X1  g623(.A1(new_n821), .A2(new_n822), .A3(new_n385), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT56), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n822), .B1(new_n812), .B2(new_n587), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(new_n827), .ZN(G1343gat));
  NOR3_X1   g627(.A1(new_n670), .A2(new_n458), .A3(new_n415), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n477), .B1(new_n808), .B2(new_n810), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(KEYINPUT57), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  AOI211_X1 g631(.A(new_n832), .B(new_n477), .C1(new_n808), .C2(new_n810), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n829), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G141gat), .B1(new_n834), .B2(new_n650), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n821), .A2(KEYINPUT115), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT115), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n670), .A2(new_n477), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n836), .A2(new_n453), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n649), .A2(new_n323), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT58), .ZN(G1344gat));
  AND2_X1   g641(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n803), .B1(new_n806), .B2(KEYINPUT117), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n643), .A2(new_n648), .B1(new_n796), .B2(new_n795), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n845), .A2(new_n794), .B1(new_n622), .B2(new_n803), .ZN(new_n846));
  OAI22_X1  g645(.A1(new_n843), .A2(new_n844), .B1(new_n846), .B2(new_n587), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n809), .B1(new_n847), .B2(new_n539), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n832), .B1(new_n848), .B2(new_n477), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n830), .A2(KEYINPUT57), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n622), .A4(new_n829), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G148gat), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n623), .B1(new_n849), .B2(new_n850), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n852), .B1(new_n855), .B2(new_n829), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT59), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n622), .B(new_n829), .C1(new_n831), .C2(new_n833), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n320), .A2(new_n321), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT116), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n858), .A2(new_n863), .A3(new_n859), .A4(new_n860), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n857), .A2(new_n865), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n839), .A2(new_n860), .A3(new_n623), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1345gat));
  OAI21_X1  g667(.A(G155gat), .B1(new_n834), .B2(new_n539), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n539), .A2(G155gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n839), .B2(new_n870), .ZN(G1346gat));
  OR2_X1    g670(.A1(new_n834), .A2(new_n676), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G162gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n874));
  INV_X1    g673(.A(G162gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n824), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n874), .B2(new_n876), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n453), .A2(new_n652), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n811), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n650), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(G169gat), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n223), .A2(new_n224), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n880), .ZN(G1348gat));
  INV_X1    g682(.A(new_n879), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n622), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n259), .A3(new_n744), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n879), .A2(new_n539), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(G183gat), .B2(new_n888), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n889), .B(KEYINPUT60), .Z(G1350gat));
  NAND2_X1  g689(.A1(new_n884), .A2(new_n587), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(G190gat), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n892), .A2(KEYINPUT61), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n891), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n891), .A2(G190gat), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(KEYINPUT119), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n895), .A2(KEYINPUT119), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n893), .B(new_n894), .C1(new_n896), .C2(new_n897), .ZN(G1351gat));
  NOR3_X1   g697(.A1(new_n670), .A2(new_n652), .A3(new_n453), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n830), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n830), .A2(KEYINPUT120), .A3(new_n899), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n649), .A3(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(G197gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n899), .B(KEYINPUT121), .Z(new_n907));
  NAND3_X1  g706(.A1(new_n851), .A2(G197gat), .A3(new_n649), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n909), .B(new_n910), .ZN(G1352gat));
  XNOR2_X1  g710(.A(KEYINPUT123), .B(G204gat), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n900), .A2(new_n623), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT62), .ZN(new_n914));
  INV_X1    g713(.A(new_n855), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n915), .B2(new_n907), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1353gat));
  NOR2_X1   g716(.A1(new_n539), .A2(G211gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920));
  OAI21_X1  g719(.A(G211gat), .B1(new_n920), .B2(KEYINPUT63), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n899), .A2(new_n744), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n851), .B2(new_n922), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n923), .A2(new_n920), .A3(KEYINPUT63), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n920), .B2(KEYINPUT63), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(G1354gat));
  NAND3_X1  g725(.A1(new_n902), .A2(new_n587), .A3(new_n903), .ZN(new_n927));
  INV_X1    g726(.A(G218gat), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n587), .A2(G218gat), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT125), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n851), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n907), .B2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n933), .B(new_n934), .ZN(G1355gat));
endmodule


