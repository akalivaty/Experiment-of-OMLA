

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(n626), .A2(n1004), .ZN(n629) );
  AND2_X1 U552 ( .A1(G2104), .A2(G2105), .ZN(n983) );
  BUF_X2 U553 ( .A(n589), .Z(n986) );
  NOR2_X1 U554 ( .A1(n611), .A2(n610), .ZN(n613) );
  XNOR2_X1 U555 ( .A(n660), .B(n659), .ZN(n679) );
  XNOR2_X1 U556 ( .A(n695), .B(n694), .ZN(n696) );
  INV_X1 U557 ( .A(KEYINPUT5), .ZN(n527) );
  INV_X1 U558 ( .A(KEYINPUT23), .ZN(n534) );
  AND2_X1 U559 ( .A1(G138), .A2(n987), .ZN(n594) );
  XOR2_X1 U560 ( .A(n662), .B(KEYINPUT30), .Z(n517) );
  AND2_X1 U561 ( .A1(n591), .A2(n590), .ZN(n518) );
  OR2_X1 U562 ( .A1(n607), .A2(n606), .ZN(n608) );
  INV_X1 U563 ( .A(KEYINPUT96), .ZN(n612) );
  XNOR2_X1 U564 ( .A(n613), .B(n612), .ZN(n626) );
  INV_X1 U565 ( .A(KEYINPUT97), .ZN(n662) );
  XNOR2_X1 U566 ( .A(n663), .B(n517), .ZN(n664) );
  OR2_X1 U567 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U568 ( .A1(n658), .A2(G2084), .ZN(n660) );
  NOR2_X1 U569 ( .A1(G1966), .A2(n706), .ZN(n685) );
  XNOR2_X1 U570 ( .A(KEYINPUT70), .B(KEYINPUT12), .ZN(n615) );
  XNOR2_X1 U571 ( .A(n616), .B(n615), .ZN(n618) );
  INV_X1 U572 ( .A(KEYINPUT101), .ZN(n694) );
  NOR2_X1 U573 ( .A1(G651), .A2(G543), .ZN(n800) );
  INV_X1 U574 ( .A(KEYINPUT17), .ZN(n538) );
  XNOR2_X1 U575 ( .A(n527), .B(KEYINPUT74), .ZN(n528) );
  NOR2_X1 U576 ( .A1(n566), .A2(n524), .ZN(n801) );
  NOR2_X1 U577 ( .A1(G651), .A2(n566), .ZN(n806) );
  XNOR2_X1 U578 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U579 ( .A(n535), .B(n534), .ZN(n537) );
  XNOR2_X1 U580 ( .A(KEYINPUT8), .B(KEYINPUT75), .ZN(n544) );
  XNOR2_X1 U581 ( .A(G168), .B(n544), .ZN(G286) );
  INV_X1 U582 ( .A(G651), .ZN(n524) );
  NOR2_X1 U583 ( .A1(G543), .A2(n524), .ZN(n519) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n519), .Z(n805) );
  NAND2_X1 U585 ( .A1(G63), .A2(n805), .ZN(n521) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n566) );
  NAND2_X1 U587 ( .A1(G51), .A2(n806), .ZN(n520) );
  NAND2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(KEYINPUT6), .B(n522), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n800), .A2(G89), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n523), .B(KEYINPUT4), .ZN(n526) );
  NAND2_X1 U592 ( .A1(G76), .A2(n801), .ZN(n525) );
  NAND2_X1 U593 ( .A1(n526), .A2(n525), .ZN(n529) );
  NOR2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U595 ( .A(KEYINPUT7), .B(n532), .Z(G168) );
  INV_X1 U596 ( .A(G2104), .ZN(n533) );
  NOR2_X2 U597 ( .A1(G2105), .A2(n533), .ZN(n589) );
  NAND2_X1 U598 ( .A1(G101), .A2(n589), .ZN(n535) );
  AND2_X2 U599 ( .A1(n533), .A2(G2105), .ZN(n982) );
  NAND2_X1 U600 ( .A1(n982), .A2(G125), .ZN(n536) );
  NAND2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n543) );
  NOR2_X2 U602 ( .A1(G2104), .A2(G2105), .ZN(n539) );
  XNOR2_X2 U603 ( .A(n539), .B(n538), .ZN(n987) );
  NAND2_X1 U604 ( .A1(n987), .A2(G137), .ZN(n541) );
  NAND2_X1 U605 ( .A1(G113), .A2(n983), .ZN(n540) );
  NAND2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X2 U607 ( .A1(n543), .A2(n542), .ZN(G160) );
  NAND2_X1 U608 ( .A1(G91), .A2(n800), .ZN(n546) );
  NAND2_X1 U609 ( .A1(G78), .A2(n801), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n805), .A2(G65), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT68), .B(n547), .Z(n548) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n806), .A2(G53), .ZN(n550) );
  NAND2_X1 U615 ( .A1(n551), .A2(n550), .ZN(G299) );
  NAND2_X1 U616 ( .A1(G64), .A2(n805), .ZN(n553) );
  NAND2_X1 U617 ( .A1(G52), .A2(n806), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G90), .A2(n800), .ZN(n555) );
  NAND2_X1 U620 ( .A1(G77), .A2(n801), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(G171) );
  NAND2_X1 U624 ( .A1(G50), .A2(n806), .ZN(n560) );
  NAND2_X1 U625 ( .A1(G75), .A2(n801), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G62), .A2(n805), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G88), .A2(n800), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT83), .ZN(G303) );
  NAND2_X1 U632 ( .A1(G87), .A2(n566), .ZN(n568) );
  NAND2_X1 U633 ( .A1(G74), .A2(G651), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U635 ( .A1(n805), .A2(n569), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G49), .A2(n806), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT81), .B(n570), .Z(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(G288) );
  NAND2_X1 U639 ( .A1(G61), .A2(n805), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G86), .A2(n800), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(KEYINPUT82), .B(n575), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n801), .A2(G73), .ZN(n576) );
  XOR2_X1 U644 ( .A(KEYINPUT2), .B(n576), .Z(n577) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n806), .A2(G48), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(G305) );
  NAND2_X1 U648 ( .A1(G60), .A2(n805), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G47), .A2(n806), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U651 ( .A(KEYINPUT67), .B(n583), .Z(n586) );
  NAND2_X1 U652 ( .A1(G85), .A2(n800), .ZN(n584) );
  XOR2_X1 U653 ( .A(KEYINPUT66), .B(n584), .Z(n585) );
  NOR2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n801), .A2(G72), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(G290) );
  NAND2_X1 U657 ( .A1(G160), .A2(G40), .ZN(n714) );
  INV_X1 U658 ( .A(n714), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G102), .A2(n986), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G114), .A2(n983), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G126), .A2(n982), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n592), .A2(n518), .ZN(n593) );
  NOR2_X1 U663 ( .A1(n594), .A2(n593), .ZN(G164) );
  NOR2_X2 U664 ( .A1(G164), .A2(G1384), .ZN(n715) );
  NAND2_X1 U665 ( .A1(n595), .A2(n715), .ZN(n596) );
  XNOR2_X1 U666 ( .A(n596), .B(KEYINPUT64), .ZN(n606) );
  BUF_X2 U667 ( .A(n606), .Z(n658) );
  NAND2_X1 U668 ( .A1(n658), .A2(G8), .ZN(n706) );
  NAND2_X1 U669 ( .A1(G92), .A2(n800), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G66), .A2(n805), .ZN(n598) );
  NAND2_X1 U671 ( .A1(G54), .A2(n806), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U673 ( .A1(G79), .A2(n801), .ZN(n599) );
  XNOR2_X1 U674 ( .A(KEYINPUT73), .B(n599), .ZN(n600) );
  NOR2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n604), .B(KEYINPUT15), .ZN(n1001) );
  INV_X1 U678 ( .A(n1001), .ZN(n628) );
  NAND2_X1 U679 ( .A1(n658), .A2(G1341), .ZN(n605) );
  XNOR2_X1 U680 ( .A(KEYINPUT95), .B(n605), .ZN(n611) );
  INV_X1 U681 ( .A(G1996), .ZN(n607) );
  XNOR2_X1 U682 ( .A(n608), .B(KEYINPUT26), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n609), .B(KEYINPUT65), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n805), .A2(G56), .ZN(n614) );
  XNOR2_X1 U685 ( .A(KEYINPUT14), .B(n614), .ZN(n621) );
  NAND2_X1 U686 ( .A1(G81), .A2(n800), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G68), .A2(n801), .ZN(n617) );
  NAND2_X1 U688 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U689 ( .A(KEYINPUT13), .B(n619), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U691 ( .A(n622), .B(KEYINPUT71), .ZN(n624) );
  NAND2_X1 U692 ( .A1(G43), .A2(n806), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X2 U694 ( .A(KEYINPUT72), .B(n625), .ZN(n1004) );
  INV_X1 U695 ( .A(n629), .ZN(n627) );
  NAND2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n635) );
  NAND2_X1 U697 ( .A1(n1001), .A2(n629), .ZN(n633) );
  NOR2_X1 U698 ( .A1(G2067), .A2(n658), .ZN(n631) );
  INV_X1 U699 ( .A(n658), .ZN(n648) );
  NOR2_X1 U700 ( .A1(n648), .A2(G1348), .ZN(n630) );
  NOR2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n635), .A2(n634), .ZN(n642) );
  INV_X1 U704 ( .A(G299), .ZN(n815) );
  INV_X1 U705 ( .A(G2072), .ZN(n876) );
  NOR2_X1 U706 ( .A1(n658), .A2(n876), .ZN(n637) );
  XOR2_X1 U707 ( .A(KEYINPUT93), .B(KEYINPUT27), .Z(n636) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n658), .A2(G1956), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U711 ( .A(KEYINPUT94), .B(n640), .Z(n643) );
  NAND2_X1 U712 ( .A1(n815), .A2(n643), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n646) );
  NOR2_X1 U714 ( .A1(n815), .A2(n643), .ZN(n644) );
  XOR2_X1 U715 ( .A(n644), .B(KEYINPUT28), .Z(n645) );
  NAND2_X1 U716 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n647), .B(KEYINPUT29), .ZN(n681) );
  NAND2_X1 U718 ( .A1(n658), .A2(G1961), .ZN(n650) );
  XOR2_X1 U719 ( .A(G2078), .B(KEYINPUT25), .Z(n915) );
  NAND2_X1 U720 ( .A1(n915), .A2(n648), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U722 ( .A(KEYINPUT92), .B(n651), .Z(n665) );
  AND2_X1 U723 ( .A1(n665), .A2(G171), .ZN(n680) );
  NOR2_X1 U724 ( .A1(G1971), .A2(n706), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(KEYINPUT98), .ZN(n654) );
  NOR2_X1 U726 ( .A1(n658), .A2(G2090), .ZN(n653) );
  NOR2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n655), .A2(G303), .ZN(n670) );
  INV_X1 U729 ( .A(n670), .ZN(n656) );
  NOR2_X1 U730 ( .A1(n656), .A2(G286), .ZN(n672) );
  OR2_X1 U731 ( .A1(n680), .A2(n672), .ZN(n657) );
  OR2_X1 U732 ( .A1(n681), .A2(n657), .ZN(n674) );
  INV_X1 U733 ( .A(KEYINPUT31), .ZN(n669) );
  INV_X1 U734 ( .A(KEYINPUT91), .ZN(n659) );
  NOR2_X1 U735 ( .A1(n685), .A2(n679), .ZN(n661) );
  AND2_X1 U736 ( .A1(n661), .A2(G8), .ZN(n663) );
  NOR2_X1 U737 ( .A1(n664), .A2(G168), .ZN(n667) );
  NOR2_X1 U738 ( .A1(G171), .A2(n665), .ZN(n666) );
  NOR2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n669), .B(n668), .ZN(n682) );
  AND2_X1 U741 ( .A1(n682), .A2(n670), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U743 ( .A(n675), .B(KEYINPUT99), .ZN(n677) );
  INV_X1 U744 ( .A(G8), .ZN(n676) );
  OR2_X2 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n678), .B(KEYINPUT32), .ZN(n689) );
  NAND2_X1 U747 ( .A1(G8), .A2(n679), .ZN(n687) );
  OR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n683) );
  AND2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U751 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n699) );
  NOR2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n949) );
  NOR2_X1 U754 ( .A1(G1971), .A2(G303), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n949), .A2(n690), .ZN(n691) );
  NAND2_X1 U756 ( .A1(n699), .A2(n691), .ZN(n692) );
  XNOR2_X1 U757 ( .A(n692), .B(KEYINPUT100), .ZN(n693) );
  NAND2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n950) );
  NAND2_X1 U759 ( .A1(n693), .A2(n950), .ZN(n695) );
  NOR2_X1 U760 ( .A1(n706), .A2(n696), .ZN(n705) );
  NOR2_X1 U761 ( .A1(G2090), .A2(G303), .ZN(n697) );
  NAND2_X1 U762 ( .A1(G8), .A2(n697), .ZN(n698) );
  NAND2_X1 U763 ( .A1(n699), .A2(n698), .ZN(n700) );
  AND2_X1 U764 ( .A1(n700), .A2(n706), .ZN(n711) );
  OR2_X2 U765 ( .A1(KEYINPUT33), .A2(n711), .ZN(n703) );
  NOR2_X1 U766 ( .A1(G1981), .A2(G305), .ZN(n701) );
  XOR2_X1 U767 ( .A(n701), .B(KEYINPUT24), .Z(n702) );
  NOR2_X1 U768 ( .A1(n706), .A2(n702), .ZN(n713) );
  OR2_X2 U769 ( .A1(n703), .A2(n713), .ZN(n704) );
  OR2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n749) );
  NAND2_X1 U771 ( .A1(n949), .A2(KEYINPUT33), .ZN(n707) );
  NOR2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n709) );
  XOR2_X1 U773 ( .A(G1981), .B(G305), .Z(n938) );
  INV_X1 U774 ( .A(n938), .ZN(n708) );
  NOR2_X1 U775 ( .A1(n709), .A2(n708), .ZN(n710) );
  OR2_X1 U776 ( .A1(n711), .A2(n710), .ZN(n712) );
  OR2_X1 U777 ( .A1(n713), .A2(n712), .ZN(n745) );
  NOR2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n760) );
  NAND2_X1 U779 ( .A1(n987), .A2(G140), .ZN(n716) );
  XNOR2_X1 U780 ( .A(n716), .B(KEYINPUT88), .ZN(n718) );
  NAND2_X1 U781 ( .A1(G104), .A2(n986), .ZN(n717) );
  NAND2_X1 U782 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U783 ( .A(KEYINPUT34), .B(n719), .ZN(n724) );
  NAND2_X1 U784 ( .A1(G128), .A2(n982), .ZN(n721) );
  NAND2_X1 U785 ( .A1(G116), .A2(n983), .ZN(n720) );
  NAND2_X1 U786 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U787 ( .A(KEYINPUT35), .B(n722), .Z(n723) );
  NOR2_X1 U788 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U789 ( .A(KEYINPUT36), .B(n725), .ZN(n996) );
  XNOR2_X1 U790 ( .A(G2067), .B(KEYINPUT37), .ZN(n758) );
  NOR2_X1 U791 ( .A1(n996), .A2(n758), .ZN(n885) );
  NAND2_X1 U792 ( .A1(n760), .A2(n885), .ZN(n756) );
  NAND2_X1 U793 ( .A1(n987), .A2(G131), .ZN(n728) );
  NAND2_X1 U794 ( .A1(G107), .A2(n983), .ZN(n726) );
  XOR2_X1 U795 ( .A(KEYINPUT89), .B(n726), .Z(n727) );
  NAND2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n732) );
  NAND2_X1 U797 ( .A1(G95), .A2(n986), .ZN(n730) );
  NAND2_X1 U798 ( .A1(G119), .A2(n982), .ZN(n729) );
  NAND2_X1 U799 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n979) );
  XOR2_X1 U801 ( .A(G1991), .B(KEYINPUT90), .Z(n916) );
  NOR2_X1 U802 ( .A1(n979), .A2(n916), .ZN(n741) );
  NAND2_X1 U803 ( .A1(n986), .A2(G105), .ZN(n733) );
  XNOR2_X1 U804 ( .A(n733), .B(KEYINPUT38), .ZN(n735) );
  NAND2_X1 U805 ( .A1(G117), .A2(n983), .ZN(n734) );
  NAND2_X1 U806 ( .A1(n735), .A2(n734), .ZN(n739) );
  NAND2_X1 U807 ( .A1(G141), .A2(n987), .ZN(n737) );
  NAND2_X1 U808 ( .A1(G129), .A2(n982), .ZN(n736) );
  NAND2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U810 ( .A1(n739), .A2(n738), .ZN(n974) );
  NOR2_X1 U811 ( .A1(n974), .A2(n607), .ZN(n740) );
  NOR2_X1 U812 ( .A1(n741), .A2(n740), .ZN(n866) );
  INV_X1 U813 ( .A(n760), .ZN(n742) );
  NOR2_X1 U814 ( .A1(n866), .A2(n742), .ZN(n752) );
  INV_X1 U815 ( .A(n752), .ZN(n743) );
  AND2_X1 U816 ( .A1(n756), .A2(n743), .ZN(n744) );
  NAND2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n747) );
  XNOR2_X1 U818 ( .A(G1986), .B(G290), .ZN(n954) );
  AND2_X1 U819 ( .A1(n954), .A2(n760), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n763) );
  AND2_X1 U822 ( .A1(n979), .A2(n916), .ZN(n855) );
  NOR2_X1 U823 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U824 ( .A1(n855), .A2(n750), .ZN(n751) );
  NOR2_X1 U825 ( .A1(n752), .A2(n751), .ZN(n754) );
  AND2_X1 U826 ( .A1(n974), .A2(n607), .ZN(n753) );
  XNOR2_X1 U827 ( .A(n753), .B(KEYINPUT102), .ZN(n858) );
  NOR2_X1 U828 ( .A1(n754), .A2(n858), .ZN(n755) );
  XNOR2_X1 U829 ( .A(n755), .B(KEYINPUT39), .ZN(n757) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U831 ( .A1(n996), .A2(n758), .ZN(n882) );
  NAND2_X1 U832 ( .A1(n759), .A2(n882), .ZN(n761) );
  NAND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U834 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U835 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U836 ( .A(G2443), .B(G2451), .Z(n766) );
  XNOR2_X1 U837 ( .A(G2454), .B(G2435), .ZN(n765) );
  XNOR2_X1 U838 ( .A(n766), .B(n765), .ZN(n773) );
  XOR2_X1 U839 ( .A(G2427), .B(G2446), .Z(n768) );
  XNOR2_X1 U840 ( .A(G1341), .B(G2430), .ZN(n767) );
  XNOR2_X1 U841 ( .A(n768), .B(n767), .ZN(n769) );
  XOR2_X1 U842 ( .A(n769), .B(G2438), .Z(n771) );
  XNOR2_X1 U843 ( .A(G1348), .B(KEYINPUT103), .ZN(n770) );
  XNOR2_X1 U844 ( .A(n771), .B(n770), .ZN(n772) );
  XNOR2_X1 U845 ( .A(n773), .B(n772), .ZN(n774) );
  AND2_X1 U846 ( .A1(n774), .A2(G14), .ZN(G401) );
  AND2_X1 U847 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U848 ( .A(G57), .ZN(G237) );
  INV_X1 U849 ( .A(G132), .ZN(G219) );
  INV_X1 U850 ( .A(G82), .ZN(G220) );
  NAND2_X1 U851 ( .A1(G7), .A2(G661), .ZN(n776) );
  XNOR2_X1 U852 ( .A(n776), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U853 ( .A(G223), .ZN(n843) );
  NAND2_X1 U854 ( .A1(n843), .A2(G567), .ZN(n777) );
  XNOR2_X1 U855 ( .A(n777), .B(KEYINPUT11), .ZN(n778) );
  XNOR2_X1 U856 ( .A(KEYINPUT69), .B(n778), .ZN(G234) );
  INV_X1 U857 ( .A(G860), .ZN(n783) );
  OR2_X1 U858 ( .A1(n783), .A2(n1004), .ZN(G153) );
  INV_X1 U859 ( .A(G171), .ZN(G301) );
  NAND2_X1 U860 ( .A1(G868), .A2(G301), .ZN(n780) );
  OR2_X1 U861 ( .A1(n1001), .A2(G868), .ZN(n779) );
  NAND2_X1 U862 ( .A1(n780), .A2(n779), .ZN(G284) );
  INV_X1 U863 ( .A(G868), .ZN(n824) );
  NOR2_X1 U864 ( .A1(G286), .A2(n824), .ZN(n782) );
  NOR2_X1 U865 ( .A1(G868), .A2(G299), .ZN(n781) );
  NOR2_X1 U866 ( .A1(n782), .A2(n781), .ZN(G297) );
  NAND2_X1 U867 ( .A1(n783), .A2(G559), .ZN(n784) );
  NAND2_X1 U868 ( .A1(n784), .A2(n1001), .ZN(n785) );
  XNOR2_X1 U869 ( .A(n785), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U870 ( .A1(n1004), .A2(G868), .ZN(n788) );
  NAND2_X1 U871 ( .A1(n1001), .A2(G868), .ZN(n786) );
  NOR2_X1 U872 ( .A1(G559), .A2(n786), .ZN(n787) );
  NOR2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U874 ( .A(KEYINPUT76), .B(n789), .ZN(G282) );
  NAND2_X1 U875 ( .A1(G123), .A2(n982), .ZN(n790) );
  XNOR2_X1 U876 ( .A(n790), .B(KEYINPUT18), .ZN(n793) );
  NAND2_X1 U877 ( .A1(G111), .A2(n983), .ZN(n791) );
  XOR2_X1 U878 ( .A(KEYINPUT77), .B(n791), .Z(n792) );
  NAND2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n797) );
  NAND2_X1 U880 ( .A1(G99), .A2(n986), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G135), .A2(n987), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n973) );
  XNOR2_X1 U884 ( .A(n973), .B(G2096), .ZN(n799) );
  INV_X1 U885 ( .A(G2100), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(G156) );
  NAND2_X1 U887 ( .A1(G93), .A2(n800), .ZN(n803) );
  NAND2_X1 U888 ( .A1(G80), .A2(n801), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U890 ( .A(KEYINPUT80), .B(n804), .ZN(n810) );
  NAND2_X1 U891 ( .A1(G67), .A2(n805), .ZN(n808) );
  NAND2_X1 U892 ( .A1(G55), .A2(n806), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n808), .A2(n807), .ZN(n809) );
  OR2_X1 U894 ( .A1(n810), .A2(n809), .ZN(n825) );
  XOR2_X1 U895 ( .A(KEYINPUT78), .B(n1004), .Z(n812) );
  NAND2_X1 U896 ( .A1(G559), .A2(n1001), .ZN(n811) );
  XNOR2_X1 U897 ( .A(n812), .B(n811), .ZN(n822) );
  XNOR2_X1 U898 ( .A(KEYINPUT79), .B(n822), .ZN(n813) );
  NOR2_X1 U899 ( .A1(G860), .A2(n813), .ZN(n814) );
  XOR2_X1 U900 ( .A(n825), .B(n814), .Z(G145) );
  INV_X1 U901 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U902 ( .A(n815), .B(G166), .ZN(n821) );
  XOR2_X1 U903 ( .A(n825), .B(G290), .Z(n816) );
  XNOR2_X1 U904 ( .A(n816), .B(G305), .ZN(n817) );
  XNOR2_X1 U905 ( .A(KEYINPUT84), .B(n817), .ZN(n819) );
  XNOR2_X1 U906 ( .A(G288), .B(KEYINPUT19), .ZN(n818) );
  XNOR2_X1 U907 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U908 ( .A(n821), .B(n820), .ZN(n1000) );
  XOR2_X1 U909 ( .A(n1000), .B(n822), .Z(n823) );
  NOR2_X1 U910 ( .A1(n824), .A2(n823), .ZN(n827) );
  NOR2_X1 U911 ( .A1(G868), .A2(n825), .ZN(n826) );
  NOR2_X1 U912 ( .A1(n827), .A2(n826), .ZN(G295) );
  NAND2_X1 U913 ( .A1(G2078), .A2(G2084), .ZN(n828) );
  XNOR2_X1 U914 ( .A(n828), .B(KEYINPUT85), .ZN(n829) );
  XNOR2_X1 U915 ( .A(n829), .B(KEYINPUT20), .ZN(n830) );
  NAND2_X1 U916 ( .A1(n830), .A2(G2090), .ZN(n831) );
  XNOR2_X1 U917 ( .A(n831), .B(KEYINPUT86), .ZN(n832) );
  XNOR2_X1 U918 ( .A(n832), .B(KEYINPUT21), .ZN(n833) );
  NAND2_X1 U919 ( .A1(n833), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U920 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U921 ( .A1(G220), .A2(G219), .ZN(n834) );
  XOR2_X1 U922 ( .A(KEYINPUT22), .B(n834), .Z(n835) );
  NOR2_X1 U923 ( .A1(G218), .A2(n835), .ZN(n836) );
  NAND2_X1 U924 ( .A1(G96), .A2(n836), .ZN(n967) );
  NAND2_X1 U925 ( .A1(n967), .A2(G2106), .ZN(n840) );
  NAND2_X1 U926 ( .A1(G69), .A2(G120), .ZN(n837) );
  NOR2_X1 U927 ( .A1(G237), .A2(n837), .ZN(n838) );
  NAND2_X1 U928 ( .A1(G108), .A2(n838), .ZN(n968) );
  NAND2_X1 U929 ( .A1(n968), .A2(G567), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(n969) );
  NAND2_X1 U931 ( .A1(G661), .A2(G483), .ZN(n841) );
  XOR2_X1 U932 ( .A(KEYINPUT87), .B(n841), .Z(n842) );
  NOR2_X1 U933 ( .A1(n969), .A2(n842), .ZN(n846) );
  NAND2_X1 U934 ( .A1(n846), .A2(G36), .ZN(G176) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U937 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U939 ( .A1(n846), .A2(n845), .ZN(G188) );
  XOR2_X1 U940 ( .A(G96), .B(KEYINPUT104), .Z(G221) );
  NAND2_X1 U942 ( .A1(G124), .A2(n982), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n847), .B(KEYINPUT108), .ZN(n848) );
  XNOR2_X1 U944 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U945 ( .A1(G112), .A2(n983), .ZN(n849) );
  NAND2_X1 U946 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U947 ( .A1(G100), .A2(n986), .ZN(n852) );
  NAND2_X1 U948 ( .A1(G136), .A2(n987), .ZN(n851) );
  NAND2_X1 U949 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U950 ( .A1(n854), .A2(n853), .ZN(G162) );
  NOR2_X1 U951 ( .A1(n855), .A2(n973), .ZN(n861) );
  XOR2_X1 U952 ( .A(G2090), .B(G162), .Z(n856) );
  XNOR2_X1 U953 ( .A(KEYINPUT116), .B(n856), .ZN(n857) );
  NOR2_X1 U954 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U955 ( .A(KEYINPUT51), .B(n859), .Z(n860) );
  NAND2_X1 U956 ( .A1(n861), .A2(n860), .ZN(n864) );
  XNOR2_X1 U957 ( .A(G2084), .B(G160), .ZN(n862) );
  XNOR2_X1 U958 ( .A(KEYINPUT115), .B(n862), .ZN(n863) );
  NOR2_X1 U959 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U960 ( .A1(n866), .A2(n865), .ZN(n881) );
  XOR2_X1 U961 ( .A(G164), .B(G2078), .Z(n878) );
  NAND2_X1 U962 ( .A1(G103), .A2(n986), .ZN(n868) );
  NAND2_X1 U963 ( .A1(G139), .A2(n987), .ZN(n867) );
  NAND2_X1 U964 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U965 ( .A1(n983), .A2(G115), .ZN(n869) );
  XOR2_X1 U966 ( .A(KEYINPUT111), .B(n869), .Z(n871) );
  NAND2_X1 U967 ( .A1(n982), .A2(G127), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U969 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U970 ( .A1(n874), .A2(n873), .ZN(n970) );
  XOR2_X1 U971 ( .A(n970), .B(KEYINPUT117), .Z(n875) );
  XNOR2_X1 U972 ( .A(n876), .B(n875), .ZN(n877) );
  NOR2_X1 U973 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U974 ( .A(KEYINPUT50), .B(n879), .Z(n880) );
  NOR2_X1 U975 ( .A1(n881), .A2(n880), .ZN(n883) );
  NAND2_X1 U976 ( .A1(n883), .A2(n882), .ZN(n884) );
  NOR2_X1 U977 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U978 ( .A(KEYINPUT52), .B(n886), .Z(n887) );
  XNOR2_X1 U979 ( .A(n887), .B(KEYINPUT118), .ZN(n888) );
  NAND2_X1 U980 ( .A1(n888), .A2(G29), .ZN(n937) );
  XNOR2_X1 U981 ( .A(G1971), .B(G22), .ZN(n890) );
  XNOR2_X1 U982 ( .A(G23), .B(G1976), .ZN(n889) );
  NOR2_X1 U983 ( .A1(n890), .A2(n889), .ZN(n892) );
  XOR2_X1 U984 ( .A(G1986), .B(G24), .Z(n891) );
  NAND2_X1 U985 ( .A1(n892), .A2(n891), .ZN(n894) );
  XOR2_X1 U986 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n893) );
  XNOR2_X1 U987 ( .A(n894), .B(n893), .ZN(n898) );
  XNOR2_X1 U988 ( .A(G1966), .B(G21), .ZN(n896) );
  XNOR2_X1 U989 ( .A(G5), .B(G1961), .ZN(n895) );
  NOR2_X1 U990 ( .A1(n896), .A2(n895), .ZN(n897) );
  NAND2_X1 U991 ( .A1(n898), .A2(n897), .ZN(n908) );
  XOR2_X1 U992 ( .A(G1348), .B(KEYINPUT59), .Z(n899) );
  XNOR2_X1 U993 ( .A(G4), .B(n899), .ZN(n901) );
  XNOR2_X1 U994 ( .A(G20), .B(G1956), .ZN(n900) );
  NOR2_X1 U995 ( .A1(n901), .A2(n900), .ZN(n905) );
  XNOR2_X1 U996 ( .A(G1341), .B(G19), .ZN(n903) );
  XNOR2_X1 U997 ( .A(G1981), .B(G6), .ZN(n902) );
  NOR2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n904) );
  NAND2_X1 U999 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(KEYINPUT60), .B(n906), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n909), .B(KEYINPUT61), .ZN(n911) );
  XNOR2_X1 U1003 ( .A(G16), .B(KEYINPUT125), .ZN(n910) );
  NAND2_X1 U1004 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1005 ( .A1(G11), .A2(n912), .ZN(n935) );
  XNOR2_X1 U1006 ( .A(G1996), .B(G32), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(G2072), .B(G33), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(n914), .A2(n913), .ZN(n925) );
  XOR2_X1 U1009 ( .A(n915), .B(G27), .Z(n920) );
  XNOR2_X1 U1010 ( .A(n916), .B(G25), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(n917), .A2(G28), .ZN(n918) );
  XNOR2_X1 U1012 ( .A(n918), .B(KEYINPUT119), .ZN(n919) );
  NAND2_X1 U1013 ( .A1(n920), .A2(n919), .ZN(n923) );
  XNOR2_X1 U1014 ( .A(KEYINPUT120), .B(G2067), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(G26), .B(n921), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1017 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1018 ( .A(n926), .B(KEYINPUT53), .ZN(n929) );
  XOR2_X1 U1019 ( .A(G2084), .B(KEYINPUT54), .Z(n927) );
  XNOR2_X1 U1020 ( .A(G34), .B(n927), .ZN(n928) );
  NAND2_X1 U1021 ( .A1(n929), .A2(n928), .ZN(n931) );
  XNOR2_X1 U1022 ( .A(G35), .B(G2090), .ZN(n930) );
  NOR2_X1 U1023 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1024 ( .A1(G29), .A2(n932), .ZN(n933) );
  XOR2_X1 U1025 ( .A(KEYINPUT55), .B(n933), .Z(n934) );
  NOR2_X1 U1026 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1027 ( .A1(n937), .A2(n936), .ZN(n965) );
  XNOR2_X1 U1028 ( .A(G1966), .B(G168), .ZN(n939) );
  NAND2_X1 U1029 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1030 ( .A(KEYINPUT57), .B(n940), .Z(n961) );
  XNOR2_X1 U1031 ( .A(G1348), .B(n1001), .ZN(n942) );
  XNOR2_X1 U1032 ( .A(G171), .B(G1961), .ZN(n941) );
  NAND2_X1 U1033 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1034 ( .A(KEYINPUT121), .B(n943), .ZN(n947) );
  XNOR2_X1 U1035 ( .A(G299), .B(G1956), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(G303), .B(G1971), .ZN(n944) );
  NOR2_X1 U1037 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n958) );
  XNOR2_X1 U1039 ( .A(G1341), .B(n1004), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(n948), .B(KEYINPUT123), .ZN(n956) );
  INV_X1 U1041 ( .A(n949), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1043 ( .A(KEYINPUT122), .B(n952), .ZN(n953) );
  NOR2_X1 U1044 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1045 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1046 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1047 ( .A(KEYINPUT124), .B(n959), .Z(n960) );
  NOR2_X1 U1048 ( .A1(n961), .A2(n960), .ZN(n963) );
  XOR2_X1 U1049 ( .A(G16), .B(KEYINPUT56), .Z(n962) );
  NOR2_X1 U1050 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1051 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1052 ( .A(n966), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1053 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1054 ( .A(G120), .ZN(G236) );
  INV_X1 U1055 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1056 ( .A1(n968), .A2(n967), .ZN(G325) );
  INV_X1 U1057 ( .A(G325), .ZN(G261) );
  INV_X1 U1058 ( .A(n969), .ZN(G319) );
  XOR2_X1 U1059 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n972) );
  XNOR2_X1 U1060 ( .A(n970), .B(KEYINPUT46), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(n972), .B(n971), .ZN(n978) );
  XOR2_X1 U1062 ( .A(n973), .B(G162), .Z(n976) );
  XNOR2_X1 U1063 ( .A(G160), .B(n974), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(n976), .B(n975), .ZN(n977) );
  XOR2_X1 U1065 ( .A(n978), .B(n977), .Z(n981) );
  XNOR2_X1 U1066 ( .A(G164), .B(n979), .ZN(n980) );
  XNOR2_X1 U1067 ( .A(n981), .B(n980), .ZN(n998) );
  NAND2_X1 U1068 ( .A1(G130), .A2(n982), .ZN(n985) );
  NAND2_X1 U1069 ( .A1(G118), .A2(n983), .ZN(n984) );
  NAND2_X1 U1070 ( .A1(n985), .A2(n984), .ZN(n994) );
  XNOR2_X1 U1071 ( .A(KEYINPUT45), .B(KEYINPUT110), .ZN(n992) );
  NAND2_X1 U1072 ( .A1(n986), .A2(G106), .ZN(n990) );
  NAND2_X1 U1073 ( .A1(n987), .A2(G142), .ZN(n988) );
  XOR2_X1 U1074 ( .A(KEYINPUT109), .B(n988), .Z(n989) );
  NAND2_X1 U1075 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1076 ( .A(n992), .B(n991), .Z(n993) );
  NOR2_X1 U1077 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1078 ( .A(n996), .B(n995), .Z(n997) );
  XNOR2_X1 U1079 ( .A(n998), .B(n997), .ZN(n999) );
  NOR2_X1 U1080 ( .A1(G37), .A2(n999), .ZN(G395) );
  XOR2_X1 U1081 ( .A(KEYINPUT113), .B(n1000), .Z(n1003) );
  XNOR2_X1 U1082 ( .A(G171), .B(n1001), .ZN(n1002) );
  XNOR2_X1 U1083 ( .A(n1003), .B(n1002), .ZN(n1006) );
  XOR2_X1 U1084 ( .A(G286), .B(n1004), .Z(n1005) );
  XNOR2_X1 U1085 ( .A(n1006), .B(n1005), .ZN(n1007) );
  NOR2_X1 U1086 ( .A1(G37), .A2(n1007), .ZN(G397) );
  XOR2_X1 U1087 ( .A(KEYINPUT105), .B(G2474), .Z(n1009) );
  XNOR2_X1 U1088 ( .A(G1966), .B(G1981), .ZN(n1008) );
  XNOR2_X1 U1089 ( .A(n1009), .B(n1008), .ZN(n1019) );
  XOR2_X1 U1090 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n1011) );
  XNOR2_X1 U1091 ( .A(G1991), .B(G1986), .ZN(n1010) );
  XNOR2_X1 U1092 ( .A(n1011), .B(n1010), .ZN(n1015) );
  XOR2_X1 U1093 ( .A(G1976), .B(G1971), .Z(n1013) );
  XNOR2_X1 U1094 ( .A(G1961), .B(G1956), .ZN(n1012) );
  XNOR2_X1 U1095 ( .A(n1013), .B(n1012), .ZN(n1014) );
  XOR2_X1 U1096 ( .A(n1015), .B(n1014), .Z(n1017) );
  XNOR2_X1 U1097 ( .A(G1996), .B(KEYINPUT106), .ZN(n1016) );
  XNOR2_X1 U1098 ( .A(n1017), .B(n1016), .ZN(n1018) );
  XOR2_X1 U1099 ( .A(n1019), .B(n1018), .Z(G229) );
  XOR2_X1 U1100 ( .A(G2100), .B(G2096), .Z(n1021) );
  XNOR2_X1 U1101 ( .A(G2067), .B(G2090), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(n1021), .B(n1020), .ZN(n1025) );
  XOR2_X1 U1103 ( .A(G2678), .B(KEYINPUT42), .Z(n1023) );
  XNOR2_X1 U1104 ( .A(G2072), .B(KEYINPUT43), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(n1023), .B(n1022), .ZN(n1024) );
  XOR2_X1 U1106 ( .A(n1025), .B(n1024), .Z(n1027) );
  XNOR2_X1 U1107 ( .A(G2078), .B(G2084), .ZN(n1026) );
  XNOR2_X1 U1108 ( .A(n1027), .B(n1026), .ZN(G227) );
  NOR2_X1 U1109 ( .A1(G395), .A2(G397), .ZN(n1028) );
  XNOR2_X1 U1110 ( .A(n1028), .B(KEYINPUT114), .ZN(n1029) );
  NAND2_X1 U1111 ( .A1(G319), .A2(n1029), .ZN(n1030) );
  NOR2_X1 U1112 ( .A1(G401), .A2(n1030), .ZN(n1033) );
  NOR2_X1 U1113 ( .A1(G229), .A2(G227), .ZN(n1031) );
  XOR2_X1 U1114 ( .A(KEYINPUT49), .B(n1031), .Z(n1032) );
  NAND2_X1 U1115 ( .A1(n1033), .A2(n1032), .ZN(G225) );
  INV_X1 U1116 ( .A(G225), .ZN(G308) );
  INV_X1 U1117 ( .A(G108), .ZN(G238) );
endmodule

