//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT66), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n226), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT64), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n231));
  NAND4_X1  g0031(.A1(new_n227), .A2(new_n228), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(new_n209), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n218), .B1(new_n212), .B2(new_n211), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n202), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n206), .A2(G20), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT70), .ZN(new_n257));
  INV_X1    g0057(.A(new_n213), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n258), .B1(new_n208), .B2(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n259), .A3(new_n254), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n255), .B1(new_n261), .B2(new_n202), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n207), .A2(G33), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT69), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT8), .B(G58), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n259), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT9), .ZN(new_n274));
  INV_X1    g0074(.A(G200), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G33), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n276), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G222), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G77), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G223), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n287), .B1(new_n288), .B2(new_n285), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n294));
  INV_X1    g0094(.A(G274), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G41), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n258), .B1(new_n277), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n294), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n296), .B1(new_n300), .B2(G226), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n274), .B1(new_n275), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  OR3_X1    g0106(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT10), .B1(new_n304), .B2(new_n306), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n302), .A2(G169), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n302), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n273), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n254), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n266), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n260), .B2(new_n266), .ZN(new_n317));
  INV_X1    g0117(.A(G58), .ZN(new_n318));
  INV_X1    g0118(.A(G68), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n320), .A2(new_n201), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(G20), .B1(G159), .B2(new_n268), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT75), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n277), .ZN(new_n324));
  NAND2_X1  g0124(.A1(KEYINPUT75), .A2(G33), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(KEYINPUT3), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(G20), .B1(new_n326), .B2(new_n282), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT7), .ZN(new_n328));
  OAI21_X1  g0128(.A(G68), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT75), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT75), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n278), .B1(new_n332), .B2(KEYINPUT3), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n333), .A2(KEYINPUT7), .A3(G20), .ZN(new_n334));
  OAI211_X1 g0134(.A(KEYINPUT16), .B(new_n322), .C1(new_n329), .C2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n335), .A2(new_n271), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n281), .A2(new_n207), .A3(new_n284), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n283), .B1(new_n332), .B2(KEYINPUT3), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n328), .A2(G20), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n337), .A2(new_n328), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n322), .B1(new_n340), .B2(new_n319), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n317), .B1(new_n336), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G226), .A2(G1698), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n290), .B2(G1698), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n333), .A2(new_n346), .B1(G33), .B2(G87), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT77), .B1(new_n347), .B2(new_n298), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n296), .B1(new_n300), .B2(G232), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n326), .A2(new_n282), .A3(new_n346), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n277), .B2(new_n221), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT77), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(new_n292), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n348), .A2(new_n311), .A3(new_n349), .A4(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n349), .B1(new_n298), .B2(new_n347), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT18), .B1(new_n344), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n355), .A2(new_n275), .ZN(new_n360));
  INV_X1    g0160(.A(new_n296), .ZN(new_n361));
  INV_X1    g0161(.A(G232), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(new_n299), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(G190), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n348), .A2(new_n353), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n317), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n341), .A2(new_n342), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n335), .A2(new_n271), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT17), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT18), .ZN(new_n374));
  INV_X1    g0174(.A(new_n358), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n344), .A2(KEYINPUT17), .A3(new_n366), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n359), .A2(new_n372), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n261), .A2(G77), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT15), .B(G87), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n380), .A2(new_n263), .B1(new_n207), .B2(new_n288), .ZN(new_n381));
  INV_X1    g0181(.A(new_n268), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n265), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n271), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n315), .A2(new_n288), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n379), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G244), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n361), .B1(new_n299), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n285), .A2(G232), .A3(new_n286), .ZN(new_n389));
  INV_X1    g0189(.A(G107), .ZN(new_n390));
  INV_X1    g0190(.A(G238), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n389), .B1(new_n390), .B2(new_n285), .C1(new_n289), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n392), .B2(new_n292), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n386), .B1(new_n393), .B2(G169), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT71), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT71), .B(new_n386), .C1(new_n393), .C2(G169), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n311), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n386), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n393), .A2(new_n305), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n393), .A2(G200), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n314), .A2(new_n378), .A3(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n264), .A2(G77), .B1(G20), .B2(new_n319), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT74), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n202), .B2(new_n382), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n406), .A2(new_n407), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n271), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT11), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(KEYINPUT11), .B(new_n271), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n206), .A2(G13), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n415), .A2(new_n207), .A3(G68), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT12), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n261), .B2(G68), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n413), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT68), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT68), .B1(new_n282), .B2(new_n283), .ZN(new_n421));
  OAI211_X1 g0221(.A(G226), .B(new_n286), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(G232), .B(G1698), .C1(new_n420), .C2(new_n421), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G97), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n292), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT13), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n296), .B1(new_n300), .B2(G238), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT73), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n428), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT13), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT73), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n426), .A2(new_n433), .A3(new_n427), .A4(new_n428), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n430), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n435), .A2(new_n311), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT72), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n426), .A2(KEYINPUT72), .A3(new_n427), .A4(new_n428), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n439), .A3(new_n432), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n440), .A2(G169), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT14), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n436), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n440), .A2(new_n442), .A3(G169), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n419), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n419), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n440), .A2(G200), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n446), .B(new_n447), .C1(new_n305), .C2(new_n435), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n405), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G257), .A2(G1698), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n222), .B2(G1698), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n326), .A2(new_n282), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n324), .A2(new_n325), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G294), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT84), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n453), .A2(KEYINPUT84), .A3(new_n455), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n292), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  AND2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n465), .A2(new_n295), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n298), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G264), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n460), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G169), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n311), .B2(new_n470), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n206), .A2(G33), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n259), .A2(new_n254), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n390), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n253), .A2(G20), .A3(new_n390), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT25), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT83), .B1(new_n207), .B2(G107), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT23), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  OR2_X1    g0282(.A1(KEYINPUT79), .A2(G116), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT79), .A2(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n454), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n481), .B(new_n482), .C1(new_n486), .C2(G20), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n221), .A2(KEYINPUT22), .A3(G20), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n285), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n326), .A2(new_n207), .A3(G87), .A4(new_n282), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT22), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n487), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT24), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n271), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n492), .A2(KEYINPUT24), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n478), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n472), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT21), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G264), .A2(G1698), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n224), .B2(G1698), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n333), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n281), .A2(G303), .A3(new_n284), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n298), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G270), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n466), .B1(new_n504), .B2(new_n467), .ZN(new_n505));
  OAI21_X1  g0305(.A(G169), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G116), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n474), .A2(new_n507), .B1(new_n254), .B2(new_n485), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT20), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n207), .B1(new_n483), .B2(new_n484), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n277), .A2(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  AOI21_X1  g0312(.A(G20), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n509), .B1(new_n514), .B2(new_n259), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n271), .B(KEYINPUT20), .C1(new_n513), .C2(new_n510), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n508), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n498), .B1(new_n506), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT82), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT82), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(new_n498), .C1(new_n506), .C2(new_n517), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n506), .A2(new_n517), .A3(new_n498), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n503), .A2(new_n505), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G179), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(new_n517), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n524), .A2(G200), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n503), .A2(new_n505), .A3(G190), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n517), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n497), .A2(new_n522), .A3(new_n527), .A4(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n333), .A2(new_n207), .A3(G68), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G87), .A2(G97), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(new_n390), .B1(new_n424), .B2(new_n207), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n207), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n534), .A2(new_n535), .B1(new_n424), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n271), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n315), .A2(new_n380), .ZN(new_n540));
  INV_X1    g0340(.A(new_n474), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G87), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT80), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n326), .A2(G244), .A3(G1698), .A4(new_n282), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n391), .A2(G1698), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n326), .A2(new_n282), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n486), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n292), .ZN(new_n549));
  OAI21_X1  g0349(.A(G250), .B1(new_n461), .B2(G1), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n462), .A2(G274), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n292), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n544), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  AOI211_X1 g0354(.A(KEYINPUT80), .B(new_n552), .C1(new_n548), .C2(new_n292), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n543), .B1(new_n556), .B2(G200), .ZN(new_n557));
  OAI21_X1  g0357(.A(G190), .B1(new_n554), .B2(new_n555), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT81), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n560), .B(G190), .C1(new_n554), .C2(new_n555), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n556), .A2(new_n356), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n311), .B1(new_n554), .B2(new_n555), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n539), .B(new_n540), .C1(new_n380), .C2(new_n474), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n531), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n315), .A2(new_n223), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n474), .B2(new_n223), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n390), .A2(KEYINPUT6), .A3(G97), .ZN(new_n571));
  XOR2_X1   g0371(.A(G97), .B(G107), .Z(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(KEYINPUT6), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(G20), .B1(G77), .B2(new_n268), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n340), .B2(new_n390), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n570), .B1(new_n575), .B2(new_n271), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n466), .B1(new_n224), .B2(new_n467), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n326), .A2(G244), .A3(new_n286), .A4(new_n282), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G250), .B(G1698), .C1(new_n420), .C2(new_n421), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n580), .A2(new_n387), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n286), .B(new_n583), .C1(new_n420), .C2(new_n421), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n581), .A2(new_n582), .A3(new_n584), .A4(new_n512), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n578), .B1(new_n585), .B2(new_n292), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G179), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n586), .A2(new_n356), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n577), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n586), .A2(G190), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(KEYINPUT78), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT78), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n586), .B2(G190), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n576), .B1(new_n275), .B2(new_n586), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n470), .A2(new_n275), .ZN(new_n598));
  INV_X1    g0398(.A(new_n470), .ZN(new_n599));
  AOI22_X1  g0399(.A1(KEYINPUT85), .A2(new_n598), .B1(new_n599), .B2(new_n305), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n598), .A2(KEYINPUT85), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n496), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n450), .A2(new_n568), .A3(new_n603), .ZN(G372));
  NAND2_X1  g0404(.A1(new_n445), .A2(new_n399), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n372), .A2(new_n377), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n448), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT89), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n344), .A2(KEYINPUT18), .A3(new_n358), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n374), .B1(new_n373), .B2(new_n375), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n359), .A2(new_n376), .A3(KEYINPUT89), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n607), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n613), .A2(new_n309), .B1(new_n273), .B2(new_n312), .ZN(new_n614));
  INV_X1    g0414(.A(new_n586), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G169), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n576), .B1(new_n616), .B2(new_n587), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n592), .A2(new_n594), .ZN(new_n618));
  INV_X1    g0418(.A(new_n596), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n600), .A2(new_n601), .ZN(new_n621));
  INV_X1    g0421(.A(new_n496), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n543), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n552), .B(KEYINPUT86), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n549), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G200), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n558), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n356), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n564), .A2(new_n565), .A3(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n497), .A2(new_n522), .A3(new_n527), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n620), .A2(new_n623), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n562), .A2(KEYINPUT26), .A3(new_n566), .A4(new_n617), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n617), .A2(new_n630), .A3(new_n628), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n634), .A2(KEYINPUT87), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n549), .A2(new_n553), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT80), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n549), .A2(new_n544), .A3(new_n553), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G200), .A3(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n561), .A2(new_n641), .A3(new_n624), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n564), .A2(new_n565), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n642), .A2(new_n559), .B1(new_n643), .B2(new_n563), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT87), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT26), .A4(new_n617), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n637), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT88), .B1(new_n647), .B2(new_n630), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT88), .ZN(new_n649));
  INV_X1    g0449(.A(new_n630), .ZN(new_n650));
  AOI211_X1 g0450(.A(new_n649), .B(new_n650), .C1(new_n637), .C2(new_n646), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n633), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n614), .B1(new_n653), .B2(new_n449), .ZN(G369));
  AND2_X1   g0454(.A1(new_n522), .A2(new_n527), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n530), .ZN(new_n656));
  OR3_X1    g0456(.A1(new_n415), .A2(KEYINPUT27), .A3(G20), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT27), .B1(new_n415), .B2(G20), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT90), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g0463(.A(KEYINPUT91), .B(G343), .Z(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n517), .ZN(new_n667));
  MUX2_X1   g0467(.A(new_n656), .B(new_n655), .S(new_n667), .Z(new_n668));
  INV_X1    g0468(.A(G330), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n622), .A2(new_n666), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n497), .B1(new_n602), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n497), .A2(new_n665), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n655), .A2(new_n665), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n674), .B1(new_n679), .B2(new_n673), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n210), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n533), .A2(new_n390), .A3(new_n507), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(G1), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n216), .B2(new_n684), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n460), .A2(new_n469), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n525), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n639), .A2(new_n640), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n691), .A2(KEYINPUT30), .A3(new_n692), .A4(new_n586), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n524), .A2(G179), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n470), .A3(new_n626), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n693), .B1(new_n586), .B2(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n556), .A2(new_n525), .A3(new_n690), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT30), .B1(new_n697), .B2(new_n586), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n665), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT31), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT92), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n568), .A2(new_n603), .A3(new_n666), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT31), .B(new_n665), .C1(new_n696), .C2(new_n698), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n699), .A2(KEYINPUT92), .A3(new_n700), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n652), .A2(new_n666), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n644), .A2(new_n635), .A3(new_n617), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n650), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n633), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(KEYINPUT29), .A3(new_n666), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n709), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n689), .B1(new_n717), .B2(G1), .ZN(G364));
  NOR2_X1   g0518(.A1(new_n207), .A2(new_n305), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n275), .A2(G179), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G303), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g0523(.A(KEYINPUT33), .B(G317), .Z(new_n724));
  NOR2_X1   g0524(.A1(new_n311), .A2(new_n275), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n207), .A2(G190), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n311), .A2(G200), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G311), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n724), .A2(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n719), .A2(new_n728), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n723), .B(new_n731), .C1(G322), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n719), .A2(new_n725), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G326), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n726), .A2(new_n720), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n726), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(G283), .A2(new_n739), .B1(new_n742), .B2(G329), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n207), .B1(new_n740), .B2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n285), .B1(G294), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n734), .A2(new_n737), .A3(new_n743), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(G159), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT94), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT32), .Z(new_n750));
  NOR2_X1   g0550(.A1(new_n738), .A2(new_n390), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n732), .A2(new_n318), .B1(new_n729), .B2(new_n288), .ZN(new_n752));
  INV_X1    g0552(.A(new_n721), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n751), .B(new_n752), .C1(G87), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n745), .A2(G97), .ZN(new_n755));
  INV_X1    g0555(.A(new_n727), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G50), .A2(new_n736), .B1(new_n756), .B2(G68), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n754), .A2(new_n285), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n747), .B1(new_n750), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n213), .B1(G20), .B2(new_n356), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n682), .A2(new_n333), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n247), .A2(new_n461), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n217), .A2(G45), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G355), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n285), .A2(new_n210), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n765), .B1(G116), .B2(new_n210), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n760), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n252), .A2(G20), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G45), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n684), .A2(G1), .A3(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT93), .Z(new_n777));
  NAND3_X1  g0577(.A1(new_n761), .A2(new_n773), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT95), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n771), .B(KEYINPUT96), .Z(new_n780));
  AOI21_X1  g0580(.A(new_n779), .B1(new_n668), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n776), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n670), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n668), .A2(new_n669), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  NOR2_X1   g0586(.A1(new_n666), .A2(new_n400), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n403), .B1(KEYINPUT98), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n789), .A2(new_n399), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT98), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n787), .B1(new_n399), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n710), .B(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n782), .B1(new_n794), .B2(new_n709), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT99), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n794), .A2(new_n709), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n795), .B2(KEYINPUT99), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n793), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n769), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n760), .A2(new_n769), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT97), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n777), .B1(G77), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n738), .A2(new_n221), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n732), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n729), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n805), .B(new_n807), .C1(new_n485), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n285), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n735), .A2(new_n722), .B1(new_n721), .B2(new_n390), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n727), .A2(new_n812), .B1(new_n741), .B2(new_n730), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n809), .A2(new_n810), .A3(new_n755), .A4(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n736), .A2(G137), .B1(new_n808), .B2(G159), .ZN(new_n816));
  INV_X1    g0616(.A(G143), .ZN(new_n817));
  INV_X1    g0617(.A(G150), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n816), .B1(new_n817), .B2(new_n732), .C1(new_n818), .C2(new_n727), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n721), .A2(new_n202), .B1(new_n741), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n333), .B1(new_n318), .B2(new_n744), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(G68), .C2(new_n739), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n819), .A2(new_n820), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n815), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n804), .B1(new_n760), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n801), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n799), .A2(new_n830), .ZN(G384));
  OAI211_X1 g0631(.A(G116), .B(new_n214), .C1(new_n573), .C2(KEYINPUT35), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(KEYINPUT35), .B2(new_n573), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT36), .ZN(new_n834));
  OR3_X1    g0634(.A1(new_n216), .A2(new_n288), .A3(new_n320), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n202), .A2(G68), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n206), .B(G13), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n712), .A2(new_n450), .A3(new_n716), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n839), .A2(new_n614), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n611), .A2(new_n612), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n663), .B(KEYINPUT101), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n342), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT7), .B1(new_n333), .B2(G20), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n327), .A2(new_n328), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n846), .A2(G68), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n845), .B1(new_n848), .B2(new_n322), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n367), .B1(new_n369), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n663), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n375), .A2(new_n850), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n852), .A3(new_n370), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n373), .A2(new_n375), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n373), .A2(new_n842), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n857), .A2(new_n858), .A3(new_n859), .A4(new_n370), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n378), .A2(new_n853), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT102), .B1(new_n861), .B2(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n378), .A2(new_n853), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n856), .A2(new_n860), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT102), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n861), .A2(KEYINPUT38), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n862), .A2(new_n868), .A3(KEYINPUT39), .A4(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n869), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n857), .A2(new_n858), .A3(new_n370), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n860), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n611), .A2(new_n606), .A3(new_n612), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n858), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n871), .B1(new_n876), .B2(new_n867), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n870), .B1(new_n877), .B2(KEYINPUT39), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n445), .A2(new_n665), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n844), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT100), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n442), .B1(new_n440), .B2(G169), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n435), .A2(new_n311), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n444), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n448), .B(new_n882), .C1(new_n885), .C2(new_n446), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n446), .A2(new_n666), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n445), .A2(new_n882), .A3(new_n448), .A4(new_n887), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n652), .A2(new_n666), .A3(new_n793), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n399), .A2(new_n665), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n891), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n862), .A2(new_n868), .A3(new_n869), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n881), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n840), .B(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n889), .A2(new_n890), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n704), .A2(new_n705), .A3(new_n701), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n899), .A2(new_n793), .A3(new_n896), .A4(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n876), .A2(new_n867), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n902), .B1(new_n903), .B2(new_n869), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n889), .A2(new_n900), .A3(new_n890), .A4(new_n793), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n901), .A2(new_n902), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  AND4_X1   g0707(.A1(new_n445), .A2(new_n405), .A3(new_n448), .A4(new_n900), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n907), .B(new_n908), .Z(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(G330), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n898), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n206), .B2(new_n774), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n898), .A2(new_n910), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n838), .B1(new_n912), .B2(new_n913), .ZN(G367));
  NOR2_X1   g0714(.A1(new_n666), .A2(new_n624), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n630), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n631), .B2(new_n915), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n780), .ZN(new_n918));
  INV_X1    g0718(.A(new_n760), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT46), .B1(new_n753), .B2(new_n485), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n333), .B(new_n920), .C1(G107), .C2(new_n745), .ZN(new_n921));
  XNOR2_X1  g0721(.A(KEYINPUT105), .B(G311), .ZN(new_n922));
  XOR2_X1   g0722(.A(KEYINPUT106), .B(G317), .Z(new_n923));
  OAI22_X1  g0723(.A1(new_n735), .A2(new_n922), .B1(new_n923), .B2(new_n741), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n727), .A2(new_n806), .B1(new_n738), .B2(new_n223), .ZN(new_n925));
  NAND2_X1  g0725(.A1(KEYINPUT46), .A2(G116), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n721), .A2(new_n926), .B1(new_n729), .B2(new_n812), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n732), .A2(new_n722), .ZN(new_n928));
  NOR4_X1   g0728(.A1(new_n924), .A2(new_n925), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(G159), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n735), .A2(new_n817), .B1(new_n727), .B2(new_n930), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n721), .A2(new_n318), .B1(new_n729), .B2(new_n202), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n744), .A2(new_n319), .ZN(new_n933));
  NOR4_X1   g0733(.A1(new_n810), .A2(new_n931), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(KEYINPUT107), .B(G137), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n738), .A2(new_n288), .B1(new_n741), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G150), .B2(new_n733), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n921), .A2(new_n929), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n919), .B1(new_n938), .B2(KEYINPUT47), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(KEYINPUT47), .B2(new_n938), .ZN(new_n940));
  INV_X1    g0740(.A(new_n762), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n772), .B1(new_n210), .B2(new_n380), .C1(new_n243), .C2(new_n941), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n918), .A2(new_n777), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT108), .Z(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n676), .B(new_n679), .Z(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(new_n670), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n717), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n620), .B1(new_n576), .B2(new_n666), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n617), .A2(new_n665), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(new_n680), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT44), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT103), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n951), .B2(new_n680), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(new_n680), .A3(new_n954), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(KEYINPUT45), .A3(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT45), .ZN(new_n959));
  INV_X1    g0759(.A(new_n957), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n960), .B2(new_n955), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n953), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n677), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n678), .A2(new_n958), .A3(new_n961), .A4(new_n953), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n717), .B1(new_n948), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT104), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n683), .B(KEYINPUT41), .Z(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n967), .B1(new_n966), .B2(new_n969), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n775), .A2(G1), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n677), .A2(new_n951), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT43), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n917), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n975), .B(new_n977), .Z(new_n978));
  AND2_X1   g0778(.A1(new_n949), .A2(new_n950), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n679), .A2(new_n673), .A3(new_n675), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT42), .ZN(new_n981));
  OAI21_X1  g0781(.A(KEYINPUT42), .B1(new_n979), .B2(new_n980), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n590), .B1(new_n949), .B2(new_n497), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n666), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n976), .B2(new_n917), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n978), .B(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n945), .B1(new_n974), .B2(new_n987), .ZN(G387));
  INV_X1    g0788(.A(new_n777), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n265), .A2(G50), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT50), .ZN(new_n991));
  AOI211_X1 g0791(.A(G45), .B(new_n685), .C1(G68), .C2(G77), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n941), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT109), .Z(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n239), .B2(new_n461), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(G107), .B2(new_n210), .C1(new_n686), .C2(new_n767), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n989), .B1(new_n996), .B2(new_n772), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n756), .A2(new_n266), .B1(new_n808), .B2(G68), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n223), .B2(new_n738), .C1(new_n930), .C2(new_n735), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G50), .A2(new_n733), .B1(new_n742), .B2(G150), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n288), .B2(new_n721), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n326), .A2(new_n282), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n744), .A2(new_n380), .ZN(new_n1003));
  NOR4_X1   g0803(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n736), .A2(G322), .B1(new_n808), .B2(G303), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n732), .B2(new_n923), .C1(new_n727), .C2(new_n922), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT48), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n753), .A2(G294), .B1(new_n745), .B2(G283), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1006), .A2(new_n1007), .B1(KEYINPUT110), .B2(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(KEYINPUT110), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(new_n1007), .C2(new_n1006), .ZN(new_n1011));
  XOR2_X1   g0811(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n485), .A2(new_n739), .B1(new_n742), .B2(G326), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n1002), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1004), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n997), .B1(new_n919), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n676), .B2(new_n780), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n947), .B2(new_n973), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n948), .A2(new_n683), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n717), .A2(new_n947), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(G393));
  INV_X1    g0823(.A(new_n948), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n965), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n948), .A2(new_n965), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n683), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1025), .A2(new_n973), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n979), .A2(new_n771), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT112), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G317), .A2(new_n736), .B1(new_n733), .B2(G311), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT52), .Z(new_n1033));
  OAI22_X1  g0833(.A1(new_n721), .A2(new_n812), .B1(new_n729), .B2(new_n806), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G303), .B2(new_n756), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n745), .A2(new_n485), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n751), .B(new_n285), .C1(G322), .C2(new_n742), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n735), .A2(new_n818), .B1(new_n732), .B2(new_n930), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT51), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n202), .A2(new_n727), .B1(new_n721), .B2(new_n319), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G143), .B2(new_n742), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n745), .A2(G77), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1002), .B(new_n805), .C1(new_n266), .C2(new_n808), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n919), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n772), .B1(new_n223), .B2(new_n210), .C1(new_n941), .C2(new_n250), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n777), .A2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT113), .Z(new_n1049));
  OR3_X1    g0849(.A1(new_n1031), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1028), .A2(new_n1029), .A3(new_n1050), .ZN(G390));
  NAND2_X1  g0851(.A1(new_n908), .A2(G330), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n839), .A2(new_n1052), .A3(new_n614), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n892), .A2(new_n894), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n891), .B1(new_n708), .B2(new_n800), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n790), .A2(new_n669), .A3(new_n792), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n899), .A2(new_n900), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n889), .A2(new_n890), .A3(new_n793), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n708), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n715), .A2(new_n793), .A3(new_n666), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1063), .A2(new_n894), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n900), .A2(new_n1057), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n891), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1060), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1054), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n878), .B1(new_n895), .B2(new_n879), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1064), .A2(new_n891), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1071), .A2(new_n879), .A3(new_n877), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1062), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n1070), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1058), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1069), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1070), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1067), .A2(new_n1062), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1053), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1055), .A2(new_n899), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n880), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1072), .B1(new_n1083), .B2(new_n878), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1078), .B(new_n1081), .C1(new_n1084), .C2(new_n1058), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1077), .A2(new_n1085), .A3(new_n683), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G283), .A2(new_n736), .B1(new_n733), .B2(G116), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n390), .B2(new_n727), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n810), .B1(new_n221), .B2(new_n721), .C1(new_n223), .C2(new_n729), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G77), .C2(new_n745), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n738), .A2(new_n319), .B1(new_n741), .B2(new_n806), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT115), .Z(new_n1092));
  INV_X1    g0892(.A(G128), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n735), .A2(new_n1093), .B1(new_n732), .B2(new_n822), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT114), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n753), .A2(G150), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT53), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n727), .A2(new_n935), .B1(new_n729), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(G125), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n738), .A2(new_n202), .B1(new_n741), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n285), .B1(new_n930), .B2(new_n744), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1097), .A2(new_n1099), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1090), .A2(new_n1092), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n777), .B1(new_n266), .B2(new_n803), .C1(new_n1104), .C2(new_n919), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n878), .B2(new_n769), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n973), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1086), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT116), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1086), .A2(new_n1108), .A3(KEYINPUT116), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(G378));
  INV_X1    g0913(.A(KEYINPUT118), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1115));
  NAND2_X1  g0915(.A1(new_n273), .A2(new_n851), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n309), .A2(new_n313), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1116), .B1(new_n309), .B2(new_n313), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1115), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1119), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1115), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n907), .A2(new_n1114), .A3(G330), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n904), .A2(new_n906), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n862), .A2(new_n868), .A3(new_n869), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n902), .B1(new_n1127), .B2(new_n905), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1126), .A2(new_n1128), .A3(G330), .A4(new_n1124), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT118), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1124), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n907), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n669), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n897), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1131), .A2(new_n897), .A3(new_n1134), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1132), .A2(new_n769), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n782), .B1(new_n803), .B2(G50), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n333), .A2(G41), .ZN(new_n1142));
  AOI211_X1 g0942(.A(G50), .B(new_n1142), .C1(new_n277), .C2(new_n297), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n729), .A2(new_n380), .B1(new_n741), .B2(new_n812), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1145), .B(new_n1142), .C1(new_n223), .C2(new_n727), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n721), .A2(new_n288), .B1(new_n738), .B2(new_n318), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n735), .A2(new_n507), .B1(new_n732), .B2(new_n390), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1146), .A2(new_n933), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1143), .B1(new_n1149), .B2(KEYINPUT58), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n735), .A2(new_n1100), .B1(new_n727), .B2(new_n822), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n808), .A2(G137), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n1093), .B2(new_n732), .C1(new_n721), .C2(new_n1098), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(G150), .C2(new_n745), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G33), .B(G41), .C1(new_n739), .C2(G159), .ZN(new_n1157));
  INV_X1    g0957(.A(G124), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n741), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT117), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT59), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1160), .B1(new_n1154), .B2(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1150), .B1(KEYINPUT58), .B2(new_n1149), .C1(new_n1156), .C2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1141), .B1(new_n1163), .B2(new_n760), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1139), .A2(new_n973), .B1(new_n1140), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1053), .B1(new_n1107), .B2(new_n1081), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1131), .A2(new_n897), .A3(new_n1134), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n897), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT57), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n683), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1085), .A2(new_n1054), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT57), .B1(new_n1171), .B2(new_n1139), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1165), .B1(new_n1170), .B2(new_n1172), .ZN(G375));
  INV_X1    g0973(.A(new_n803), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n989), .B1(new_n319), .B2(new_n1174), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n333), .B1(new_n318), .B2(new_n738), .C1(new_n727), .C2(new_n1098), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n732), .A2(new_n935), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n735), .A2(new_n822), .B1(new_n729), .B2(new_n818), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n744), .A2(new_n202), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n721), .A2(new_n930), .B1(new_n741), .B2(new_n1093), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT119), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n721), .A2(new_n223), .B1(new_n741), .B2(new_n722), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n485), .B2(new_n756), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n735), .A2(new_n806), .B1(new_n732), .B2(new_n812), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n288), .A2(new_n738), .B1(new_n729), .B2(new_n390), .ZN(new_n1186));
  NOR4_X1   g0986(.A1(new_n1185), .A2(new_n1186), .A3(new_n285), .A4(new_n1003), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1180), .A2(new_n1182), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1175), .B1(new_n919), .B2(new_n1188), .C1(new_n899), .C2(new_n770), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1068), .B2(new_n973), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1081), .A2(new_n968), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1053), .A2(new_n1080), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(G381));
  INV_X1    g0996(.A(G384), .ZN(new_n1197));
  INV_X1    g0997(.A(G390), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(G393), .A2(G396), .ZN(new_n1200));
  NOR4_X1   g1000(.A1(G387), .A2(new_n1199), .A3(G381), .A4(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT120), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1109), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1171), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1085), .A2(new_n1054), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n683), .C1(KEYINPUT57), .C2(new_n1207), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1202), .A2(new_n1203), .A3(new_n1208), .A4(new_n1165), .ZN(G407));
  NAND2_X1  g1009(.A1(new_n1139), .A2(new_n973), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1140), .A2(new_n1164), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1171), .A2(new_n1139), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n1204), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n684), .B1(new_n1205), .B2(new_n1171), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1212), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n664), .A2(G213), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1203), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(G407), .A2(G213), .A3(new_n1219), .ZN(G409));
  OAI21_X1  g1020(.A(new_n1165), .B1(new_n1213), .B2(new_n968), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1203), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1222), .B1(new_n1223), .B2(G375), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1194), .A2(KEYINPUT60), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT60), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1053), .A2(new_n1226), .A3(new_n1080), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n684), .B(new_n1081), .C1(new_n1225), .C2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1197), .B1(new_n1228), .B2(new_n1192), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1228), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(G384), .A3(new_n1191), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1224), .A2(new_n1217), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT62), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1208), .A2(new_n1111), .A3(new_n1112), .A4(new_n1165), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1218), .B1(new_n1236), .B2(new_n1222), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT62), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1233), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1218), .A2(G2897), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1229), .A2(new_n1231), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1207), .A2(new_n969), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1109), .B1(new_n1244), .B2(new_n1165), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G378), .B2(new_n1216), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1243), .B1(new_n1246), .B2(new_n1218), .ZN(new_n1247));
  XOR2_X1   g1047(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1248));
  NAND4_X1  g1048(.A1(new_n1235), .A2(new_n1239), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n972), .A2(new_n973), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n987), .B1(new_n1250), .B2(new_n970), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1198), .B1(new_n1251), .B2(new_n944), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n945), .B(G390), .C1(new_n974), .C2(new_n987), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G393), .B(new_n785), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(KEYINPUT123), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1198), .B1(new_n1254), .B2(KEYINPUT123), .C1(new_n1251), .C2(new_n944), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1251), .A2(new_n944), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(G390), .A3(new_n1254), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT126), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1249), .A2(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1224), .A2(KEYINPUT63), .A3(new_n1217), .A4(new_n1233), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT124), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1237), .A2(new_n1265), .A3(KEYINPUT63), .A4(new_n1233), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1260), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1237), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1269), .B1(new_n1270), .B2(new_n1243), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  XOR2_X1   g1072(.A(KEYINPUT121), .B(KEYINPUT63), .Z(new_n1273));
  AND3_X1   g1073(.A1(new_n1234), .A2(KEYINPUT122), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT122), .B1(new_n1234), .B2(new_n1273), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1262), .B1(new_n1272), .B2(new_n1276), .ZN(G405));
  NOR2_X1   g1077(.A1(new_n1223), .A2(G375), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1216), .A2(new_n1109), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1232), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1236), .B(new_n1233), .C1(new_n1109), .C2(new_n1216), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1260), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1260), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .ZN(G402));
endmodule


