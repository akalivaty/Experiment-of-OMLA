//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G116), .ZN(new_n211));
  INV_X1    g0011(.A(G270), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n214), .B1(new_n202), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n213), .B(new_n218), .C1(G97), .C2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(new_n206), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT64), .B(KEYINPUT1), .Z(new_n222));
  XNOR2_X1  g0022(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n209), .B(new_n223), .C1(new_n226), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n224), .B1(new_n206), .B2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G58), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(new_n216), .ZN(new_n249));
  OR2_X1    g0049(.A1(new_n249), .A2(new_n201), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n250), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT7), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT77), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT76), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n245), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT76), .A2(G33), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n256), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n225), .B(new_n255), .C1(new_n260), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT77), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT7), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n216), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT76), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT76), .A2(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT3), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n261), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n271), .A2(new_n225), .A3(new_n255), .A4(new_n265), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n253), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n247), .B1(new_n273), .B2(KEYINPUT16), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT79), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(KEYINPUT7), .B(new_n225), .C1(new_n278), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n254), .B1(new_n282), .B2(G20), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n216), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n275), .B(new_n277), .C1(new_n284), .C2(new_n253), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n261), .A2(new_n279), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT7), .B1(new_n287), .B2(new_n225), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n258), .A2(new_n256), .A3(new_n259), .ZN(new_n289));
  AOI21_X1  g0089(.A(G20), .B1(new_n289), .B2(new_n279), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n290), .B2(KEYINPUT7), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n252), .B1(new_n291), .B2(new_n216), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n275), .B1(new_n292), .B2(new_n277), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n274), .B1(new_n286), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT80), .ZN(new_n295));
  INV_X1    g0095(.A(G1), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT66), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT66), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n300), .A2(new_n296), .A3(G13), .A4(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT8), .B(G58), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n246), .B1(new_n299), .B2(new_n301), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n305), .A2(new_n297), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n304), .B1(new_n306), .B2(new_n303), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n277), .B1(new_n284), .B2(new_n253), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT79), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n285), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT80), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(new_n274), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n295), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n296), .B1(G41), .B2(G45), .ZN(new_n314));
  INV_X1    g0114(.A(G274), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT65), .B(G1698), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n317), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n318));
  INV_X1    g0118(.A(G87), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n318), .A2(new_n271), .B1(new_n245), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G232), .ZN(new_n323));
  INV_X1    g0123(.A(new_n321), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n314), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n322), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G190), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(G200), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n313), .A2(KEYINPUT17), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT17), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n295), .A2(new_n330), .A3(new_n307), .A4(new_n312), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n328), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n295), .A2(new_n307), .A3(new_n312), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n326), .A2(G169), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n326), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(KEYINPUT18), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT18), .B1(new_n335), .B2(new_n338), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n331), .B(new_n334), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n325), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G244), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G238), .A2(G1698), .ZN(new_n345));
  AND2_X1   g0145(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n282), .B(new_n345), .C1(new_n348), .C2(new_n323), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(new_n321), .C1(G107), .C2(new_n282), .ZN(new_n350));
  INV_X1    g0150(.A(new_n316), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n344), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n352), .A2(new_n327), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n306), .A2(G77), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n245), .A2(G20), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n251), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n355), .A2(new_n357), .B1(new_n303), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G77), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n225), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n246), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n354), .B(new_n362), .C1(G77), .C2(new_n302), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(G200), .B2(new_n352), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n342), .B1(new_n353), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n203), .A2(G20), .ZN(new_n366));
  INV_X1    g0166(.A(G150), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n366), .B1(new_n367), .B2(new_n358), .C1(new_n357), .C2(new_n303), .ZN(new_n368));
  INV_X1    g0168(.A(new_n302), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n368), .A2(new_n246), .B1(new_n202), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n297), .A2(G50), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(KEYINPUT67), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(KEYINPUT67), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n305), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(KEYINPUT9), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT9), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n370), .B2(new_n374), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G223), .A2(G1698), .ZN(new_n380));
  INV_X1    g0180(.A(G222), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n282), .B(new_n380), .C1(new_n348), .C2(new_n381), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n382), .B(new_n321), .C1(G77), .C2(new_n282), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(new_n351), .C1(new_n215), .C2(new_n325), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n327), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT70), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n384), .A2(KEYINPUT69), .A3(G200), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n384), .A2(G200), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT69), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT10), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n386), .A2(new_n387), .A3(new_n388), .A4(new_n391), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n388), .B1(new_n327), .B2(new_n384), .C1(new_n376), .C2(new_n378), .ZN(new_n393));
  INV_X1    g0193(.A(new_n391), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT70), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n386), .A2(new_n389), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n392), .A2(new_n395), .B1(new_n396), .B2(KEYINPUT10), .ZN(new_n397));
  INV_X1    g0197(.A(G169), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n384), .A2(new_n398), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n384), .A2(G179), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n400), .A2(KEYINPUT68), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(KEYINPUT68), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n375), .B(new_n399), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT74), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  OAI21_X1  g0209(.A(G226), .B1(new_n346), .B2(new_n347), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(new_n287), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n261), .A2(new_n279), .A3(G232), .A4(G1698), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT71), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n282), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n411), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n408), .B1(new_n416), .B2(new_n324), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n415), .ZN(new_n418));
  OR2_X1    g0218(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n419));
  NAND2_X1  g0219(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n215), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n282), .B1(G33), .B2(G97), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(KEYINPUT72), .A3(new_n321), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n343), .A2(G238), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n417), .A2(new_n424), .A3(new_n351), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT13), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(new_n321), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n316), .B1(new_n428), .B2(new_n408), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n425), .A4(new_n424), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n407), .B1(new_n432), .B2(new_n398), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n406), .A2(KEYINPUT74), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n398), .B1(new_n427), .B2(new_n431), .ZN(new_n436));
  INV_X1    g0236(.A(new_n407), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n427), .A2(new_n431), .A3(G179), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n433), .A2(new_n435), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n369), .A2(new_n216), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT12), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n356), .A2(G77), .B1(new_n251), .B2(G50), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n225), .B2(G68), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n246), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT11), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n306), .A2(G68), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n442), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT73), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT73), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n442), .A2(new_n446), .A3(new_n450), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT75), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n449), .A2(KEYINPUT75), .A3(new_n451), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n440), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n427), .A2(new_n431), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n452), .B1(new_n459), .B2(new_n327), .ZN(new_n460));
  INV_X1    g0260(.A(G200), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n432), .A2(new_n461), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n352), .A2(new_n398), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n363), .B(new_n464), .C1(G179), .C2(new_n352), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n405), .A2(new_n458), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n365), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n302), .A2(G116), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT87), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n296), .A2(G33), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n305), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G116), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n225), .C1(G33), .C2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n478), .B(new_n246), .C1(new_n225), .C2(G116), .ZN(new_n479));
  XOR2_X1   g0279(.A(new_n479), .B(KEYINPUT20), .Z(new_n480));
  NAND3_X1  g0280(.A1(new_n472), .A2(new_n475), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G45), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(G1), .ZN(new_n484));
  AND2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  NOR2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n324), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G270), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n487), .A2(new_n315), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G264), .A2(G1698), .ZN(new_n492));
  INV_X1    g0292(.A(G257), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n348), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT76), .B(G33), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n262), .B1(new_n495), .B2(KEYINPUT3), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n494), .A2(new_n496), .B1(G303), .B2(new_n287), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n490), .B(new_n491), .C1(new_n497), .C2(new_n324), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G200), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n482), .B(new_n499), .C1(new_n327), .C2(new_n498), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n481), .A2(G169), .A3(new_n498), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT21), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n498), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n481), .A2(G179), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n481), .A2(KEYINPUT21), .A3(G169), .A4(new_n498), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n500), .A2(new_n503), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n324), .A2(new_n487), .A3(G264), .ZN(new_n508));
  OAI21_X1  g0308(.A(G250), .B1(new_n346), .B2(new_n347), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G257), .A2(G1698), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n495), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n496), .A2(new_n511), .B1(G294), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n508), .B(new_n491), .C1(new_n513), .C2(new_n324), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G179), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n398), .B2(new_n514), .ZN(new_n516));
  OR3_X1    g0316(.A1(new_n319), .A2(KEYINPUT22), .A3(G20), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(new_n287), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n270), .A2(new_n225), .A3(G87), .A4(new_n261), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT22), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT88), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT88), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(new_n522), .A3(KEYINPUT22), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n518), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n512), .A2(new_n225), .A3(G116), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n225), .A2(G107), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n526), .B(KEYINPUT23), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT24), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  INV_X1    g0330(.A(new_n528), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n519), .A2(new_n522), .A3(KEYINPUT22), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n522), .B1(new_n519), .B2(KEYINPUT22), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n530), .B(new_n531), .C1(new_n534), .C2(new_n518), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n247), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n369), .A2(KEYINPUT25), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT25), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n302), .B2(G107), .ZN(new_n540));
  AOI22_X1  g0340(.A1(G107), .A2(new_n474), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n516), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT89), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT89), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(new_n516), .C1(new_n536), .C2(new_n542), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n507), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n537), .B1(new_n281), .B2(new_n283), .ZN(new_n548));
  XNOR2_X1  g0348(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n537), .A2(G97), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(G97), .B(G107), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(G20), .C1(new_n552), .C2(new_n549), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n251), .A2(G77), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n246), .B1(new_n548), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT82), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT83), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n302), .A2(new_n477), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n560), .C1(new_n474), .C2(new_n477), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n477), .B1(new_n305), .B2(new_n473), .ZN(new_n562));
  INV_X1    g0362(.A(new_n560), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT83), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(KEYINPUT82), .B(new_n246), .C1(new_n548), .C2(new_n555), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n558), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n270), .A2(G244), .A3(new_n261), .A4(new_n317), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT4), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(KEYINPUT4), .B(G244), .C1(new_n346), .C2(new_n347), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G250), .A2(G1698), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n282), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(new_n476), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n321), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n491), .B1(new_n488), .B2(new_n493), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n398), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n577), .B1(new_n575), .B2(new_n321), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n337), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n567), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT85), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n496), .A2(new_n584), .A3(G244), .A4(G1698), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n270), .A2(G244), .A3(G1698), .A4(new_n261), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT85), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n496), .A2(G238), .A3(new_n317), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n512), .A2(G116), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n585), .A2(new_n587), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n321), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n321), .A2(new_n484), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(G250), .B1(G274), .B2(new_n484), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(G190), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n474), .A2(G87), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT19), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n225), .B1(new_n409), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT86), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n319), .A2(new_n477), .A3(new_n537), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT86), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n600), .B(new_n225), .C1(new_n409), .C2(new_n596), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n270), .A2(new_n225), .A3(G68), .A4(new_n261), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n596), .B1(new_n357), .B2(new_n477), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n246), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n369), .A2(new_n355), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n595), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n593), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n590), .B2(new_n321), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n594), .B(new_n609), .C1(new_n461), .C2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT84), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n579), .B2(new_n327), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n581), .A2(KEYINPUT84), .A3(G190), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n579), .A2(G200), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(new_n565), .A3(new_n566), .A4(new_n558), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n583), .B(new_n612), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n514), .A2(new_n327), .ZN(new_n620));
  INV_X1    g0420(.A(new_n514), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(new_n461), .ZN(new_n622));
  NOR4_X1   g0422(.A1(new_n536), .A2(new_n542), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n355), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n474), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n606), .A2(new_n625), .A3(new_n607), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n611), .B2(G169), .ZN(new_n627));
  AOI211_X1 g0427(.A(G179), .B(new_n610), .C1(new_n590), .C2(new_n321), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n619), .A2(new_n623), .A3(new_n629), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n469), .A2(new_n547), .A3(new_n630), .ZN(G372));
  XNOR2_X1  g0431(.A(new_n543), .B(KEYINPUT90), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n612), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT91), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n583), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n567), .A2(KEYINPUT91), .A3(new_n580), .A4(new_n582), .ZN(new_n638));
  AOI211_X1 g0438(.A(KEYINPUT26), .B(new_n635), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n594), .A2(new_n609), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n611), .A2(new_n461), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n640), .A2(new_n641), .B1(new_n627), .B2(new_n628), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT26), .B1(new_n642), .B2(new_n583), .ZN(new_n643));
  INV_X1    g0443(.A(new_n629), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT92), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n639), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n583), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n644), .A3(new_n612), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n629), .B1(new_n649), .B2(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n637), .A2(new_n638), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(new_n612), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT92), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n634), .B1(new_n647), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n469), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n460), .A2(new_n462), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n458), .B1(new_n657), .B2(new_n465), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n331), .A2(new_n334), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n341), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n339), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n397), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n404), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n656), .A2(new_n665), .ZN(G369));
  AOI21_X1  g0466(.A(new_n623), .B1(new_n544), .B2(new_n546), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n536), .A2(new_n542), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n298), .A2(G20), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n296), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n667), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n675), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n543), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n482), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n633), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n507), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n633), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n675), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n667), .A2(new_n687), .B1(new_n632), .B2(new_n678), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n207), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n599), .A2(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n227), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n646), .B1(new_n639), .B2(new_n645), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n650), .A2(new_n653), .A3(KEYINPUT92), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n675), .B1(new_n699), .B2(new_n634), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n651), .A2(new_n612), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n629), .B1(new_n703), .B2(KEYINPUT26), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n649), .A2(KEYINPUT26), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n619), .A2(new_n623), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n633), .B1(new_n544), .B2(new_n546), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n704), .B(new_n705), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n678), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n702), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n630), .A2(new_n547), .A3(new_n678), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n504), .A2(G179), .ZN(new_n713));
  INV_X1    g0513(.A(new_n611), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT93), .B1(new_n579), .B2(new_n514), .ZN(new_n715));
  INV_X1    g0515(.A(new_n476), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n568), .B2(new_n569), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n324), .B1(new_n717), .B2(new_n574), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n514), .B(KEYINPUT93), .C1(new_n718), .C2(new_n577), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n713), .B(new_n714), .C1(new_n715), .C2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT94), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n611), .A2(new_n581), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n508), .B1(new_n513), .B2(new_n324), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n317), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n728));
  INV_X1    g0528(.A(G303), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n728), .A2(new_n271), .B1(new_n729), .B2(new_n282), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n730), .A2(new_n321), .B1(G270), .B2(new_n489), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n727), .A2(new_n731), .A3(G179), .A4(new_n491), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n724), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n498), .A2(new_n726), .A3(new_n337), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(KEYINPUT30), .A3(new_n611), .A4(new_n581), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT93), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n621), .B2(new_n581), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n611), .B1(new_n738), .B2(new_n719), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(KEYINPUT94), .A3(new_n713), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n723), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n675), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n736), .A2(new_n721), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n712), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n711), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n696), .B1(new_n749), .B2(G1), .ZN(G364));
  NAND2_X1  g0550(.A1(new_n669), .A2(G45), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n692), .A2(G1), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n684), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G330), .B2(new_n682), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n224), .B1(G20), .B2(new_n398), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n496), .A2(new_n690), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G45), .B2(new_n227), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(G45), .B2(new_n240), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n211), .B2(new_n690), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n282), .A2(G355), .A3(new_n207), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n761), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n225), .A2(new_n337), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(new_n327), .A3(G200), .ZN(new_n769));
  XOR2_X1   g0569(.A(KEYINPUT33), .B(G317), .Z(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n768), .A2(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G200), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n225), .B1(new_n776), .B2(G190), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n774), .A2(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n772), .A2(new_n461), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n771), .B(new_n779), .C1(G326), .C2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n768), .A2(new_n327), .A3(new_n461), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G311), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n461), .A2(G179), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(G20), .A3(G190), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n287), .B1(new_n786), .B2(new_n729), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT96), .Z(new_n788));
  NAND3_X1  g0588(.A1(new_n776), .A2(G20), .A3(new_n327), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT97), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n785), .A2(G20), .A3(new_n327), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n791), .A2(G329), .B1(G283), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n781), .A2(new_n784), .A3(new_n788), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n777), .A2(new_n477), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  OAI21_X1  g0597(.A(KEYINPUT32), .B1(new_n789), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n774), .B2(new_n248), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n796), .B(new_n799), .C1(G50), .C2(new_n780), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n793), .A2(G107), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n783), .A2(KEYINPUT95), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n783), .A2(KEYINPUT95), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G77), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n789), .A2(KEYINPUT32), .A3(new_n797), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n786), .A2(new_n319), .ZN(new_n808));
  INV_X1    g0608(.A(new_n769), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n807), .B(new_n808), .C1(G68), .C2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n800), .A2(new_n801), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n795), .B1(new_n811), .B2(new_n287), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n767), .B1(new_n812), .B2(new_n759), .ZN(new_n813));
  INV_X1    g0613(.A(new_n758), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n753), .B(new_n813), .C1(new_n682), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n755), .A2(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n364), .A2(new_n353), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n363), .A2(new_n675), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n465), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n465), .A2(new_n675), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n700), .B(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(new_n748), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n752), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n287), .B1(new_n792), .B2(new_n319), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n791), .B2(G311), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n796), .B1(new_n780), .B2(G303), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(new_n778), .C2(new_n774), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT98), .ZN(new_n831));
  INV_X1    g0631(.A(G283), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n804), .A2(new_n211), .B1(new_n832), .B2(new_n769), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n830), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n834), .B1(new_n831), .B2(new_n833), .C1(new_n537), .C2(new_n786), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G137), .A2(new_n780), .B1(new_n773), .B2(G143), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n836), .B1(new_n367), .B2(new_n769), .C1(new_n804), .C2(new_n797), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT34), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n792), .A2(new_n216), .ZN(new_n841));
  INV_X1    g0641(.A(new_n777), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(G58), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n496), .B1(new_n202), .B2(new_n786), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n791), .B2(G132), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n839), .A2(new_n840), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n835), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n759), .A2(new_n756), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n847), .A2(new_n759), .B1(new_n360), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n823), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n849), .B(new_n753), .C1(new_n850), .C2(new_n757), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n826), .A2(new_n851), .ZN(G384));
  NAND3_X1  g0652(.A1(new_n454), .A2(new_n455), .A3(new_n675), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n439), .B1(new_n436), .B2(new_n437), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n398), .B(new_n407), .C1(new_n427), .C2(new_n431), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n854), .A2(new_n434), .A3(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n463), .B(new_n853), .C1(new_n856), .C2(new_n456), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n457), .B(new_n675), .C1(new_n440), .C2(new_n657), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n712), .A2(new_n744), .A3(new_n860), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n859), .A2(new_n861), .A3(new_n850), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n264), .B(KEYINPUT7), .C1(new_n496), .C2(G20), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(G68), .A3(new_n272), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n252), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT16), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n246), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n273), .A2(new_n276), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n307), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT101), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT101), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n872), .B(new_n307), .C1(new_n868), .C2(new_n869), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n338), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n673), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n871), .A2(new_n875), .A3(new_n873), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n874), .B(new_n876), .C1(new_n333), .C2(new_n328), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n310), .A2(new_n311), .A3(new_n274), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n311), .B1(new_n310), .B2(new_n274), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n881), .A2(new_n329), .A3(new_n330), .A4(new_n307), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n335), .B1(new_n338), .B2(new_n875), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n876), .ZN(new_n886));
  AOI221_X4 g0686(.A(new_n863), .B1(new_n878), .B2(new_n885), .C1(new_n342), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n342), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n878), .A2(new_n885), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n862), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n313), .A2(new_n673), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n342), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n882), .A2(new_n883), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n885), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n862), .B(KEYINPUT40), .C1(new_n887), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n469), .A2(new_n861), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n901), .B(new_n902), .Z(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(G330), .ZN(new_n904));
  INV_X1    g0704(.A(new_n859), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n655), .A2(new_n678), .A3(new_n850), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n906), .B2(new_n822), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n887), .B2(new_n890), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n887), .B2(new_n899), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n876), .B1(new_n659), .B2(new_n662), .ZN(new_n911));
  INV_X1    g0711(.A(new_n889), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n863), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n458), .A2(new_n675), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n910), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n661), .A2(new_n339), .A3(new_n673), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n908), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n665), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n468), .B1(new_n702), .B2(new_n710), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n919), .B(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n904), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n296), .B2(new_n669), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n551), .B1(new_n552), .B2(new_n549), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT35), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(G116), .A3(new_n226), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT99), .Z(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n927), .B2(new_n926), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n249), .A2(new_n227), .A3(new_n360), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT100), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(G50), .B2(new_n216), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(G1), .A3(new_n298), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n925), .A2(new_n932), .A3(new_n936), .ZN(G367));
  NAND2_X1  g0737(.A1(new_n780), .A2(G143), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n797), .B2(new_n769), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n282), .B1(new_n774), .B2(new_n367), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n792), .A2(new_n360), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n805), .A2(G50), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n842), .A2(G68), .ZN(new_n944));
  INV_X1    g0744(.A(G137), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n786), .A2(new_n248), .B1(new_n945), .B2(new_n789), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT106), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n942), .A2(new_n943), .A3(new_n944), .A4(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT107), .Z(new_n949));
  OAI22_X1  g0749(.A1(new_n774), .A2(new_n729), .B1(new_n777), .B2(new_n537), .ZN(new_n950));
  INV_X1    g0750(.A(new_n789), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n496), .B(new_n950), .C1(G317), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n805), .A2(G283), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n793), .A2(G97), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT46), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n786), .A2(new_n955), .A3(new_n211), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n786), .B2(new_n211), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n778), .B2(new_n769), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n956), .B(new_n958), .C1(G311), .C2(new_n780), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n949), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT108), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT47), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n752), .B1(new_n963), .B2(new_n759), .ZN(new_n964));
  INV_X1    g0764(.A(new_n762), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n965), .A2(new_n236), .B1(new_n207), .B2(new_n355), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n964), .B1(new_n761), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT109), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n609), .A2(new_n678), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n629), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n642), .B2(new_n969), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n968), .B1(new_n814), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n616), .A2(new_n618), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(new_n648), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n567), .A2(new_n675), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n583), .B2(new_n678), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT103), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n544), .A2(new_n546), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n583), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n678), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n667), .A2(new_n687), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT42), .B1(new_n983), .B2(new_n976), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n983), .A2(KEYINPUT42), .A3(new_n976), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT104), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n982), .A2(new_n984), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT102), .ZN(new_n992));
  INV_X1    g0792(.A(new_n979), .ZN(new_n993));
  INV_X1    g0793(.A(new_n685), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n994), .A3(new_n992), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n991), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n989), .A2(new_n990), .A3(new_n996), .A4(new_n997), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(new_n1003), .A3(new_n1000), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n751), .A2(G1), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n983), .B1(new_n679), .B2(new_n687), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(new_n684), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n749), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n688), .A2(new_n977), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT45), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n688), .A2(KEYINPUT44), .A3(new_n974), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT44), .B1(new_n688), .B2(new_n974), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OR3_X1    g0814(.A1(new_n1011), .A2(new_n1014), .A3(new_n994), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n994), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n749), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n691), .B(new_n1019), .Z(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1006), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n972), .B1(new_n1005), .B2(new_n1022), .ZN(G387));
  XOR2_X1   g0823(.A(new_n691), .B(KEYINPUT111), .Z(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n749), .B2(new_n1008), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n749), .B2(new_n1008), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n842), .A2(new_n624), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n780), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1027), .B1(new_n303), .B2(new_n769), .C1(new_n1028), .C2(new_n797), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n496), .B1(new_n360), .B2(new_n786), .C1(new_n774), .C2(new_n202), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n954), .B1(new_n367), .B2(new_n789), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n216), .B2(new_n782), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G322), .A2(new_n780), .B1(new_n809), .B2(G311), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n804), .B2(new_n729), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G317), .B2(new_n773), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT48), .Z(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n832), .B2(new_n777), .C1(new_n778), .C2(new_n786), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT49), .Z(new_n1039));
  NAND2_X1  g0839(.A1(new_n951), .A2(G326), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1040), .B(new_n271), .C1(new_n211), .C2(new_n792), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT110), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1033), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1043), .A2(new_n759), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n679), .A2(new_n814), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n762), .B1(new_n233), .B2(new_n483), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n693), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1047), .A2(new_n207), .A3(new_n282), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n216), .A2(new_n360), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n303), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n202), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1047), .B1(new_n1052), .B2(KEYINPUT50), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n483), .C1(KEYINPUT50), .C2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1049), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n690), .A2(new_n537), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n761), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1044), .A2(new_n1045), .A3(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1058), .A2(new_n753), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1026), .A2(new_n1059), .ZN(G393));
  NAND3_X1  g0860(.A1(new_n1015), .A2(new_n1006), .A3(new_n1016), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n760), .B1(new_n477), .B2(new_n207), .C1(new_n965), .C2(new_n243), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G311), .A2(new_n773), .B1(new_n780), .B2(G317), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT52), .Z(new_n1064));
  OAI22_X1  g0864(.A1(new_n778), .A2(new_n782), .B1(new_n769), .B2(new_n729), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n282), .B(new_n1065), .C1(G116), .C2(new_n842), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n786), .A2(new_n832), .B1(new_n775), .B2(new_n789), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT112), .Z(new_n1068));
  NAND4_X1  g0868(.A1(new_n1064), .A2(new_n801), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G150), .A2(new_n780), .B1(new_n773), .B2(G159), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1070), .A2(KEYINPUT51), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n805), .A2(new_n1051), .B1(KEYINPUT51), .B2(new_n1070), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n271), .B1(G50), .B2(new_n809), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n777), .A2(new_n360), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n792), .A2(new_n319), .B1(new_n786), .B2(new_n216), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(G143), .C2(new_n951), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1072), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1069), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n752), .B1(new_n1078), .B2(new_n759), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1062), .B(new_n1079), .C1(new_n993), .C2(new_n814), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1061), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1009), .A2(new_n1017), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n1024), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1009), .A2(new_n1017), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G390));
  NAND2_X1  g0886(.A1(new_n910), .A2(new_n915), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n756), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1074), .B1(new_n773), .B2(G116), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n832), .B2(new_n1028), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n841), .B(new_n1090), .C1(G107), .C2(new_n809), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n282), .B(new_n808), .C1(new_n791), .C2(G294), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(new_n477), .C2(new_n804), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n792), .A2(new_n202), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G128), .A2(new_n780), .B1(new_n773), .B2(G132), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT116), .Z(new_n1096));
  NOR2_X1   g0896(.A1(new_n786), .A2(new_n367), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT53), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n797), .B2(new_n777), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G137), .B2(new_n809), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n282), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G125), .B2(new_n791), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT54), .B(G143), .Z(new_n1104));
  NAND2_X1  g0904(.A1(new_n805), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1096), .A2(new_n1101), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1093), .B1(new_n1094), .B2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1107), .A2(new_n759), .B1(new_n303), .B2(new_n848), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1088), .A2(new_n753), .A3(new_n1108), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n887), .A2(new_n890), .A3(new_n909), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n894), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n659), .B2(new_n662), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n885), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n884), .B1(new_n882), .B2(new_n883), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n863), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT39), .B1(new_n1116), .B2(new_n914), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1110), .A2(new_n1117), .B1(new_n907), .B2(new_n916), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n916), .B1(new_n1116), .B2(new_n914), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n708), .A2(new_n678), .A3(new_n820), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n822), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n859), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n850), .A2(G330), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n859), .A2(new_n747), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n861), .A2(new_n1124), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1125), .B1(new_n1127), .B2(KEYINPUT113), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1118), .A2(new_n1123), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n916), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n821), .B1(new_n700), .B2(new_n850), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n905), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1087), .A2(new_n1133), .B1(new_n1122), .B2(new_n1119), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1127), .A2(new_n859), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(KEYINPUT113), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1130), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1006), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1109), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT117), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AND4_X1   g0942(.A1(G330), .A2(new_n365), .A3(new_n467), .A4(new_n861), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1144), .B(new_n665), .C1(new_n711), .C2(new_n468), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1126), .A2(new_n905), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1147), .A2(new_n822), .A3(new_n1120), .A4(new_n1125), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT115), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n747), .A2(new_n1124), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n905), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1152), .A2(KEYINPUT114), .B1(new_n1127), .B2(new_n859), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1152), .A2(KEYINPUT114), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1132), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1146), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1138), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1148), .B(KEYINPUT115), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1132), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1145), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n1136), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1130), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1024), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1157), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(KEYINPUT117), .B(new_n1109), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1142), .A2(new_n1167), .A3(new_n1168), .ZN(G378));
  XNOR2_X1  g0969(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n397), .A2(KEYINPUT55), .A3(new_n404), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(KEYINPUT55), .B1(new_n397), .B2(new_n404), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n375), .A2(new_n875), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1171), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1174), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n375), .B(new_n875), .C1(new_n1179), .C2(new_n1172), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1170), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1178), .A2(new_n1182), .A3(new_n756), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n848), .A2(new_n202), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G125), .A2(new_n780), .B1(new_n773), .B2(G128), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G132), .B2(new_n809), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n786), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1188), .A2(new_n1104), .B1(new_n842), .B2(G150), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(new_n945), .C2(new_n782), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n951), .A2(G124), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(G33), .A2(G41), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT118), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G159), .B2(new_n793), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n496), .A2(G41), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n793), .A2(G58), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1199), .B(new_n944), .C1(new_n360), .C2(new_n786), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(G283), .C2(new_n791), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n809), .A2(G97), .B1(new_n783), .B2(new_n624), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n211), .B2(new_n1028), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1201), .B(new_n1204), .C1(new_n537), .C2(new_n774), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT58), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1198), .A2(new_n202), .A3(new_n1195), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1197), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n752), .B1(new_n1208), .B2(new_n759), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1183), .A2(new_n1184), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n859), .A2(new_n861), .A3(new_n850), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n913), .B2(new_n914), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n900), .B(G330), .C1(new_n1212), .C2(KEYINPUT40), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT120), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1178), .A2(new_n1182), .A3(KEYINPUT120), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1213), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1178), .A2(new_n1182), .A3(KEYINPUT120), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1219), .A2(new_n893), .A3(G330), .A4(new_n900), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1218), .A2(new_n919), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n919), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1210), .B1(new_n1223), .B2(new_n1139), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n919), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1218), .A2(new_n919), .A3(new_n1220), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1146), .B1(new_n1138), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1024), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1229), .A2(new_n1231), .A3(KEYINPUT57), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1224), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(G375));
  OAI221_X1 g1037(.A(new_n1027), .B1(new_n1028), .B2(new_n778), .C1(new_n832), .C2(new_n774), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n790), .A2(new_n729), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n287), .B1(new_n786), .B2(new_n477), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n941), .A4(new_n1240), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n537), .B2(new_n804), .C1(new_n211), .C2(new_n769), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT121), .Z(new_n1243));
  NOR2_X1   g1043(.A1(new_n777), .A2(new_n202), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n773), .A2(G137), .B1(new_n809), .B2(new_n1104), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n780), .A2(G132), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n367), .C2(new_n782), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1244), .B(new_n1247), .C1(G128), .C2(new_n791), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1199), .A2(new_n496), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT122), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1248), .B(new_n1250), .C1(new_n797), .C2(new_n786), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1243), .A2(new_n1251), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT123), .Z(new_n1253));
  AOI21_X1  g1053(.A(new_n752), .B1(new_n1253), .B2(new_n759), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n757), .B2(new_n859), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n216), .B2(new_n848), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1230), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1257), .B2(new_n1006), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1158), .A2(new_n1161), .A3(new_n1145), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1156), .A2(new_n1021), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(G381));
  AOI221_X4 g1061(.A(new_n1128), .B1(new_n1119), .B2(new_n1122), .C1(new_n1087), .C2(new_n1133), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1137), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1145), .B1(new_n1264), .B2(new_n1257), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1233), .B1(new_n1265), .B2(new_n1223), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(new_n1166), .A3(new_n1235), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1142), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1224), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1085), .B(new_n972), .C1(new_n1005), .C2(new_n1022), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1272), .A2(G384), .A3(G381), .ZN(new_n1273));
  OR2_X1    g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1271), .A2(new_n1273), .A3(new_n1275), .ZN(G407));
  OAI211_X1 g1076(.A(G407), .B(G213), .C1(G343), .C2(new_n1270), .ZN(G409));
  NAND2_X1  g1077(.A1(G387), .A2(G390), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1272), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n1274), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1274), .A2(new_n1280), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1278), .A2(new_n1272), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1268), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1230), .A2(KEYINPUT60), .A3(new_n1145), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT60), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1259), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1286), .A2(new_n1288), .A3(new_n1166), .A4(new_n1156), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(G384), .A3(new_n1258), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT125), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1258), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n826), .A3(new_n851), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1289), .A2(new_n1294), .A3(G384), .A4(new_n1258), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1291), .A2(new_n1293), .A3(KEYINPUT62), .A4(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1229), .A2(new_n1231), .A3(new_n1021), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(G378), .A2(new_n1298), .A3(new_n1224), .ZN(new_n1299));
  INV_X1    g1099(.A(G213), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1300), .A2(G343), .ZN(new_n1301));
  NOR4_X1   g1101(.A1(new_n1285), .A2(new_n1296), .A3(new_n1299), .A4(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT124), .B1(new_n1285), .B2(new_n1299), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1301), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT124), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1268), .A2(new_n1269), .A3(new_n1297), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1305), .B(new_n1306), .C1(new_n1236), .C2(new_n1268), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1291), .A2(new_n1293), .A3(new_n1295), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1303), .A2(new_n1304), .A3(new_n1307), .A4(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1302), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT61), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1301), .A2(G2897), .ZN(new_n1314));
  OR2_X1    g1114(.A1(new_n1314), .A2(KEYINPUT127), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1291), .A2(new_n1293), .A3(new_n1315), .A4(new_n1295), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(KEYINPUT127), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1316), .B(new_n1317), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1285), .A2(new_n1299), .A3(new_n1301), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1313), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1284), .B1(new_n1312), .B2(new_n1320), .ZN(new_n1321));
  XOR2_X1   g1121(.A(new_n1316), .B(new_n1317), .Z(new_n1322));
  NAND3_X1  g1122(.A1(new_n1303), .A2(new_n1304), .A3(new_n1307), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT61), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1309), .A2(KEYINPUT63), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1284), .B1(new_n1319), .B2(new_n1325), .ZN(new_n1326));
  XOR2_X1   g1126(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1327));
  NAND2_X1  g1127(.A1(new_n1310), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1324), .A2(new_n1326), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1321), .A2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(new_n1284), .A2(new_n1309), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1281), .A2(new_n1308), .A3(new_n1283), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1271), .A2(new_n1285), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1333), .B(new_n1334), .ZN(G402));
endmodule


