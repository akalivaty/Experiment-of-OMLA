

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n702), .A2(n923), .ZN(n696) );
  BUF_X1 U549 ( .A(n875), .Z(n517) );
  XOR2_X1 U550 ( .A(KEYINPUT17), .B(n540), .Z(n875) );
  NAND2_X1 U551 ( .A1(n765), .A2(n763), .ZN(n709) );
  AND2_X1 U552 ( .A1(n730), .A2(n725), .ZN(n724) );
  INV_X1 U553 ( .A(G2105), .ZN(n536) );
  XNOR2_X1 U554 ( .A(n526), .B(KEYINPUT70), .ZN(n527) );
  XOR2_X1 U555 ( .A(G543), .B(KEYINPUT0), .Z(n518) );
  NOR2_X1 U556 ( .A1(n709), .A2(n944), .ZN(n692) );
  XNOR2_X1 U557 ( .A(n706), .B(KEYINPUT27), .ZN(n707) );
  XNOR2_X1 U558 ( .A(n708), .B(n707), .ZN(n711) );
  XNOR2_X1 U559 ( .A(n723), .B(KEYINPUT94), .ZN(n731) );
  NOR2_X1 U560 ( .A1(n733), .A2(n732), .ZN(n736) );
  AND2_X1 U561 ( .A1(n742), .A2(n741), .ZN(n743) );
  INV_X1 U562 ( .A(KEYINPUT9), .ZN(n526) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n540) );
  NAND2_X1 U564 ( .A1(n808), .A2(n795), .ZN(n796) );
  XNOR2_X1 U565 ( .A(n528), .B(n527), .ZN(n529) );
  NOR2_X1 U566 ( .A1(n522), .A2(n630), .ZN(n635) );
  OR2_X1 U567 ( .A1(n797), .A2(n796), .ZN(n814) );
  NOR2_X1 U568 ( .A1(G651), .A2(n630), .ZN(n640) );
  OR2_X1 U569 ( .A1(n548), .A2(n547), .ZN(n550) );
  INV_X1 U570 ( .A(G651), .ZN(n522) );
  NOR2_X1 U571 ( .A1(G543), .A2(n522), .ZN(n520) );
  XNOR2_X1 U572 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n519) );
  XNOR2_X1 U573 ( .A(n520), .B(n519), .ZN(n639) );
  NAND2_X1 U574 ( .A1(n639), .A2(G64), .ZN(n521) );
  XNOR2_X1 U575 ( .A(KEYINPUT69), .B(n521), .ZN(n530) );
  XNOR2_X1 U576 ( .A(KEYINPUT66), .B(n518), .ZN(n630) );
  NAND2_X1 U577 ( .A1(n635), .A2(G77), .ZN(n525) );
  NOR2_X1 U578 ( .A1(G543), .A2(G651), .ZN(n523) );
  XNOR2_X1 U579 ( .A(n523), .B(KEYINPUT64), .ZN(n636) );
  NAND2_X1 U580 ( .A1(G90), .A2(n636), .ZN(n524) );
  NAND2_X1 U581 ( .A1(n525), .A2(n524), .ZN(n528) );
  NOR2_X1 U582 ( .A1(n530), .A2(n529), .ZN(n532) );
  NAND2_X1 U583 ( .A1(n640), .A2(G52), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U585 ( .A(KEYINPUT71), .B(n533), .Z(G301) );
  NOR2_X1 U586 ( .A1(G2104), .A2(n536), .ZN(n879) );
  NAND2_X1 U587 ( .A1(G125), .A2(n879), .ZN(n535) );
  AND2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n882) );
  NAND2_X1 U589 ( .A1(G113), .A2(n882), .ZN(n534) );
  AND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n673) );
  INV_X1 U591 ( .A(KEYINPUT23), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n536), .A2(G2104), .ZN(n537) );
  XNOR2_X2 U593 ( .A(n537), .B(KEYINPUT65), .ZN(n873) );
  NAND2_X1 U594 ( .A1(G101), .A2(n873), .ZN(n538) );
  XNOR2_X1 U595 ( .A(n539), .B(n538), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n517), .A2(G137), .ZN(n541) );
  AND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n674) );
  AND2_X1 U598 ( .A1(n673), .A2(n674), .ZN(G160) );
  INV_X1 U599 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U600 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U601 ( .A1(G138), .A2(n875), .ZN(n544) );
  NAND2_X1 U602 ( .A1(G126), .A2(n879), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U604 ( .A1(G114), .A2(n882), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G102), .A2(n873), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n547) );
  INV_X1 U607 ( .A(KEYINPUT82), .ZN(n549) );
  XNOR2_X1 U608 ( .A(n550), .B(n549), .ZN(n672) );
  BUF_X1 U609 ( .A(n672), .Z(G164) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  NAND2_X1 U612 ( .A1(G63), .A2(n639), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G51), .A2(n640), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U615 ( .A(KEYINPUT6), .B(n553), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G89), .A2(n636), .ZN(n554) );
  XNOR2_X1 U617 ( .A(n554), .B(KEYINPUT4), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G76), .A2(n635), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U620 ( .A(n557), .B(KEYINPUT5), .Z(n558) );
  NOR2_X1 U621 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT75), .B(n560), .Z(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT7), .B(n561), .Z(G168) );
  XOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U627 ( .A(G223), .ZN(n816) );
  NAND2_X1 U628 ( .A1(n816), .A2(G567), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U630 ( .A1(G81), .A2(n636), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G68), .A2(n635), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT13), .B(n567), .Z(n571) );
  NAND2_X1 U635 ( .A1(G56), .A2(n639), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(KEYINPUT14), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(KEYINPUT73), .ZN(n570) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n640), .A2(G43), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n920) );
  INV_X1 U641 ( .A(G860), .ZN(n823) );
  NOR2_X1 U642 ( .A1(n920), .A2(n823), .ZN(n574) );
  XOR2_X1 U643 ( .A(KEYINPUT74), .B(n574), .Z(G153) );
  NAND2_X1 U644 ( .A1(G868), .A2(G301), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G66), .A2(n639), .ZN(n576) );
  NAND2_X1 U646 ( .A1(G54), .A2(n640), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n635), .A2(G79), .ZN(n578) );
  NAND2_X1 U649 ( .A1(G92), .A2(n636), .ZN(n577) );
  NAND2_X1 U650 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U652 ( .A(n581), .B(KEYINPUT15), .ZN(n923) );
  INV_X1 U653 ( .A(G868), .ZN(n652) );
  NAND2_X1 U654 ( .A1(n923), .A2(n652), .ZN(n582) );
  NAND2_X1 U655 ( .A1(n583), .A2(n582), .ZN(G284) );
  NAND2_X1 U656 ( .A1(G65), .A2(n639), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G53), .A2(n640), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n635), .A2(G78), .ZN(n587) );
  NAND2_X1 U660 ( .A1(G91), .A2(n636), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n913) );
  XOR2_X1 U663 ( .A(n913), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U664 ( .A1(G299), .A2(G868), .ZN(n591) );
  NOR2_X1 U665 ( .A1(G286), .A2(n652), .ZN(n590) );
  NOR2_X1 U666 ( .A1(n591), .A2(n590), .ZN(G297) );
  NAND2_X1 U667 ( .A1(n823), .A2(G559), .ZN(n592) );
  INV_X1 U668 ( .A(n923), .ZN(n633) );
  NAND2_X1 U669 ( .A1(n592), .A2(n633), .ZN(n593) );
  XNOR2_X1 U670 ( .A(n593), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U671 ( .A1(n633), .A2(G868), .ZN(n594) );
  NOR2_X1 U672 ( .A1(G559), .A2(n594), .ZN(n595) );
  XNOR2_X1 U673 ( .A(n595), .B(KEYINPUT76), .ZN(n597) );
  NOR2_X1 U674 ( .A1(n920), .A2(G868), .ZN(n596) );
  NOR2_X1 U675 ( .A1(n597), .A2(n596), .ZN(G282) );
  NAND2_X1 U676 ( .A1(n879), .A2(G123), .ZN(n598) );
  XNOR2_X1 U677 ( .A(n598), .B(KEYINPUT18), .ZN(n600) );
  NAND2_X1 U678 ( .A1(G111), .A2(n882), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U680 ( .A1(G135), .A2(n517), .ZN(n602) );
  NAND2_X1 U681 ( .A1(G99), .A2(n873), .ZN(n601) );
  NAND2_X1 U682 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U683 ( .A1(n604), .A2(n603), .ZN(n975) );
  XNOR2_X1 U684 ( .A(n975), .B(G2096), .ZN(n606) );
  INV_X1 U685 ( .A(G2100), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n606), .A2(n605), .ZN(G156) );
  NAND2_X1 U687 ( .A1(n639), .A2(G61), .ZN(n608) );
  NAND2_X1 U688 ( .A1(G86), .A2(n636), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n635), .A2(G73), .ZN(n609) );
  XOR2_X1 U691 ( .A(KEYINPUT2), .B(n609), .Z(n610) );
  NOR2_X1 U692 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n640), .A2(G48), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(G305) );
  NAND2_X1 U695 ( .A1(n635), .A2(G75), .ZN(n615) );
  NAND2_X1 U696 ( .A1(G88), .A2(n636), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G62), .A2(n639), .ZN(n617) );
  NAND2_X1 U699 ( .A1(G50), .A2(n640), .ZN(n616) );
  NAND2_X1 U700 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U701 ( .A1(n619), .A2(n618), .ZN(G166) );
  NAND2_X1 U702 ( .A1(n635), .A2(G72), .ZN(n621) );
  NAND2_X1 U703 ( .A1(G85), .A2(n636), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G60), .A2(n639), .ZN(n623) );
  NAND2_X1 U706 ( .A1(G47), .A2(n640), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U708 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U709 ( .A(KEYINPUT68), .B(n626), .Z(G290) );
  NAND2_X1 U710 ( .A1(G49), .A2(n640), .ZN(n628) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U713 ( .A1(n639), .A2(n629), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G87), .A2(n630), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U716 ( .A1(G559), .A2(n633), .ZN(n634) );
  XOR2_X1 U717 ( .A(n920), .B(n634), .Z(n822) );
  NAND2_X1 U718 ( .A1(n635), .A2(G80), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G93), .A2(n636), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G67), .A2(n639), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G55), .A2(n640), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U725 ( .A(KEYINPUT77), .B(n645), .ZN(n824) );
  XOR2_X1 U726 ( .A(G299), .B(n824), .Z(n647) );
  XNOR2_X1 U727 ( .A(G305), .B(G166), .ZN(n646) );
  XNOR2_X1 U728 ( .A(n647), .B(n646), .ZN(n650) );
  XNOR2_X1 U729 ( .A(G290), .B(KEYINPUT19), .ZN(n648) );
  XNOR2_X1 U730 ( .A(n648), .B(G288), .ZN(n649) );
  XNOR2_X1 U731 ( .A(n650), .B(n649), .ZN(n891) );
  XNOR2_X1 U732 ( .A(n822), .B(n891), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n651), .A2(G868), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n652), .A2(n824), .ZN(n653) );
  NAND2_X1 U735 ( .A1(n654), .A2(n653), .ZN(G295) );
  XOR2_X1 U736 ( .A(KEYINPUT78), .B(KEYINPUT20), .Z(n656) );
  NAND2_X1 U737 ( .A1(G2078), .A2(G2084), .ZN(n655) );
  XNOR2_X1 U738 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n657), .ZN(n658) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n658), .ZN(n659) );
  NAND2_X1 U741 ( .A1(n659), .A2(G2072), .ZN(G158) );
  NAND2_X1 U742 ( .A1(G120), .A2(G108), .ZN(n660) );
  NOR2_X1 U743 ( .A1(G237), .A2(n660), .ZN(n661) );
  NAND2_X1 U744 ( .A1(n661), .A2(G69), .ZN(n662) );
  XNOR2_X1 U745 ( .A(n662), .B(KEYINPUT80), .ZN(n820) );
  NAND2_X1 U746 ( .A1(n820), .A2(G567), .ZN(n663) );
  XNOR2_X1 U747 ( .A(n663), .B(KEYINPUT81), .ZN(n669) );
  NAND2_X1 U748 ( .A1(G132), .A2(G82), .ZN(n664) );
  XNOR2_X1 U749 ( .A(n664), .B(KEYINPUT79), .ZN(n665) );
  XNOR2_X1 U750 ( .A(KEYINPUT22), .B(n665), .ZN(n666) );
  NAND2_X1 U751 ( .A1(n666), .A2(G96), .ZN(n667) );
  OR2_X1 U752 ( .A1(G218), .A2(n667), .ZN(n821) );
  AND2_X1 U753 ( .A1(G2106), .A2(n821), .ZN(n668) );
  NOR2_X1 U754 ( .A1(n669), .A2(n668), .ZN(G319) );
  INV_X1 U755 ( .A(G319), .ZN(n671) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n670) );
  NOR2_X1 U757 ( .A1(n671), .A2(n670), .ZN(n819) );
  NAND2_X1 U758 ( .A1(n819), .A2(G36), .ZN(G176) );
  INV_X1 U759 ( .A(G166), .ZN(G303) );
  NOR2_X1 U760 ( .A1(G1384), .A2(n672), .ZN(n765) );
  AND2_X1 U761 ( .A1(n673), .A2(G40), .ZN(n675) );
  AND2_X1 U762 ( .A1(n675), .A2(n674), .ZN(n763) );
  NAND2_X1 U763 ( .A1(G8), .A2(n709), .ZN(n758) );
  NOR2_X1 U764 ( .A1(G1966), .A2(n758), .ZN(n733) );
  NOR2_X1 U765 ( .A1(G2084), .A2(n709), .ZN(n734) );
  NOR2_X1 U766 ( .A1(n733), .A2(n734), .ZN(n676) );
  NAND2_X1 U767 ( .A1(G8), .A2(n676), .ZN(n677) );
  XNOR2_X1 U768 ( .A(KEYINPUT30), .B(n677), .ZN(n678) );
  NOR2_X1 U769 ( .A1(G168), .A2(n678), .ZN(n683) );
  XOR2_X1 U770 ( .A(KEYINPUT88), .B(G1961), .Z(n998) );
  NAND2_X1 U771 ( .A1(n998), .A2(n709), .ZN(n680) );
  INV_X1 U772 ( .A(n709), .ZN(n705) );
  XNOR2_X1 U773 ( .A(G2078), .B(KEYINPUT25), .ZN(n945) );
  NAND2_X1 U774 ( .A1(n705), .A2(n945), .ZN(n679) );
  NAND2_X1 U775 ( .A1(n680), .A2(n679), .ZN(n720) );
  INV_X1 U776 ( .A(n720), .ZN(n681) );
  AND2_X1 U777 ( .A1(G301), .A2(n681), .ZN(n682) );
  NOR2_X1 U778 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U779 ( .A(n684), .B(KEYINPUT31), .ZN(n685) );
  XNOR2_X1 U780 ( .A(n685), .B(KEYINPUT95), .ZN(n730) );
  INV_X1 U781 ( .A(G8), .ZN(n691) );
  NOR2_X1 U782 ( .A1(G2090), .A2(n709), .ZN(n686) );
  XNOR2_X1 U783 ( .A(n686), .B(KEYINPUT96), .ZN(n688) );
  NOR2_X1 U784 ( .A1(n758), .A2(G1971), .ZN(n687) );
  NOR2_X1 U785 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U786 ( .A1(n689), .A2(G303), .ZN(n690) );
  OR2_X1 U787 ( .A1(n691), .A2(n690), .ZN(n725) );
  XOR2_X1 U788 ( .A(G1996), .B(KEYINPUT90), .Z(n944) );
  XNOR2_X1 U789 ( .A(n692), .B(KEYINPUT26), .ZN(n693) );
  NOR2_X1 U790 ( .A1(n920), .A2(n693), .ZN(n695) );
  NAND2_X1 U791 ( .A1(G1341), .A2(n709), .ZN(n694) );
  NAND2_X1 U792 ( .A1(n695), .A2(n694), .ZN(n702) );
  XNOR2_X1 U793 ( .A(n696), .B(KEYINPUT91), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n709), .A2(G1348), .ZN(n697) );
  XNOR2_X1 U795 ( .A(n697), .B(KEYINPUT92), .ZN(n699) );
  NAND2_X1 U796 ( .A1(n705), .A2(G2067), .ZN(n698) );
  NAND2_X1 U797 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U798 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U799 ( .A1(n923), .A2(n702), .ZN(n703) );
  NAND2_X1 U800 ( .A1(n704), .A2(n703), .ZN(n713) );
  NAND2_X1 U801 ( .A1(G2072), .A2(n705), .ZN(n708) );
  INV_X1 U802 ( .A(KEYINPUT89), .ZN(n706) );
  AND2_X1 U803 ( .A1(n709), .A2(G1956), .ZN(n710) );
  NOR2_X1 U804 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U805 ( .A1(n913), .A2(n714), .ZN(n712) );
  NAND2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U807 ( .A1(n913), .A2(n714), .ZN(n715) );
  XOR2_X1 U808 ( .A(n715), .B(KEYINPUT28), .Z(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n719) );
  XNOR2_X1 U810 ( .A(KEYINPUT29), .B(KEYINPUT93), .ZN(n718) );
  XNOR2_X1 U811 ( .A(n719), .B(n718), .ZN(n722) );
  NAND2_X1 U812 ( .A1(G171), .A2(n720), .ZN(n721) );
  NAND2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n724), .A2(n731), .ZN(n728) );
  INV_X1 U815 ( .A(n725), .ZN(n726) );
  OR2_X1 U816 ( .A1(n726), .A2(G286), .ZN(n727) );
  NAND2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U818 ( .A(n729), .B(KEYINPUT32), .ZN(n738) );
  AND2_X1 U819 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U820 ( .A1(G8), .A2(n734), .ZN(n735) );
  NAND2_X1 U821 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U822 ( .A1(n738), .A2(n737), .ZN(n752) );
  NOR2_X1 U823 ( .A1(G1976), .A2(G288), .ZN(n744) );
  NOR2_X1 U824 ( .A1(G1971), .A2(G303), .ZN(n739) );
  NOR2_X1 U825 ( .A1(n744), .A2(n739), .ZN(n917) );
  NAND2_X1 U826 ( .A1(n752), .A2(n917), .ZN(n742) );
  INV_X1 U827 ( .A(n758), .ZN(n740) );
  NAND2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n916) );
  AND2_X1 U829 ( .A1(n740), .A2(n916), .ZN(n741) );
  NOR2_X1 U830 ( .A1(KEYINPUT33), .A2(n743), .ZN(n747) );
  NAND2_X1 U831 ( .A1(n744), .A2(KEYINPUT33), .ZN(n745) );
  NOR2_X1 U832 ( .A1(n745), .A2(n758), .ZN(n746) );
  NOR2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n749) );
  XNOR2_X1 U834 ( .A(KEYINPUT97), .B(G1981), .ZN(n748) );
  XNOR2_X1 U835 ( .A(n748), .B(G305), .ZN(n932) );
  NAND2_X1 U836 ( .A1(n749), .A2(n932), .ZN(n755) );
  NOR2_X1 U837 ( .A1(G2090), .A2(G303), .ZN(n750) );
  NAND2_X1 U838 ( .A1(G8), .A2(n750), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U840 ( .A1(n753), .A2(n758), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n761) );
  NOR2_X1 U842 ( .A1(G1981), .A2(G305), .ZN(n756) );
  XOR2_X1 U843 ( .A(n756), .B(KEYINPUT24), .Z(n757) );
  NOR2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U845 ( .A(KEYINPUT87), .B(n759), .Z(n760) );
  NOR2_X1 U846 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U847 ( .A(n762), .B(KEYINPUT98), .ZN(n797) );
  INV_X1 U848 ( .A(n763), .ZN(n764) );
  NOR2_X1 U849 ( .A1(n765), .A2(n764), .ZN(n811) );
  NAND2_X1 U850 ( .A1(n517), .A2(G140), .ZN(n766) );
  XOR2_X1 U851 ( .A(KEYINPUT83), .B(n766), .Z(n768) );
  NAND2_X1 U852 ( .A1(n873), .A2(G104), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U854 ( .A(KEYINPUT34), .B(n769), .ZN(n775) );
  NAND2_X1 U855 ( .A1(G128), .A2(n879), .ZN(n771) );
  NAND2_X1 U856 ( .A1(G116), .A2(n882), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U858 ( .A(KEYINPUT84), .B(n772), .Z(n773) );
  XNOR2_X1 U859 ( .A(KEYINPUT35), .B(n773), .ZN(n774) );
  NOR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U861 ( .A(KEYINPUT36), .B(n776), .ZN(n887) );
  XNOR2_X1 U862 ( .A(KEYINPUT37), .B(G2067), .ZN(n798) );
  NOR2_X1 U863 ( .A1(n887), .A2(n798), .ZN(n982) );
  NAND2_X1 U864 ( .A1(n811), .A2(n982), .ZN(n777) );
  XOR2_X1 U865 ( .A(KEYINPUT85), .B(n777), .Z(n808) );
  NAND2_X1 U866 ( .A1(G129), .A2(n879), .ZN(n779) );
  NAND2_X1 U867 ( .A1(G117), .A2(n882), .ZN(n778) );
  NAND2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n873), .A2(G105), .ZN(n780) );
  XOR2_X1 U870 ( .A(KEYINPUT38), .B(n780), .Z(n781) );
  NOR2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n517), .A2(G141), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n870) );
  NAND2_X1 U874 ( .A1(G1996), .A2(n870), .ZN(n785) );
  XOR2_X1 U875 ( .A(KEYINPUT86), .B(n785), .Z(n793) );
  NAND2_X1 U876 ( .A1(G119), .A2(n879), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G131), .A2(n517), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G107), .A2(n882), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G95), .A2(n873), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n869) );
  INV_X1 U883 ( .A(G1991), .ZN(n800) );
  NOR2_X1 U884 ( .A1(n869), .A2(n800), .ZN(n792) );
  NOR2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n803) );
  XOR2_X1 U886 ( .A(G1986), .B(G290), .Z(n922) );
  NAND2_X1 U887 ( .A1(n803), .A2(n922), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n794), .A2(n811), .ZN(n795) );
  AND2_X1 U889 ( .A1(n887), .A2(n798), .ZN(n799) );
  XNOR2_X1 U890 ( .A(KEYINPUT101), .B(n799), .ZN(n987) );
  NOR2_X1 U891 ( .A1(G1996), .A2(n870), .ZN(n972) );
  AND2_X1 U892 ( .A1(n800), .A2(n869), .ZN(n976) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n801) );
  XOR2_X1 U894 ( .A(n801), .B(KEYINPUT99), .Z(n802) );
  NOR2_X1 U895 ( .A1(n976), .A2(n802), .ZN(n804) );
  INV_X1 U896 ( .A(n803), .ZN(n978) );
  NOR2_X1 U897 ( .A1(n804), .A2(n978), .ZN(n805) );
  NOR2_X1 U898 ( .A1(n972), .A2(n805), .ZN(n806) );
  XNOR2_X1 U899 ( .A(KEYINPUT39), .B(n806), .ZN(n807) );
  XNOR2_X1 U900 ( .A(n807), .B(KEYINPUT100), .ZN(n809) );
  NAND2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n987), .A2(n810), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U905 ( .A(n815), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U907 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U908 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(G188) );
  XNOR2_X1 U911 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  INV_X1 U913 ( .A(G132), .ZN(G219) );
  INV_X1 U914 ( .A(G120), .ZN(G236) );
  INV_X1 U915 ( .A(G96), .ZN(G221) );
  INV_X1 U916 ( .A(G82), .ZN(G220) );
  NOR2_X1 U917 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U918 ( .A(G325), .ZN(G261) );
  NAND2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n825) );
  XNOR2_X1 U920 ( .A(n825), .B(n824), .ZN(G145) );
  XOR2_X1 U921 ( .A(KEYINPUT42), .B(G2072), .Z(n827) );
  XNOR2_X1 U922 ( .A(G2084), .B(G2078), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U924 ( .A(n828), .B(G2100), .Z(n830) );
  XNOR2_X1 U925 ( .A(G2067), .B(G2090), .ZN(n829) );
  XNOR2_X1 U926 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U927 ( .A(G2096), .B(KEYINPUT43), .Z(n832) );
  XNOR2_X1 U928 ( .A(G2678), .B(KEYINPUT103), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U930 ( .A(n834), .B(n833), .Z(G227) );
  XOR2_X1 U931 ( .A(G1956), .B(G1971), .Z(n836) );
  XNOR2_X1 U932 ( .A(G1986), .B(G1976), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U934 ( .A(n837), .B(G2474), .Z(n839) );
  XNOR2_X1 U935 ( .A(G1996), .B(G1991), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U937 ( .A(KEYINPUT41), .B(G1961), .Z(n841) );
  XNOR2_X1 U938 ( .A(G1981), .B(G1966), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(G229) );
  NAND2_X1 U941 ( .A1(G124), .A2(n879), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n844), .B(KEYINPUT44), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n845), .B(KEYINPUT104), .ZN(n847) );
  NAND2_X1 U944 ( .A1(G136), .A2(n517), .ZN(n846) );
  NAND2_X1 U945 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n848), .B(KEYINPUT105), .ZN(n850) );
  NAND2_X1 U947 ( .A1(G112), .A2(n882), .ZN(n849) );
  NAND2_X1 U948 ( .A1(n850), .A2(n849), .ZN(n853) );
  NAND2_X1 U949 ( .A1(n873), .A2(G100), .ZN(n851) );
  XOR2_X1 U950 ( .A(KEYINPUT106), .B(n851), .Z(n852) );
  NOR2_X1 U951 ( .A1(n853), .A2(n852), .ZN(G162) );
  NAND2_X1 U952 ( .A1(G139), .A2(n517), .ZN(n855) );
  NAND2_X1 U953 ( .A1(G103), .A2(n873), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n862) );
  NAND2_X1 U955 ( .A1(n879), .A2(G127), .ZN(n856) );
  XNOR2_X1 U956 ( .A(KEYINPUT109), .B(n856), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n882), .A2(G115), .ZN(n857) );
  XOR2_X1 U958 ( .A(KEYINPUT110), .B(n857), .Z(n858) );
  NOR2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n860), .B(KEYINPUT47), .ZN(n861) );
  NOR2_X1 U961 ( .A1(n862), .A2(n861), .ZN(n966) );
  XOR2_X1 U962 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n864) );
  XNOR2_X1 U963 ( .A(n975), .B(KEYINPUT46), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U965 ( .A(G162), .B(n865), .ZN(n867) );
  XNOR2_X1 U966 ( .A(G164), .B(G160), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n966), .B(n868), .ZN(n872) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n872), .B(n871), .ZN(n889) );
  NAND2_X1 U971 ( .A1(n873), .A2(G106), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n874), .B(KEYINPUT108), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G142), .A2(n517), .ZN(n876) );
  NAND2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U975 ( .A(n878), .B(KEYINPUT45), .ZN(n881) );
  NAND2_X1 U976 ( .A1(G130), .A2(n879), .ZN(n880) );
  NAND2_X1 U977 ( .A1(n881), .A2(n880), .ZN(n885) );
  NAND2_X1 U978 ( .A1(G118), .A2(n882), .ZN(n883) );
  XNOR2_X1 U979 ( .A(KEYINPUT107), .B(n883), .ZN(n884) );
  NOR2_X1 U980 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U981 ( .A(n887), .B(n886), .Z(n888) );
  XNOR2_X1 U982 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U983 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U984 ( .A(n891), .B(KEYINPUT112), .ZN(n893) );
  XNOR2_X1 U985 ( .A(n923), .B(G286), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n893), .B(n892), .ZN(n895) );
  XOR2_X1 U987 ( .A(n920), .B(G171), .Z(n894) );
  XNOR2_X1 U988 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U989 ( .A1(G37), .A2(n896), .ZN(G397) );
  XOR2_X1 U990 ( .A(G2438), .B(G2435), .Z(n898) );
  XNOR2_X1 U991 ( .A(G2443), .B(KEYINPUT102), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U993 ( .A(n899), .B(G2454), .Z(n901) );
  XNOR2_X1 U994 ( .A(G1348), .B(G1341), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U996 ( .A(G2451), .B(G2427), .Z(n903) );
  XNOR2_X1 U997 ( .A(G2430), .B(G2446), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U999 ( .A(n905), .B(n904), .Z(n906) );
  NAND2_X1 U1000 ( .A1(G14), .A2(n906), .ZN(n912) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n912), .ZN(n909) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(n909), .A2(n908), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G69), .ZN(G235) );
  INV_X1 U1009 ( .A(n912), .ZN(G401) );
  XOR2_X1 U1010 ( .A(G16), .B(KEYINPUT56), .Z(n939) );
  XNOR2_X1 U1011 ( .A(G1956), .B(n913), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(G1971), .A2(G303), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n931) );
  XOR2_X1 U1016 ( .A(G1341), .B(n920), .Z(n921) );
  NAND2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n929) );
  XNOR2_X1 U1018 ( .A(G1348), .B(KEYINPUT120), .ZN(n924) );
  XNOR2_X1 U1019 ( .A(n924), .B(n923), .ZN(n926) );
  XNOR2_X1 U1020 ( .A(G1961), .B(G301), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(n927), .B(KEYINPUT121), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n936) );
  XNOR2_X1 U1025 ( .A(G1966), .B(G168), .ZN(n933) );
  NAND2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1027 ( .A(KEYINPUT57), .B(n934), .Z(n935) );
  NOR2_X1 U1028 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1029 ( .A(KEYINPUT122), .B(n937), .ZN(n938) );
  NOR2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n965) );
  XOR2_X1 U1031 ( .A(G2090), .B(G35), .Z(n943) );
  XOR2_X1 U1032 ( .A(G2084), .B(G34), .Z(n940) );
  XNOR2_X1 U1033 ( .A(KEYINPUT118), .B(n940), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n941), .B(KEYINPUT54), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n959) );
  XOR2_X1 U1036 ( .A(n944), .B(G32), .Z(n947) );
  XOR2_X1 U1037 ( .A(n945), .B(G27), .Z(n946) );
  NOR2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n955) );
  XNOR2_X1 U1039 ( .A(G2067), .B(G26), .ZN(n949) );
  XNOR2_X1 U1040 ( .A(G1991), .B(G25), .ZN(n948) );
  NOR2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1042 ( .A1(G28), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(KEYINPUT116), .B(G2072), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(G33), .B(n951), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(n956), .B(KEYINPUT117), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(n957), .B(KEYINPUT53), .ZN(n958) );
  NOR2_X1 U1049 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1050 ( .A(KEYINPUT119), .B(n960), .Z(n961) );
  NOR2_X1 U1051 ( .A1(G29), .A2(n961), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(KEYINPUT55), .B(n962), .ZN(n963) );
  NAND2_X1 U1053 ( .A1(n963), .A2(G11), .ZN(n964) );
  NOR2_X1 U1054 ( .A1(n965), .A2(n964), .ZN(n992) );
  XNOR2_X1 U1055 ( .A(G164), .B(G2078), .ZN(n969) );
  XOR2_X1 U1056 ( .A(G2072), .B(n966), .Z(n967) );
  XNOR2_X1 U1057 ( .A(KEYINPUT115), .B(n967), .ZN(n968) );
  NAND2_X1 U1058 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1059 ( .A(n970), .B(KEYINPUT50), .ZN(n986) );
  XOR2_X1 U1060 ( .A(G2090), .B(G162), .Z(n971) );
  NOR2_X1 U1061 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1062 ( .A(KEYINPUT51), .B(n973), .Z(n974) );
  XNOR2_X1 U1063 ( .A(KEYINPUT114), .B(n974), .ZN(n984) );
  NOR2_X1 U1064 ( .A1(n976), .A2(n975), .ZN(n980) );
  XOR2_X1 U1065 ( .A(G160), .B(G2084), .Z(n977) );
  NOR2_X1 U1066 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1067 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1068 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1069 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1070 ( .A1(n986), .A2(n985), .ZN(n988) );
  NAND2_X1 U1071 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1072 ( .A(KEYINPUT52), .B(n989), .ZN(n990) );
  NAND2_X1 U1073 ( .A1(n990), .A2(G29), .ZN(n991) );
  NAND2_X1 U1074 ( .A1(n992), .A2(n991), .ZN(n1021) );
  XOR2_X1 U1075 ( .A(G1976), .B(G23), .Z(n994) );
  XOR2_X1 U1076 ( .A(G1971), .B(G22), .Z(n993) );
  NAND2_X1 U1077 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1078 ( .A(G24), .B(G1986), .ZN(n995) );
  NOR2_X1 U1079 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1080 ( .A(KEYINPUT58), .B(n997), .Z(n1017) );
  XOR2_X1 U1081 ( .A(G1966), .B(G21), .Z(n1000) );
  XNOR2_X1 U1082 ( .A(G5), .B(n998), .ZN(n999) );
  NAND2_X1 U1083 ( .A1(n1000), .A2(n999), .ZN(n1014) );
  XOR2_X1 U1084 ( .A(G1981), .B(G6), .Z(n1003) );
  XNOR2_X1 U1085 ( .A(KEYINPUT123), .B(G20), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(n1001), .B(G1956), .ZN(n1002) );
  NAND2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1088 ( .A(G19), .B(G1341), .ZN(n1004) );
  NOR2_X1 U1089 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(KEYINPUT124), .B(n1006), .ZN(n1010) );
  XOR2_X1 U1091 ( .A(KEYINPUT125), .B(G4), .Z(n1008) );
  XNOR2_X1 U1092 ( .A(G1348), .B(KEYINPUT59), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(n1008), .B(n1007), .ZN(n1009) );
  NAND2_X1 U1094 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(n1011), .B(KEYINPUT60), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(n1012), .B(KEYINPUT126), .ZN(n1013) );
  NOR2_X1 U1097 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(KEYINPUT127), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1099 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1100 ( .A(KEYINPUT61), .B(n1018), .Z(n1019) );
  NOR2_X1 U1101 ( .A1(G16), .A2(n1019), .ZN(n1020) );
  NOR2_X1 U1102 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1103 ( .A(n1022), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

