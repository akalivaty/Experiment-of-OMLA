//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT64), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n454), .A2(G567), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT65), .Z(new_n461));
  NOR2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT66), .Z(G319));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI211_X1 g048(.A(KEYINPUT67), .B(G2105), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n466), .A2(new_n468), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n477), .A2(new_n472), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n477), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n482), .A2(KEYINPUT68), .A3(G124), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n485), .A2(new_n487), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NOR2_X1   g067(.A1(new_n465), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G102), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(new_n465), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT3), .B(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n494), .B1(new_n498), .B2(new_n472), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT69), .A2(G138), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n466), .A2(new_n468), .A3(new_n500), .A4(new_n472), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n497), .A2(KEYINPUT4), .A3(new_n472), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n499), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n513), .B2(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT70), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G75), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n507), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n514), .A2(G88), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n516), .A2(G62), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n518), .A2(new_n525), .ZN(G166));
  AND2_X1   g101(.A1(new_n519), .A2(new_n521), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT71), .Z(new_n529));
  NAND2_X1  g104(.A1(new_n514), .A2(new_n527), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  INV_X1    g107(.A(new_n509), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT6), .ZN(new_n534));
  OAI211_X1 g109(.A(G543), .B(new_n533), .C1(new_n516), .C2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n529), .A2(new_n532), .A3(new_n537), .A4(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  NAND2_X1  g116(.A1(new_n531), .A2(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n536), .A2(G52), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n513), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n531), .A2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n522), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n536), .A2(G43), .B1(new_n516), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT72), .B1(new_n535), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n514), .A2(new_n563), .A3(G53), .A4(G543), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n564), .A3(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n514), .A2(G91), .A3(new_n527), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n522), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  OAI211_X1 g147(.A(KEYINPUT72), .B(new_n572), .C1(new_n535), .C2(new_n561), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n565), .A2(new_n571), .A3(new_n573), .ZN(G299));
  NAND2_X1  g149(.A1(G171), .A2(KEYINPUT73), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n546), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G301));
  OR2_X1    g153(.A1(new_n518), .A2(new_n525), .ZN(G303));
  OAI21_X1  g154(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n580));
  INV_X1    g155(.A(G49), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  OAI221_X1 g157(.A(new_n580), .B1(new_n581), .B2(new_n535), .C1(new_n530), .C2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n584), .A2(G86), .A3(new_n533), .A4(new_n527), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n584), .A2(G48), .A3(G543), .A4(new_n533), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n519), .A2(new_n521), .A3(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT74), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n519), .A2(new_n521), .A3(new_n591), .A4(G61), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(new_n516), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n587), .A2(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n522), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(new_n516), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(KEYINPUT75), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n531), .A2(G85), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n536), .A2(G47), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n599), .A2(KEYINPUT75), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n600), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n530), .A2(KEYINPUT10), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n522), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n536), .A2(G54), .B1(G651), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT10), .B1(new_n530), .B2(new_n606), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n607), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT76), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n605), .B1(G868), .B2(new_n615), .ZN(G284));
  OAI21_X1  g191(.A(new_n605), .B1(G868), .B2(new_n615), .ZN(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G299), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G168), .B2(new_n618), .ZN(G280));
  XNOR2_X1  g195(.A(G280), .B(KEYINPUT77), .ZN(G297));
  XNOR2_X1  g196(.A(KEYINPUT78), .B(G559), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n615), .B1(G860), .B2(new_n623), .ZN(G148));
  NAND2_X1  g199(.A1(new_n615), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n482), .A2(G123), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n486), .A2(G135), .ZN(new_n630));
  NOR2_X1   g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(new_n472), .B2(G111), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n635));
  NOR3_X1   g210(.A1(new_n467), .A2(new_n465), .A3(G2105), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT80), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT13), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n634), .B(new_n641), .C1(KEYINPUT80), .C2(new_n638), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2435), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2438), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT81), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  XOR2_X1   g234(.A(G2067), .B(G2678), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n659), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n638), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n661), .A2(new_n662), .ZN(new_n668));
  AOI21_X1  g243(.A(KEYINPUT18), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n680), .A2(new_n672), .A3(new_n675), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n678), .B(new_n681), .C1(new_n672), .C2(new_n680), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n682), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT83), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT84), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(G229));
  NAND2_X1  g265(.A1(new_n482), .A2(G119), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n486), .A2(G131), .ZN(new_n692));
  NOR2_X1   g267(.A1(G95), .A2(G2105), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(new_n472), .B2(G107), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n691), .B(new_n692), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(G25), .B(new_n695), .S(G29), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT35), .B(G1991), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  NOR2_X1   g273(.A1(G16), .A2(G24), .ZN(new_n699));
  INV_X1    g274(.A(G290), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(G16), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT85), .B(G1986), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(G16), .A2(G23), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(G288), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT33), .ZN(new_n707));
  INV_X1    g282(.A(G1976), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(G303), .A2(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(G22), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT87), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n710), .A2(new_n714), .A3(new_n711), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n713), .A2(G1971), .A3(new_n715), .ZN(new_n719));
  MUX2_X1   g294(.A(G6), .B(G305), .S(G16), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT32), .B(G1981), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT86), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n709), .A2(new_n718), .A3(new_n719), .A4(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT34), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n698), .B(new_n703), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n728), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G33), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n493), .A2(G103), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  AOI22_X1  g313(.A1(new_n497), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n486), .A2(G139), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n740), .A2(KEYINPUT91), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(KEYINPUT91), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n738), .B1(new_n472), .B2(new_n739), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT92), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n736), .B1(new_n744), .B2(new_n735), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT93), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2072), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n724), .B(new_n725), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n748), .A2(new_n731), .A3(new_n698), .A4(new_n703), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n705), .A2(G4), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n615), .B2(new_n705), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(G1348), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n705), .A2(G19), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n554), .B2(new_n705), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G1341), .Z(new_n755));
  XOR2_X1   g330(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n735), .A2(G26), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n482), .A2(G128), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n486), .A2(G140), .ZN(new_n760));
  OR2_X1    g335(.A1(G104), .A2(G2105), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n758), .B1(new_n764), .B2(new_n735), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n751), .A2(G1348), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n752), .A2(new_n755), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT90), .ZN(new_n770));
  NAND2_X1  g345(.A1(G299), .A2(G16), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n705), .A2(KEYINPUT23), .A3(G20), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT23), .ZN(new_n773));
  INV_X1    g348(.A(G20), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(G16), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n771), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G1956), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(G168), .A2(G16), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G16), .B2(G21), .ZN(new_n780));
  INV_X1    g355(.A(G1966), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT24), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(G34), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(G29), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G160), .B2(new_n735), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G2084), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n778), .A2(new_n782), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G27), .A2(G29), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G164), .B2(G29), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G2078), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n705), .A2(G5), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G171), .B2(new_n705), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1961), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n789), .A2(G2084), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n793), .A2(G2078), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n633), .A2(new_n735), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(G28), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(G28), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n802), .A2(new_n803), .A3(new_n735), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n798), .A2(new_n799), .A3(new_n800), .A4(new_n804), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n791), .A2(new_n794), .A3(new_n797), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT31), .B(G11), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n806), .B(new_n807), .C1(new_n781), .C2(new_n780), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n770), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n734), .A2(new_n747), .A3(new_n749), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n486), .A2(G141), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT94), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n493), .A2(G105), .ZN(new_n813));
  NAND3_X1  g388(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT26), .ZN(new_n815));
  AOI211_X1 g390(.A(new_n813), .B(new_n815), .C1(G129), .C2(new_n482), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G29), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G29), .B2(G32), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT27), .B(G1996), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n735), .A2(G35), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G162), .B2(new_n735), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT29), .B(G2090), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n810), .A2(new_n822), .A3(new_n826), .ZN(G311));
  AND3_X1   g402(.A1(new_n734), .A2(new_n749), .A3(new_n809), .ZN(new_n828));
  INV_X1    g403(.A(new_n822), .ZN(new_n829));
  INV_X1    g404(.A(new_n826), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n828), .A2(new_n829), .A3(new_n830), .A4(new_n747), .ZN(G150));
  NAND2_X1  g406(.A1(new_n536), .A2(G55), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT95), .B(G93), .Z(new_n834));
  OAI221_X1 g409(.A(new_n832), .B1(new_n513), .B2(new_n833), .C1(new_n530), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT96), .B(KEYINPUT37), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n835), .B(new_n553), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n615), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n838), .B1(new_n843), .B2(G860), .ZN(G145));
  XNOR2_X1  g419(.A(new_n817), .B(new_n695), .ZN(new_n845));
  XNOR2_X1  g420(.A(G164), .B(new_n637), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n744), .A2(new_n763), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT92), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n743), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n764), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n482), .A2(G130), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n486), .A2(G142), .ZN(new_n854));
  OR2_X1    g429(.A1(G106), .A2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n849), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n849), .B2(new_n852), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n848), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n849), .A2(new_n852), .ZN(new_n861));
  INV_X1    g436(.A(new_n857), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n849), .A2(new_n852), .A3(new_n857), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n864), .A3(new_n847), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G160), .B(new_n633), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G162), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(G37), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n860), .A2(new_n865), .A3(new_n868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT97), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n860), .A2(new_n865), .A3(new_n873), .A4(new_n868), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT98), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n870), .A2(new_n872), .A3(new_n877), .A4(new_n874), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n876), .A2(KEYINPUT40), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT40), .B1(new_n876), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(G395));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n882));
  INV_X1    g457(.A(G288), .ZN(new_n883));
  NAND2_X1  g458(.A1(G290), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(G290), .A2(new_n883), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT100), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G166), .B(G305), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n700), .A2(G288), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n891), .A3(new_n884), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n888), .A2(new_n891), .A3(new_n884), .A4(new_n890), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n893), .A2(KEYINPUT101), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT101), .B1(new_n893), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT42), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n894), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n882), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n839), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n625), .B(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n613), .A2(G299), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n613), .A2(G299), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n906), .A2(KEYINPUT41), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(KEYINPUT41), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(KEYINPUT99), .A3(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(KEYINPUT99), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n625), .B(new_n839), .ZN(new_n912));
  INV_X1    g487(.A(new_n906), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n900), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(KEYINPUT102), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n901), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n898), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n893), .A2(KEYINPUT101), .A3(new_n894), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n899), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT102), .B1(new_n923), .B2(new_n917), .ZN(new_n924));
  INV_X1    g499(.A(new_n918), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n835), .A2(new_n618), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(G295));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n930), .A3(new_n928), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n916), .B1(new_n901), .B2(new_n918), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n924), .A2(new_n915), .A3(new_n925), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n618), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n928), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT103), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n936), .ZN(G331));
  NAND2_X1  g512(.A1(G286), .A2(G171), .ZN(new_n938));
  INV_X1    g513(.A(G301), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n839), .B(new_n938), .C1(new_n939), .C2(G286), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  AOI21_X1  g516(.A(G286), .B1(new_n575), .B2(new_n577), .ZN(new_n942));
  INV_X1    g517(.A(new_n938), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n902), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n902), .B(KEYINPUT105), .C1(new_n942), .C2(new_n943), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n945), .A2(new_n909), .A3(new_n910), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n921), .A2(new_n922), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n940), .A2(new_n913), .A3(new_n944), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n948), .B1(new_n947), .B2(new_n949), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n906), .B1(new_n945), .B2(new_n946), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n940), .A2(new_n944), .B1(new_n907), .B2(new_n908), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n950), .B(new_n951), .C1(new_n957), .C2(new_n948), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n954), .B1(KEYINPUT43), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n952), .A2(new_n953), .ZN(new_n963));
  OAI211_X1 g538(.A(KEYINPUT44), .B(new_n962), .C1(new_n963), .C2(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(G397));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n499), .B2(new_n505), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n497), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT67), .B1(new_n970), .B2(G2105), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n471), .A2(new_n464), .A3(new_n472), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(G40), .A3(new_n480), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G2078), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT45), .B(new_n966), .C1(new_n499), .C2(new_n505), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n969), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n505), .ZN(new_n980));
  INV_X1    g555(.A(G126), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n477), .A2(new_n981), .B1(new_n495), .B2(new_n465), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n982), .A2(G2105), .B1(G102), .B2(new_n493), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n974), .ZN(new_n988));
  INV_X1    g563(.A(G1961), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n977), .A2(new_n978), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n979), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G171), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT123), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n979), .A2(G301), .A3(new_n990), .A4(new_n991), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT123), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(new_n996), .A3(G171), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n994), .A2(KEYINPUT54), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT122), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n969), .A2(new_n974), .A3(new_n976), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n781), .ZN(new_n1001));
  INV_X1    g576(.A(G2084), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n986), .A2(new_n987), .A3(new_n974), .A4(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(G168), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n1005));
  AND2_X1   g580(.A1(KEYINPUT121), .A2(G8), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1005), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(G8), .A3(G286), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n999), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT51), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1015));
  AND4_X1   g590(.A1(new_n999), .A2(new_n1014), .A3(new_n1011), .A4(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n998), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n992), .A2(new_n939), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n995), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n973), .A2(new_n967), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n708), .B2(G288), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n883), .B2(G1976), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  AND4_X1   g605(.A1(new_n1030), .A2(new_n594), .A3(new_n585), .A4(new_n586), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n587), .B2(new_n594), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT112), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT112), .B(new_n1035), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1024), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1034), .A2(KEYINPUT113), .A3(new_n1024), .A4(new_n1036), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n1028), .B(new_n1029), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1000), .A2(new_n717), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT109), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n988), .B2(G2090), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT109), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1000), .A2(new_n1046), .A3(new_n717), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n973), .B1(KEYINPUT50), .B2(new_n967), .ZN(new_n1048));
  INV_X1    g623(.A(G2090), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1048), .A2(KEYINPUT111), .A3(new_n1049), .A4(new_n986), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G303), .A2(G8), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1052), .B(KEYINPUT55), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1051), .A2(new_n1054), .A3(G8), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n475), .A2(G40), .A3(new_n480), .A4(new_n985), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(KEYINPUT115), .C1(new_n973), .C2(new_n967), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n974), .B(new_n1058), .C1(new_n984), .C2(new_n985), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1057), .A2(new_n1059), .A3(new_n1049), .A4(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1061), .A2(new_n1042), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1053), .B1(new_n1062), .B2(new_n1023), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1021), .A2(new_n1041), .A3(new_n1055), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT124), .B1(new_n1017), .B2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT56), .B(G2072), .Z(new_n1066));
  NOR2_X1   g641(.A1(new_n1000), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1057), .A2(new_n1060), .A3(new_n1059), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n777), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n1070));
  INV_X1    g645(.A(new_n565), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n573), .A2(new_n566), .A3(new_n570), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n565), .A2(new_n571), .A3(KEYINPUT57), .A4(new_n573), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT120), .B1(new_n1069), .B2(new_n1076), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1067), .B(new_n1075), .C1(new_n1068), .C2(new_n777), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1068), .A2(new_n777), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1067), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1076), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1077), .A2(KEYINPUT61), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1075), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT61), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1069), .A2(new_n1076), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1084), .A2(KEYINPUT120), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT58), .B(G1341), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n1000), .A2(G1996), .B1(new_n1022), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n554), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT59), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1092), .A2(new_n1095), .A3(new_n554), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n973), .A2(new_n967), .A3(G2067), .ZN(new_n1098));
  INV_X1    g673(.A(G1348), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n988), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n615), .B2(KEYINPUT60), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n615), .A2(KEYINPUT60), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1101), .B(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1088), .A2(new_n1097), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n613), .A2(KEYINPUT76), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n613), .A2(KEYINPUT76), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1105), .B1(new_n1108), .B2(new_n1100), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1348), .B1(new_n1048), .B2(new_n986), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n615), .B(KEYINPUT117), .C1(new_n1110), .C2(new_n1098), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1109), .B(new_n1111), .C1(new_n1076), .C2(new_n1069), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n1086), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1113), .B1(new_n1112), .B2(new_n1086), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1104), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1029), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1028), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n1055), .A3(new_n1063), .A4(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT54), .B1(new_n1018), .B2(new_n995), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1009), .A2(new_n999), .A3(new_n1011), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1014), .A2(new_n1015), .A3(new_n1011), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT122), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1122), .A2(new_n1123), .A3(new_n1127), .A4(new_n998), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1065), .A2(new_n1117), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1055), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1041), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n883), .A2(new_n708), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1024), .B1(new_n1133), .B2(new_n1031), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT114), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT114), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1131), .A2(new_n1134), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1010), .A2(G8), .A3(G168), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT116), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1051), .A2(G8), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(new_n1053), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1141), .A2(new_n1041), .A3(new_n1055), .A4(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1142), .B1(new_n1120), .B2(new_n1140), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1136), .A2(new_n1138), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT62), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1124), .A2(new_n1126), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1127), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1120), .A2(new_n1018), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1129), .A2(new_n1147), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n969), .A2(new_n973), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(G1996), .A3(new_n817), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT107), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n763), .B(new_n766), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(G1996), .B2(new_n817), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1157), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1160), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n695), .B(new_n697), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT108), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1167), .A2(new_n1157), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(G1986), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n700), .A2(new_n1157), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1157), .A2(G1986), .A3(G290), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT106), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1169), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1156), .A2(new_n1175), .ZN(new_n1176));
  OR3_X1    g751(.A1(new_n969), .A2(G1996), .A3(new_n973), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT46), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT127), .Z(new_n1180));
  NAND2_X1  g755(.A1(new_n818), .A2(new_n1161), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1157), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT126), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1180), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT47), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n695), .A2(new_n697), .ZN(new_n1187));
  OAI22_X1  g762(.A1(new_n1165), .A2(new_n1187), .B1(G2067), .B2(new_n763), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1157), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1171), .B(KEYINPUT48), .Z(new_n1190));
  OAI211_X1 g765(.A(new_n1186), .B(new_n1189), .C1(new_n1169), .C2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1176), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g768(.A(G227), .B1(new_n655), .B2(new_n657), .ZN(new_n1195));
  AND2_X1   g769(.A1(new_n875), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g770(.A(G229), .ZN(new_n1197));
  NAND4_X1  g771(.A1(new_n959), .A2(new_n1196), .A3(new_n462), .A4(new_n1197), .ZN(G225));
  INV_X1    g772(.A(G225), .ZN(G308));
endmodule


