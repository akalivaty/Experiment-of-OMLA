//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(new_n466), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(new_n471), .B2(KEYINPUT3), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n472), .A2(KEYINPUT67), .A3(G137), .A4(new_n461), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT3), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n467), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n476), .A2(G137), .A3(new_n461), .A4(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n469), .A2(new_n461), .A3(new_n470), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT68), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n469), .A2(new_n484), .A3(new_n461), .A4(new_n470), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT69), .B1(new_n486), .B2(G101), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  INV_X1    g063(.A(G101), .ZN(new_n489));
  AOI211_X1 g064(.A(new_n488), .B(new_n489), .C1(new_n483), .C2(new_n485), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n481), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n481), .B(KEYINPUT70), .C1(new_n487), .C2(new_n490), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n465), .B1(new_n493), .B2(new_n494), .ZN(G160));
  NAND2_X1  g070(.A1(new_n472), .A2(new_n461), .ZN(new_n496));
  INV_X1    g071(.A(G136), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n461), .A2(G112), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n496), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n476), .A2(G2105), .A3(new_n477), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(G124), .B2(new_n501), .ZN(new_n502));
  XOR2_X1   g077(.A(new_n502), .B(KEYINPUT71), .Z(G162));
  NAND4_X1  g078(.A1(new_n476), .A2(G138), .A3(new_n461), .A4(new_n477), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g082(.A(G138), .B(new_n461), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(new_n462), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n476), .A2(G126), .A3(G2105), .A4(new_n477), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n461), .B2(G114), .ZN(new_n514));
  INV_X1    g089(.A(G114), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT72), .A3(G2105), .ZN(new_n516));
  OR2_X1    g091(.A1(G102), .A2(G2105), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n514), .A2(new_n516), .A3(new_n517), .A4(G2104), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(G164));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT5), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n528), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT6), .B(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G88), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G50), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n531), .A2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  XNOR2_X1  g114(.A(new_n527), .B(KEYINPUT74), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n540), .A2(G63), .A3(G651), .ZN(new_n541));
  INV_X1    g116(.A(new_n533), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G89), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n532), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G51), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n541), .A2(new_n543), .A3(new_n545), .A4(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  AOI22_X1  g124(.A1(new_n540), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n530), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n542), .A2(G90), .B1(G52), .B2(new_n546), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(G171));
  AOI22_X1  g128(.A1(new_n540), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n530), .ZN(new_n555));
  XNOR2_X1  g130(.A(KEYINPUT75), .B(G43), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n542), .A2(G81), .B1(new_n546), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(new_n546), .A2(G53), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT9), .Z(new_n567));
  AOI22_X1  g142(.A1(new_n528), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n568), .A2(new_n530), .B1(new_n533), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  OAI21_X1  g148(.A(G651), .B1(new_n540), .B2(G74), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT77), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n546), .A2(G49), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n542), .A2(G87), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT76), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(G288));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n527), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n580), .B1(new_n583), .B2(G651), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n580), .A3(G651), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n585), .A2(new_n586), .B1(G48), .B2(new_n546), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n542), .A2(G86), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n542), .A2(G85), .B1(G47), .B2(new_n546), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n540), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n530), .ZN(G290));
  AND3_X1   g167(.A1(new_n528), .A2(G92), .A3(new_n532), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT10), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n528), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(new_n530), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n546), .A2(KEYINPUT79), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n546), .A2(KEYINPUT79), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n597), .A2(G54), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n594), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G284));
  OAI21_X1  g178(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n571), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n571), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(new_n600), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n486), .A2(new_n462), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT12), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2100), .Z(new_n618));
  NAND2_X1  g193(.A1(new_n501), .A2(G123), .ZN(new_n619));
  OR2_X1    g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n620), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n621));
  INV_X1    g196(.A(G135), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n621), .C1(new_n622), .C2(new_n496), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n618), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT15), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2435), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2435), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT16), .B(G2443), .Z(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT80), .B(G2446), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT81), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n639), .A2(KEYINPUT81), .A3(G14), .A4(new_n640), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(G401));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT82), .Z(new_n647));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(KEYINPUT17), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n649), .B(new_n651), .C1(new_n647), .C2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n648), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n654), .A2(new_n646), .A3(new_n650), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT18), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n647), .A2(new_n652), .A3(new_n650), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT83), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT20), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n670), .A2(new_n662), .A3(new_n665), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n668), .B(new_n671), .C1(new_n662), .C2(new_n670), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  INV_X1    g250(.A(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n674), .B(new_n679), .ZN(G229));
  XNOR2_X1  g255(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n683), .A2(G6), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G305), .B2(G16), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT32), .B(G1981), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n685), .A2(new_n686), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n682), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(new_n681), .A3(new_n687), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n575), .A2(G16), .A3(new_n576), .A4(new_n578), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G16), .B2(G23), .ZN(new_n696));
  OR3_X1    g271(.A1(new_n695), .A2(G16), .A3(G23), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT89), .B(KEYINPUT33), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1976), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(G16), .A2(G22), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G166), .B2(G16), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT90), .B(G1971), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n694), .A2(new_n696), .A3(new_n697), .A4(new_n700), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n702), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n693), .A2(new_n708), .A3(KEYINPUT34), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT34), .B1(new_n693), .B2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G24), .ZN(new_n711));
  XOR2_X1   g286(.A(G290), .B(KEYINPUT85), .Z(new_n712));
  AOI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(new_n678), .ZN(new_n714));
  OR2_X1    g289(.A1(G95), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT84), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n501), .A2(G119), .ZN(new_n718));
  INV_X1    g293(.A(G131), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n496), .ZN(new_n720));
  MUX2_X1   g295(.A(G25), .B(new_n720), .S(G29), .Z(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT35), .B(G1991), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n721), .B(new_n722), .Z(new_n723));
  NAND4_X1  g298(.A1(new_n709), .A2(new_n710), .A3(new_n714), .A4(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT92), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT91), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n725), .B1(new_n724), .B2(new_n727), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n728), .A2(new_n729), .B1(KEYINPUT91), .B2(new_n726), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n724), .A2(new_n727), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(KEYINPUT92), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n726), .A2(KEYINPUT91), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G168), .A2(new_n683), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n683), .B2(G21), .ZN(new_n737));
  INV_X1    g312(.A(G1966), .ZN(new_n738));
  AOI22_X1  g313(.A1(G105), .A2(new_n486), .B1(new_n501), .B2(G129), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT95), .B(KEYINPUT26), .Z(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G141), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n739), .B(new_n742), .C1(new_n743), .C2(new_n496), .ZN(new_n744));
  MUX2_X1   g319(.A(G32), .B(new_n744), .S(G29), .Z(new_n745));
  XOR2_X1   g320(.A(KEYINPUT27), .B(G1996), .Z(new_n746));
  OAI22_X1  g321(.A1(new_n737), .A2(new_n738), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n683), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n683), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n745), .A2(new_n746), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  INV_X1    g328(.A(G29), .ZN(new_n754));
  NOR2_X1   g329(.A1(G164), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G27), .B2(new_n754), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n756), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n747), .B(new_n757), .C1(new_n753), .C2(new_n756), .ZN(new_n758));
  OR2_X1    g333(.A1(G29), .A2(G33), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  AOI22_X1  g336(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  INV_X1    g337(.A(G139), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n761), .B1(new_n461), .B2(new_n762), .C1(new_n496), .C2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(new_n754), .ZN(new_n765));
  INV_X1    g340(.A(G2072), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n683), .A2(KEYINPUT23), .A3(G20), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT23), .ZN(new_n769));
  INV_X1    g344(.A(G20), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(G16), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n768), .B(new_n771), .C1(new_n571), .C2(new_n683), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1956), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n765), .A2(new_n766), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT31), .B(G11), .Z(new_n775));
  NOR3_X1   g350(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n683), .A2(G19), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n559), .B2(new_n683), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1341), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n754), .A2(G26), .ZN(new_n780));
  OR2_X1    g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT94), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n501), .A2(G128), .ZN(new_n784));
  INV_X1    g359(.A(G140), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n496), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n780), .B1(new_n786), .B2(G29), .ZN(new_n787));
  MUX2_X1   g362(.A(new_n780), .B(new_n787), .S(KEYINPUT28), .Z(new_n788));
  INV_X1    g363(.A(G2067), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(KEYINPUT93), .B1(G4), .B2(G16), .ZN(new_n791));
  OR3_X1    g366(.A1(KEYINPUT93), .A2(G4), .A3(G16), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n791), .B(new_n792), .C1(new_n600), .C2(new_n683), .ZN(new_n793));
  INV_X1    g368(.A(G1348), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G28), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(KEYINPUT30), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT96), .Z(new_n798));
  AOI21_X1  g373(.A(G29), .B1(new_n796), .B2(KEYINPUT30), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n779), .A2(new_n790), .A3(new_n795), .A4(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n758), .A2(new_n767), .A3(new_n776), .A4(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G34), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n803), .A2(KEYINPUT24), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(KEYINPUT24), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n754), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G160), .B2(new_n754), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2084), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n754), .A2(G35), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G162), .B2(new_n754), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT29), .B(G2090), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n730), .A2(new_n735), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n737), .A2(new_n738), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n623), .A2(new_n754), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n814), .A2(new_n816), .A3(new_n817), .ZN(G311));
  AND3_X1   g393(.A1(new_n730), .A2(new_n735), .A3(new_n809), .ZN(new_n819));
  INV_X1    g394(.A(new_n817), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n819), .A2(new_n815), .A3(new_n820), .A4(new_n813), .ZN(G150));
  AOI22_X1  g396(.A1(new_n540), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n530), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n533), .A2(new_n824), .B1(new_n535), .B2(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G860), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(KEYINPUT98), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n823), .A2(new_n826), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n830), .A2(new_n558), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n559), .A2(new_n831), .A3(new_n832), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT39), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n600), .A2(new_n609), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n829), .B1(new_n841), .B2(G860), .ZN(G145));
  INV_X1    g417(.A(G142), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n461), .A2(G118), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n496), .A2(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G130), .B2(new_n501), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(new_n720), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT103), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n616), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n744), .B(new_n786), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT101), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n512), .A2(KEYINPUT99), .A3(new_n518), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT99), .B1(new_n512), .B2(new_n518), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n511), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n511), .B(KEYINPUT100), .C1(new_n854), .C2(new_n855), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n853), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n852), .A2(KEYINPUT101), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n852), .A2(KEYINPUT101), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n764), .B(KEYINPUT102), .Z(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n764), .A2(KEYINPUT102), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n860), .B2(new_n864), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n851), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n869), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(new_n850), .C1(new_n866), .C2(new_n865), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(G162), .B(G160), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(new_n623), .Z(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n870), .A2(new_n872), .A3(new_n875), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g456(.A1(new_n827), .A2(new_n601), .ZN(new_n882));
  XOR2_X1   g457(.A(G288), .B(G290), .Z(new_n883));
  OR2_X1    g458(.A1(new_n883), .A2(KEYINPUT108), .ZN(new_n884));
  XNOR2_X1  g459(.A(G303), .B(KEYINPUT107), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(G305), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(KEYINPUT108), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OR3_X1    g463(.A1(new_n886), .A2(new_n883), .A3(KEYINPUT108), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT42), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n571), .A2(KEYINPUT104), .A3(new_n600), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT104), .B1(new_n571), .B2(new_n600), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(G299), .A2(new_n608), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT105), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n836), .B(new_n611), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  INV_X1    g476(.A(new_n894), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(KEYINPUT106), .A3(new_n892), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n896), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n895), .A2(KEYINPUT106), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n897), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT41), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n900), .B1(new_n899), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n891), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n882), .B1(new_n911), .B2(new_n601), .ZN(G295));
  OAI21_X1  g487(.A(new_n882), .B1(new_n911), .B2(new_n601), .ZN(G331));
  XNOR2_X1  g488(.A(G171), .B(KEYINPUT110), .ZN(new_n914));
  AOI21_X1  g489(.A(G286), .B1(new_n834), .B2(new_n835), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n834), .A2(G286), .A3(new_n835), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  INV_X1    g494(.A(new_n914), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n919), .A2(new_n920), .A3(new_n915), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n907), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n920), .B1(new_n919), .B2(new_n915), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n916), .A2(new_n914), .A3(new_n917), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n906), .A2(new_n923), .A3(new_n924), .A4(new_n908), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n890), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OR3_X1    g503(.A1(new_n904), .A2(new_n905), .A3(new_n901), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n897), .A2(new_n901), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n929), .A2(new_n924), .A3(new_n923), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n898), .B1(new_n921), .B2(new_n918), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n890), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n890), .B1(new_n926), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT111), .B1(new_n922), .B2(new_n925), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n928), .B(new_n936), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n935), .A2(new_n940), .A3(KEYINPUT44), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n934), .A2(new_n936), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n928), .B(KEYINPUT43), .C1(new_n938), .C2(new_n939), .ZN(new_n943));
  XOR2_X1   g518(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n945), .ZN(G397));
  AOI21_X1  g521(.A(G1384), .B1(new_n858), .B2(new_n859), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(KEYINPUT45), .ZN(new_n948));
  INV_X1    g523(.A(G40), .ZN(new_n949));
  AOI211_X1 g524(.A(new_n949), .B(new_n465), .C1(new_n493), .C2(new_n494), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n720), .B(new_n722), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT112), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n744), .B(G1996), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n786), .B(G2067), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(G290), .B(G1986), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n952), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1956), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n493), .A2(new_n494), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n521), .A2(KEYINPUT117), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n504), .A2(KEYINPUT4), .B1(new_n509), .B2(new_n462), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n963), .B(new_n964), .C1(new_n966), .C2(new_n519), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT117), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n465), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n962), .A2(new_n970), .A3(G40), .A4(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT99), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n519), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n512), .A2(KEYINPUT99), .A3(new_n518), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n966), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n976), .A2(KEYINPUT113), .A3(G1384), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n856), .B2(new_n964), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n977), .A2(new_n979), .A3(new_n963), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n961), .B1(new_n972), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n571), .A2(KEYINPUT120), .A3(new_n982), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n982), .A2(KEYINPUT120), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(KEYINPUT120), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n984), .B(new_n985), .C1(new_n567), .C2(new_n570), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n862), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n521), .A2(new_n964), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT56), .B(G2072), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n950), .A2(new_n988), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n981), .A2(new_n987), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n981), .A2(new_n993), .ZN(new_n996));
  INV_X1    g571(.A(new_n987), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT121), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT121), .ZN(new_n999));
  AOI211_X1 g574(.A(new_n999), .B(new_n987), .C1(new_n981), .C2(new_n993), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n989), .A2(KEYINPUT50), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n962), .A2(G40), .A3(new_n971), .A4(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT113), .B1(new_n976), .B2(G1384), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n856), .A2(new_n978), .A3(new_n964), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT50), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n794), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n950), .A2(new_n789), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n608), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n995), .B1(new_n1001), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n996), .A2(new_n997), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT122), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(new_n994), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT123), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n987), .B1(new_n981), .B2(new_n993), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT61), .B1(new_n1017), .B2(KEYINPUT122), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1016), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1010), .A2(KEYINPUT60), .A3(new_n600), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1007), .A2(new_n600), .A3(new_n1009), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1011), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1024), .B2(KEYINPUT60), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT61), .B(new_n994), .C1(new_n998), .C2(new_n1000), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n950), .A2(new_n988), .A3(new_n991), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(G1996), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT58), .B(G1341), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n950), .B2(new_n1008), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n559), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT59), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1033), .B(new_n559), .C1(new_n1028), .C2(new_n1030), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1025), .A2(new_n1026), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1012), .B1(new_n1021), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G303), .A2(G8), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT55), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n972), .A2(new_n980), .A3(G2090), .ZN(new_n1040));
  INV_X1    g615(.A(G1971), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n1027), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1039), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n962), .A2(G40), .A3(new_n971), .A4(new_n991), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n990), .B(G1384), .C1(new_n858), .C2(new_n859), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1041), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1008), .A2(new_n963), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(new_n950), .A3(new_n1002), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1049), .B2(G2090), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1039), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(G8), .A3(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n575), .A2(G1976), .A3(new_n576), .A4(new_n578), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n962), .A2(G40), .A3(new_n971), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n977), .A2(new_n979), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1053), .B(G8), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT52), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n950), .A2(new_n1008), .ZN(new_n1058));
  INV_X1    g633(.A(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1058), .A2(new_n1060), .A3(G8), .A4(new_n1053), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n587), .A2(new_n676), .A3(new_n588), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n546), .A2(G48), .ZN(new_n1063));
  INV_X1    g638(.A(new_n586), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1064), .B2(new_n584), .ZN(new_n1065));
  NOR2_X1   g640(.A1(KEYINPUT114), .A2(G86), .ZN(new_n1066));
  AND2_X1   g641(.A1(KEYINPUT114), .A2(G86), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n533), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G1981), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1062), .A2(new_n1069), .A3(KEYINPUT49), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT49), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1058), .A2(new_n1072), .A3(G8), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1057), .A2(new_n1061), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1044), .A2(new_n1052), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT126), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n950), .A2(new_n988), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(G2078), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n947), .B2(KEYINPUT45), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1077), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1080), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n862), .A2(new_n964), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1083), .B1(new_n1084), .B2(new_n990), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1085), .A2(KEYINPUT126), .A3(new_n988), .A4(new_n950), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n750), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1045), .A2(new_n1046), .A3(G2078), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(KEYINPUT53), .ZN(new_n1090));
  OAI21_X1  g665(.A(G171), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1004), .A2(new_n990), .A3(new_n1005), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n521), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n950), .A2(new_n1092), .A3(new_n1093), .A4(new_n1080), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1088), .B(new_n1094), .C1(new_n1089), .C2(KEYINPUT53), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1091), .B(KEYINPUT54), .C1(G171), .C2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G168), .A2(new_n1043), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT51), .B1(new_n1097), .B2(KEYINPUT124), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1099));
  INV_X1    g674(.A(G2084), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n950), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n738), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(G8), .B(new_n1098), .C1(new_n1104), .C2(G286), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1097), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1098), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1099), .A2(new_n1100), .B1(new_n1102), .B2(new_n738), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1106), .B(new_n1107), .C1(new_n1108), .C2(new_n1043), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(G8), .A3(G286), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1105), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1087), .A2(G171), .A3(new_n1090), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1095), .A2(new_n1113), .A3(G171), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1113), .B1(new_n1095), .B2(G171), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1096), .B(new_n1111), .C1(new_n1116), .C2(KEYINPUT54), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1037), .A2(new_n1076), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1052), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1104), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n1122));
  INV_X1    g697(.A(G2090), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1099), .A2(new_n1123), .B1(new_n1027), .B2(new_n1041), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1039), .B1(new_n1124), .B2(new_n1043), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1122), .B1(new_n1125), .B2(new_n1075), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1051), .B1(new_n1050), .B2(G8), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1127), .A2(KEYINPUT118), .A3(new_n1074), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1121), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1104), .A2(G8), .A3(G168), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1076), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT119), .B(new_n1121), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1131), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(G288), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1073), .A2(new_n1059), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1062), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT116), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT116), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1138), .A2(new_n1141), .A3(new_n1062), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1058), .A2(G8), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT115), .Z(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1052), .B2(new_n1074), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1105), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1076), .B1(new_n1111), .B2(KEYINPUT62), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1146), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1136), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n960), .B1(new_n1118), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n786), .A2(G2067), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n720), .A2(new_n722), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n957), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(new_n951), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n951), .A2(G1996), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1159), .A2(KEYINPUT46), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n952), .B1(new_n744), .B2(new_n956), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(KEYINPUT46), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT47), .Z(new_n1164));
  NAND2_X1  g739(.A1(new_n958), .A2(new_n952), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n951), .A2(G1986), .A3(G290), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT127), .Z(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT48), .ZN(new_n1168));
  AOI211_X1 g743(.A(new_n1158), .B(new_n1164), .C1(new_n1165), .C2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1154), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g745(.A(new_n459), .B1(new_n643), .B2(new_n644), .ZN(new_n1172));
  NAND4_X1  g746(.A1(new_n880), .A2(new_n942), .A3(new_n943), .A4(new_n1172), .ZN(new_n1173));
  NOR2_X1   g747(.A1(G229), .A2(G227), .ZN(new_n1174));
  INV_X1    g748(.A(new_n1174), .ZN(new_n1175));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1175), .ZN(G308));
  AND2_X1   g750(.A1(new_n942), .A2(new_n943), .ZN(new_n1177));
  NAND4_X1  g751(.A1(new_n1177), .A2(new_n880), .A3(new_n1174), .A4(new_n1172), .ZN(G225));
endmodule


