//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043;
  XOR2_X1   g000(.A(G125), .B(G140), .Z(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G146), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT73), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n192), .B1(new_n189), .B2(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT24), .B(G110), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT79), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n190), .A2(KEYINPUT74), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(KEYINPUT23), .ZN(new_n200));
  OR2_X1    g014(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n199), .A2(new_n200), .B1(new_n190), .B2(new_n201), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT78), .B(G110), .Z(new_n203));
  AOI22_X1  g017(.A1(new_n197), .A2(new_n198), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n195), .A2(KEYINPUT79), .A3(new_n196), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n188), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT75), .B(G125), .ZN(new_n207));
  NOR3_X1   g021(.A1(new_n207), .A2(KEYINPUT16), .A3(G140), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT75), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT75), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G125), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n210), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(G125), .A2(G140), .ZN(new_n216));
  OAI211_X1 g030(.A(KEYINPUT76), .B(KEYINPUT16), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n216), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n207), .B2(new_n210), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT76), .B1(new_n220), .B2(KEYINPUT16), .ZN(new_n221));
  OAI211_X1 g035(.A(G146), .B(new_n209), .C1(new_n218), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n206), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n209), .B1(new_n218), .B2(new_n221), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n222), .ZN(new_n227));
  INV_X1    g041(.A(G110), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n202), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n195), .A2(new_n196), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT77), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT77), .ZN(new_n234));
  AOI211_X1 g048(.A(new_n234), .B(new_n231), .C1(new_n226), .C2(new_n222), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n223), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT22), .B(G137), .ZN(new_n237));
  INV_X1    g051(.A(G953), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n238), .A2(G221), .A3(G234), .ZN(new_n239));
  XOR2_X1   g053(.A(new_n237), .B(new_n239), .Z(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT76), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n212), .A2(new_n214), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n216), .B1(new_n244), .B2(G140), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT16), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n243), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n217), .ZN(new_n248));
  AOI21_X1  g062(.A(G146), .B1(new_n248), .B2(new_n209), .ZN(new_n249));
  AOI211_X1 g063(.A(new_n225), .B(new_n208), .C1(new_n247), .C2(new_n217), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n232), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n234), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n227), .A2(KEYINPUT77), .A3(new_n232), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n223), .A3(new_n240), .ZN(new_n255));
  INV_X1    g069(.A(G902), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n242), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n242), .A2(new_n255), .A3(KEYINPUT25), .A4(new_n256), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G217), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n262), .B1(G234), .B2(new_n256), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT80), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT80), .ZN(new_n265));
  INV_X1    g079(.A(new_n263), .ZN(new_n266));
  AOI211_X1 g080(.A(new_n265), .B(new_n266), .C1(new_n259), .C2(new_n260), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n240), .B1(new_n254), .B2(new_n223), .ZN(new_n268));
  INV_X1    g082(.A(new_n223), .ZN(new_n269));
  AOI211_X1 g083(.A(new_n269), .B(new_n241), .C1(new_n252), .C2(new_n253), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n263), .A2(G902), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n264), .A2(new_n267), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G472), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT11), .ZN(new_n278));
  INV_X1    g092(.A(G134), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(new_n279), .B2(G137), .ZN(new_n280));
  INV_X1    g094(.A(G137), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT11), .A3(G134), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(G137), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT64), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT64), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n280), .A2(new_n282), .A3(new_n286), .A4(new_n283), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(G131), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G131), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n280), .A2(new_n282), .A3(new_n289), .A4(new_n283), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT65), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n225), .A2(G143), .ZN(new_n294));
  INV_X1    g108(.A(G143), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G146), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(KEYINPUT0), .A2(G128), .ZN(new_n298));
  OR2_X1    g112(.A1(KEYINPUT0), .A2(G128), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(G143), .B(G146), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT0), .A3(G128), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n285), .A2(KEYINPUT65), .A3(G131), .A4(new_n287), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n293), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n279), .A2(G137), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n281), .A2(G134), .ZN(new_n307));
  OAI21_X1  g121(.A(G131), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G128), .ZN(new_n309));
  AND2_X1   g123(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n310));
  NOR2_X1   g124(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n294), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n309), .B1(new_n312), .B2(KEYINPUT68), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(new_n294), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n301), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n297), .A2(new_n314), .A3(new_n309), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n290), .B(new_n308), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT69), .ZN(new_n320));
  INV_X1    g134(.A(G116), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(G119), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n189), .A2(KEYINPUT69), .A3(G116), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(G119), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT2), .B(G113), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n326), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT70), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n328), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AND4_X1   g147(.A1(new_n305), .A2(new_n319), .A3(new_n330), .A4(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n277), .B1(new_n334), .B2(KEYINPUT28), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n305), .A2(new_n319), .B1(new_n330), .B2(new_n333), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT28), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n305), .A2(new_n319), .A3(new_n330), .A4(new_n333), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT28), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(KEYINPUT71), .A3(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(G237), .A2(G953), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G210), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT27), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT26), .B(G101), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n335), .A2(new_n337), .A3(new_n340), .A4(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n349), .A2(new_n256), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n290), .A2(new_n308), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT66), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT66), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n290), .A2(new_n308), .A3(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n352), .B(new_n354), .C1(new_n317), .C2(new_n318), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n329), .B1(new_n305), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT28), .B1(new_n334), .B2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n357), .A2(new_n335), .A3(new_n340), .A4(new_n345), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(new_n305), .B2(new_n319), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n305), .A2(new_n355), .A3(new_n359), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n329), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n346), .B1(new_n363), .B2(new_n334), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n358), .A2(new_n364), .A3(new_n347), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n276), .B1(new_n350), .B2(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n305), .A2(new_n355), .A3(new_n359), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n331), .B1(new_n367), .B2(new_n360), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n338), .A3(new_n345), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT31), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n368), .A2(KEYINPUT31), .A3(new_n338), .A4(new_n345), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n357), .A2(new_n335), .A3(new_n340), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n371), .A2(new_n372), .B1(new_n373), .B2(new_n346), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n374), .A2(G472), .A3(G902), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n366), .B1(new_n375), .B2(KEYINPUT32), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n372), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n346), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n276), .A3(new_n256), .ZN(new_n380));
  XOR2_X1   g194(.A(KEYINPUT72), .B(KEYINPUT32), .Z(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G221), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT9), .B(G234), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n387), .B2(new_n256), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n312), .A2(KEYINPUT68), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n316), .A3(G128), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n318), .B1(new_n390), .B2(new_n297), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT81), .B(G101), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G107), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n393), .B2(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G104), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n392), .A2(new_n394), .A3(new_n395), .A4(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n394), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n393), .A2(G107), .ZN(new_n401));
  OAI21_X1  g215(.A(G101), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(KEYINPUT10), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT82), .B1(new_n391), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n403), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT82), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n405), .B(new_n406), .C1(new_n317), .C2(new_n318), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n395), .A2(new_n398), .A3(new_n394), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G101), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n411), .B2(new_n399), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT4), .B1(new_n410), .B2(G101), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n303), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n225), .A2(G143), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT1), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n301), .B2(G128), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n318), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n399), .A2(new_n402), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n415), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n408), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n293), .A2(new_n304), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n408), .A2(KEYINPUT83), .A3(new_n422), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G110), .B(G140), .ZN(new_n430));
  INV_X1    g244(.A(G227), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(G953), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n430), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n414), .A2(new_n421), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n404), .B2(new_n407), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n433), .B1(new_n435), .B2(new_n426), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT12), .ZN(new_n438));
  OR3_X1    g252(.A1(new_n297), .A2(new_n314), .A3(new_n309), .ZN(new_n439));
  INV_X1    g253(.A(new_n418), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n420), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(new_n391), .B2(new_n420), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n438), .B1(new_n442), .B2(new_n426), .ZN(new_n443));
  INV_X1    g257(.A(new_n420), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n318), .B2(new_n418), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n390), .A2(new_n297), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n439), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n447), .B2(new_n444), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT12), .A3(new_n427), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n408), .A2(new_n426), .A3(new_n422), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n433), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n437), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G469), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n454), .A2(KEYINPUT84), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n457));
  INV_X1    g271(.A(new_n433), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n426), .B1(new_n423), .B2(new_n424), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n460), .B2(new_n428), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n458), .B1(new_n450), .B2(new_n451), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n256), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n457), .B1(new_n463), .B2(G469), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n456), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n458), .B1(new_n429), .B2(new_n451), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n442), .A2(new_n438), .A3(new_n426), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT12), .B1(new_n448), .B2(new_n427), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n443), .A2(new_n449), .A3(KEYINPUT85), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n470), .A2(new_n436), .A3(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n455), .B(new_n256), .C1(new_n466), .C2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT86), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n470), .A2(new_n436), .A3(new_n471), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n460), .A2(new_n428), .B1(new_n426), .B2(new_n435), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n458), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n478), .A2(KEYINPUT86), .A3(new_n455), .A4(new_n256), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n388), .B1(new_n465), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT15), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G478), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT96), .ZN(new_n484));
  INV_X1    g298(.A(G122), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT92), .B1(new_n485), .B2(G116), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n321), .A3(G122), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(G116), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n397), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n309), .A2(G143), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n295), .A2(G128), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n492), .A2(new_n493), .A3(new_n279), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n279), .B1(new_n492), .B2(new_n493), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n295), .A2(G128), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n309), .A2(G143), .ZN(new_n499));
  OAI21_X1  g313(.A(G134), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n492), .A2(new_n493), .A3(new_n279), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT95), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n491), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n489), .A2(KEYINPUT14), .B1(G116), .B2(new_n485), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n486), .A2(new_n488), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n397), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n484), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n489), .A2(new_n397), .A3(new_n490), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n496), .B1(new_n494), .B2(new_n495), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n500), .A2(KEYINPUT95), .A3(new_n501), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n489), .A2(KEYINPUT14), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n506), .A3(new_n490), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G107), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(KEYINPUT96), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT13), .ZN(new_n518));
  OAI211_X1 g332(.A(KEYINPUT93), .B(new_n493), .C1(new_n498), .C2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n493), .B2(new_n518), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n499), .A2(KEYINPUT94), .A3(KEYINPUT13), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n499), .B1(KEYINPUT13), .B2(new_n492), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(KEYINPUT93), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n279), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n397), .B1(new_n489), .B2(new_n490), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n501), .B1(new_n509), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n386), .A2(new_n262), .A3(G953), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n517), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(new_n517), .B2(new_n529), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n256), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT97), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n503), .A2(new_n484), .A3(new_n507), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT96), .B1(new_n512), .B2(new_n515), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n529), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n530), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n517), .A2(new_n529), .A3(new_n530), .ZN(new_n541));
  AOI21_X1  g355(.A(G902), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT97), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n483), .B1(new_n535), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n483), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n533), .B2(new_n534), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT98), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n542), .A2(KEYINPUT97), .ZN(new_n548));
  AOI211_X1 g362(.A(new_n534), .B(G902), .C1(new_n540), .C2(new_n541), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n546), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT98), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n188), .B1(G146), .B2(new_n245), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G237), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(new_n238), .A3(G214), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n295), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n341), .A2(G143), .A3(G214), .ZN(new_n560));
  NAND2_X1  g374(.A1(KEYINPUT18), .A2(G131), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n560), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(KEYINPUT18), .A3(G131), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n556), .A2(KEYINPUT89), .A3(new_n562), .A4(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT89), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n562), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n566), .B1(new_n567), .B2(new_n555), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n559), .A2(new_n289), .A3(new_n560), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT90), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n559), .A2(KEYINPUT90), .A3(new_n289), .A4(new_n560), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n563), .A2(G131), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n245), .A2(KEYINPUT19), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(KEYINPUT19), .B2(new_n187), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n222), .B(new_n575), .C1(G146), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n569), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(G113), .B(G122), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(new_n393), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT17), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n572), .A2(new_n574), .A3(new_n584), .A4(new_n573), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n563), .A2(KEYINPUT17), .A3(G131), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n226), .A2(new_n222), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n581), .A3(new_n569), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT91), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n587), .A2(new_n581), .A3(new_n569), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n581), .B1(new_n569), .B2(new_n578), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(G475), .A2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OAI22_X1  g408(.A1(KEYINPUT20), .A2(new_n589), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n583), .A2(new_n588), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT20), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n596), .A2(KEYINPUT91), .A3(new_n597), .A4(new_n593), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n581), .B1(new_n587), .B2(new_n569), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n256), .B1(new_n590), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G475), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(G110), .B(G122), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT8), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT5), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n189), .A3(G116), .ZN(new_n607));
  OAI211_X1 g421(.A(G113), .B(new_n607), .C1(new_n325), .C2(new_n606), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n444), .A2(new_n327), .A3(new_n608), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n608), .A2(new_n327), .B1(new_n402), .B2(new_n399), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n444), .A2(new_n327), .A3(new_n608), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n412), .A2(new_n413), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n604), .B(new_n612), .C1(new_n613), .C2(new_n329), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n303), .A2(new_n244), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n391), .B2(new_n244), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT87), .B(G224), .Z(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(G953), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n617), .A2(KEYINPUT7), .A3(new_n620), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n619), .B(new_n616), .C1(new_n391), .C2(new_n244), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT7), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n623), .B(new_n616), .C1(new_n391), .C2(new_n244), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT88), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n625), .B1(new_n622), .B2(new_n624), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n615), .B(new_n621), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n612), .B1(new_n613), .B2(new_n329), .ZN(new_n630));
  INV_X1    g444(.A(new_n604), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(KEYINPUT6), .A3(new_n614), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n617), .A2(new_n620), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n622), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT6), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n630), .A2(new_n636), .A3(new_n631), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n633), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n629), .A2(new_n638), .A3(new_n256), .ZN(new_n639));
  OAI21_X1  g453(.A(G210), .B1(G237), .B2(G902), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n303), .A2(new_n244), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n447), .B2(new_n207), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n644), .B(KEYINPUT88), .C1(new_n623), .C2(new_n619), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n626), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n621), .A2(new_n614), .A3(new_n611), .ZN(new_n647));
  AOI21_X1  g461(.A(G902), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n640), .A3(new_n638), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(G214), .B1(G237), .B2(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(G234), .A2(G237), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(G952), .A3(new_n238), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(G902), .A3(G953), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT21), .B(G898), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n650), .A2(new_n651), .A3(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n554), .A2(new_n603), .A3(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n275), .A2(new_n384), .A3(new_n481), .A4(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(new_n392), .Z(G3));
  AOI21_X1  g477(.A(KEYINPUT25), .B1(new_n271), .B2(new_n256), .ZN(new_n664));
  INV_X1    g478(.A(new_n260), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n263), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n265), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n261), .A2(KEYINPUT80), .A3(new_n263), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n276), .B1(new_n379), .B2(new_n256), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n375), .ZN(new_n670));
  AND4_X1   g484(.A1(new_n667), .A2(new_n668), .A3(new_n273), .A4(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(new_n481), .ZN(new_n672));
  INV_X1    g486(.A(new_n651), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n640), .B1(new_n648), .B2(new_n638), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(KEYINPUT99), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT99), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n642), .A2(new_n676), .A3(new_n649), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n659), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n540), .A2(new_n541), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n682));
  OR2_X1    g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(KEYINPUT100), .A2(KEYINPUT33), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n256), .A2(G478), .ZN(new_n687));
  OAI22_X1  g501(.A1(new_n686), .A2(new_n687), .B1(G478), .B2(new_n542), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n603), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n672), .A2(new_n680), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT34), .B(G104), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G6));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n694), .B(new_n597), .C1(new_n592), .C2(new_n594), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n597), .ZN(new_n696));
  NAND2_X1  g510(.A1(KEYINPUT101), .A2(KEYINPUT20), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n596), .A2(new_n593), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n695), .A2(new_n602), .A3(new_n698), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n554), .A2(new_n678), .A3(new_n659), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n672), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT35), .B(G107), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G9));
  NOR2_X1   g517(.A1(new_n241), .A2(KEYINPUT36), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n236), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n272), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n667), .A2(new_n668), .A3(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(new_n481), .A3(new_n661), .A4(new_n670), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT37), .B(G110), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G12));
  NAND2_X1  g524(.A1(new_n675), .A2(new_n677), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n376), .B2(new_n383), .ZN(new_n712));
  INV_X1    g526(.A(G900), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n656), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n653), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n554), .A2(new_n699), .A3(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n707), .A2(new_n712), .A3(new_n481), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  XNOR2_X1  g532(.A(new_n715), .B(KEYINPUT39), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n481), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT40), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n379), .A2(KEYINPUT32), .A3(new_n276), .A4(new_n256), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n346), .B1(new_n334), .B2(new_n336), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n369), .A2(G472), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n276), .A2(new_n256), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT102), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n383), .A2(new_n722), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n650), .B(KEYINPUT38), .Z(new_n731));
  NOR2_X1   g545(.A1(new_n264), .A2(new_n267), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n595), .A2(new_n598), .B1(G475), .B2(new_n601), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n547), .B2(new_n553), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n732), .A2(new_n651), .A3(new_n706), .A4(new_n734), .ZN(new_n735));
  AOI211_X1 g549(.A(new_n730), .B(new_n731), .C1(new_n735), .C2(KEYINPUT103), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n721), .B(new_n736), .C1(KEYINPUT103), .C2(new_n735), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G143), .ZN(G45));
  NAND3_X1  g552(.A1(new_n603), .A2(new_n688), .A3(new_n715), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n707), .A2(new_n712), .A3(new_n481), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G146), .ZN(G48));
  NAND4_X1  g556(.A1(new_n275), .A2(new_n384), .A3(new_n680), .A4(new_n690), .ZN(new_n743));
  INV_X1    g557(.A(new_n388), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n478), .A2(new_n256), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(G469), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n480), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n480), .A2(KEYINPUT104), .A3(new_n744), .A4(new_n746), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT41), .B(G113), .Z(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G15));
  NAND3_X1  g568(.A1(new_n275), .A2(new_n384), .A3(new_n700), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n751), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n321), .ZN(G18));
  AND3_X1   g571(.A1(new_n480), .A2(new_n744), .A3(new_n746), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n554), .A2(new_n603), .A3(new_n658), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n707), .A2(new_n712), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G119), .ZN(G21));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  AND4_X1   g576(.A1(new_n762), .A2(new_n554), .A3(new_n678), .A4(new_n603), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n762), .B1(new_n734), .B2(new_n678), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n659), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n335), .A2(new_n337), .A3(new_n340), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n346), .ZN(new_n767));
  AOI211_X1 g581(.A(G472), .B(G902), .C1(new_n377), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n669), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n275), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n765), .A2(new_n751), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n485), .ZN(G24));
  AND4_X1   g586(.A1(new_n744), .A2(new_n480), .A3(new_n678), .A4(new_n746), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(new_n707), .A3(new_n740), .A4(new_n769), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G125), .ZN(G27));
  NAND2_X1  g589(.A1(new_n732), .A2(new_n273), .ZN(new_n776));
  INV_X1    g590(.A(new_n366), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n383), .A2(new_n722), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n475), .A2(new_n479), .B1(G469), .B2(new_n463), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n388), .A2(new_n673), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n642), .A2(new_n649), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n739), .A2(KEYINPUT42), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n779), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n376), .B1(KEYINPUT32), .B2(new_n375), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n275), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n780), .A2(new_n739), .A3(new_n782), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT42), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G131), .ZN(G33));
  NAND4_X1  g606(.A1(new_n275), .A2(new_n384), .A3(new_n716), .A4(new_n783), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G134), .ZN(G36));
  NAND2_X1  g608(.A1(new_n733), .A2(new_n688), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT43), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n670), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(KEYINPUT44), .A3(new_n707), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT108), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n461), .B2(new_n462), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n437), .A2(new_n453), .A3(KEYINPUT45), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n802), .A3(G469), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n455), .B2(new_n256), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT46), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT107), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n480), .B1(new_n804), .B2(new_n805), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT106), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n808), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n744), .A3(new_n719), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT44), .B1(new_n797), .B2(new_n707), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n642), .A2(new_n649), .A3(new_n651), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n799), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(KEYINPUT109), .B(G137), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(G39));
  NOR4_X1   g636(.A1(new_n275), .A2(new_n384), .A3(new_n739), .A4(new_n818), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n813), .A2(KEYINPUT47), .A3(new_n744), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT47), .B1(new_n813), .B2(new_n744), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  NAND2_X1  g642(.A1(new_n758), .A2(new_n673), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT116), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n770), .A2(new_n653), .A3(new_n796), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n731), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT50), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n796), .A2(new_n653), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n747), .A2(new_n818), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n707), .A2(new_n834), .A3(new_n769), .A4(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n275), .A3(new_n654), .A4(new_n730), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n837), .A2(new_n603), .A3(new_n688), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n833), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n825), .A2(new_n826), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n480), .A2(new_n746), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n840), .B1(new_n744), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n817), .A3(new_n831), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT51), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n275), .A2(new_n834), .A3(new_n786), .A4(new_n835), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT48), .ZN(new_n846));
  INV_X1    g660(.A(G952), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n847), .B(G953), .C1(new_n831), .C2(new_n773), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n689), .B2(new_n837), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n844), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n839), .A2(KEYINPUT51), .A3(new_n843), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n774), .A2(new_n717), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n729), .B1(new_n763), .B2(new_n764), .ZN(new_n855));
  INV_X1    g669(.A(new_n780), .ZN(new_n856));
  INV_X1    g670(.A(new_n715), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n388), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n732), .A2(new_n856), .A3(new_n706), .A4(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(KEYINPUT52), .B(new_n741), .C1(new_n855), .C2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n853), .B1(new_n774), .B2(new_n717), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n854), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  XOR2_X1   g676(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n734), .A2(new_n678), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT105), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n734), .A2(new_n762), .A3(new_n678), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n730), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n858), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n707), .A2(new_n780), .A3(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n707), .A2(new_n481), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n778), .A2(new_n711), .A3(new_n739), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n868), .A2(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n774), .A2(new_n717), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n864), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT114), .B1(new_n862), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(KEYINPUT112), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n774), .A2(new_n717), .A3(new_n853), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n873), .A3(KEYINPUT52), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT114), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n741), .B1(new_n855), .B2(new_n859), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n863), .B1(new_n882), .B2(new_n874), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n877), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n660), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n671), .A2(new_n481), .A3(new_n886), .A4(new_n690), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT110), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n887), .A2(new_n888), .A3(new_n662), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n888), .B1(new_n887), .B2(new_n662), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n751), .B1(new_n743), .B2(new_n755), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n733), .B1(new_n544), .B2(new_n546), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n660), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n275), .A2(new_n894), .A3(new_n481), .A4(new_n670), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n760), .A3(new_n708), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n771), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n788), .A2(new_n707), .A3(new_n769), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n544), .A2(new_n546), .A3(new_n857), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n899), .A2(new_n699), .A3(new_n817), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n707), .A2(new_n384), .A3(new_n481), .A4(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n793), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT111), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n793), .A2(new_n898), .A3(new_n901), .A4(KEYINPUT111), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND4_X1   g720(.A1(new_n791), .A2(new_n891), .A3(new_n897), .A4(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT53), .B1(new_n885), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n904), .B2(new_n905), .ZN(new_n910));
  AND4_X1   g724(.A1(new_n791), .A2(new_n910), .A3(new_n891), .A4(new_n897), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n882), .A2(new_n874), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT52), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT54), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT53), .B1(new_n907), .B2(new_n913), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n885), .A2(KEYINPUT115), .A3(new_n911), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT115), .B1(new_n885), .B2(new_n911), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n915), .B1(new_n920), .B2(KEYINPUT54), .ZN(new_n921));
  OAI22_X1  g735(.A1(new_n852), .A2(new_n921), .B1(G952), .B2(G953), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n841), .B(KEYINPUT49), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n731), .A2(new_n733), .A3(new_n688), .A4(new_n781), .ZN(new_n924));
  OR3_X1    g738(.A1(new_n924), .A2(new_n776), .A3(new_n729), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n922), .B1(new_n923), .B2(new_n925), .ZN(G75));
  NAND2_X1  g740(.A1(new_n847), .A2(G953), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT119), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n920), .A2(G210), .A3(G902), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n633), .A2(new_n637), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n635), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT55), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n929), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT117), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n920), .A2(KEYINPUT117), .A3(G210), .A4(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n936), .A2(new_n942), .ZN(G51));
  XNOR2_X1  g757(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n455), .A2(new_n256), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT54), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT115), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n881), .B1(new_n880), .B2(new_n883), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n910), .A2(new_n891), .A3(new_n897), .A4(new_n791), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n885), .A2(new_n911), .A3(KEYINPUT115), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n947), .B1(new_n955), .B2(new_n917), .ZN(new_n956));
  AOI211_X1 g770(.A(KEYINPUT54), .B(new_n916), .C1(new_n953), .C2(new_n954), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n946), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n478), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n920), .A2(G902), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n960), .A2(new_n803), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n929), .B1(new_n959), .B2(new_n961), .ZN(G54));
  NAND2_X1  g776(.A1(KEYINPUT58), .A2(G475), .ZN(new_n963));
  OR3_X1    g777(.A1(new_n960), .A2(new_n596), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n596), .B1(new_n960), .B2(new_n963), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n929), .B1(new_n964), .B2(new_n965), .ZN(G60));
  NOR2_X1   g780(.A1(new_n956), .A2(new_n957), .ZN(new_n967));
  INV_X1    g781(.A(new_n686), .ZN(new_n968));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT59), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n928), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n968), .B1(new_n921), .B2(new_n970), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(G63));
  INV_X1    g788(.A(KEYINPUT121), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT61), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n928), .B1(new_n975), .B2(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT60), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n920), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n271), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n920), .A2(new_n705), .A3(new_n980), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n976), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n916), .B1(new_n953), .B2(new_n954), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n982), .B1(new_n986), .B2(new_n979), .ZN(new_n987));
  INV_X1    g801(.A(new_n977), .ZN(new_n988));
  AND4_X1   g802(.A1(new_n976), .A2(new_n987), .A3(new_n984), .A4(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n985), .A2(new_n989), .ZN(G66));
  NOR2_X1   g804(.A1(new_n618), .A2(new_n657), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n991), .A2(new_n238), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n891), .A2(new_n897), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(new_n238), .ZN(new_n994));
  INV_X1    g808(.A(G898), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n933), .B1(new_n995), .B2(G953), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n994), .B(new_n996), .ZN(G69));
  NAND2_X1  g811(.A1(new_n361), .A2(new_n362), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(new_n577), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n854), .A2(new_n861), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n1000), .A2(new_n741), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n785), .A2(new_n790), .A3(new_n793), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n787), .B1(new_n867), .B2(new_n866), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n815), .B2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n820), .A2(new_n1001), .A3(new_n827), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n238), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n713), .A2(G953), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n999), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n737), .A2(new_n1000), .A3(new_n741), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n818), .B1(new_n689), .B2(new_n893), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n779), .A2(new_n720), .A3(new_n1011), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n820), .A2(new_n827), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT122), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n1009), .A2(new_n1014), .A3(KEYINPUT62), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1014), .B1(new_n1009), .B2(KEYINPUT62), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1010), .B(new_n1013), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n238), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1008), .B1(new_n1018), .B2(new_n999), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n238), .B1(G227), .B2(G900), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT123), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1019), .B(new_n1021), .ZN(G72));
  INV_X1    g836(.A(KEYINPUT126), .ZN(new_n1023));
  XNOR2_X1  g837(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(new_n725), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1025), .B1(new_n1005), .B2(new_n993), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n368), .A2(new_n338), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1027), .B(KEYINPUT125), .Z(new_n1028));
  NOR2_X1   g842(.A1(new_n1028), .A2(new_n345), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1023), .B1(new_n1030), .B2(new_n928), .ZN(new_n1031));
  AOI211_X1 g845(.A(KEYINPUT126), .B(new_n929), .C1(new_n1026), .C2(new_n1029), .ZN(new_n1032));
  OR2_X1    g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT127), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1025), .B1(new_n1017), .B2(new_n993), .ZN(new_n1035));
  AND2_X1   g849(.A1(new_n1028), .A2(new_n345), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n364), .A2(new_n369), .ZN(new_n1038));
  OAI211_X1 g852(.A(new_n1025), .B(new_n1038), .C1(new_n908), .C2(new_n914), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1033), .A2(new_n1034), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1039), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1037), .ZN(new_n1042));
  OAI21_X1  g856(.A(KEYINPUT127), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1040), .A2(new_n1043), .ZN(G57));
endmodule


