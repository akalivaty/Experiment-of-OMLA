//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI22_X1  g0023(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n224), .B1(new_n227), .B2(KEYINPUT65), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT64), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n228), .B(new_n230), .C1(KEYINPUT65), .C2(new_n227), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(new_n211), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n214), .B1(new_n217), .B2(new_n219), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n202), .A2(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n220), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n247), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT87), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G257), .A3(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G294), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  OAI211_X1 g0064(.A(G250), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n260), .A2(new_n261), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G1), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT5), .A2(G41), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT5), .A2(G41), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n266), .A2(new_n267), .B1(new_n275), .B2(G264), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n272), .A2(new_n267), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n276), .A2(G179), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G169), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(new_n276), .B2(new_n279), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n254), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n266), .A2(new_n267), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n275), .A2(G264), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n279), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G169), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n276), .A2(G179), .A3(new_n279), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(KEYINPUT87), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n215), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n209), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT22), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT22), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n259), .A2(new_n294), .A3(new_n209), .A4(G87), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT86), .B(KEYINPUT24), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G116), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(G20), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT23), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n209), .B2(G107), .ZN(new_n301));
  INV_X1    g0101(.A(G107), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(KEYINPUT23), .A3(G20), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n299), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n296), .A2(new_n297), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n297), .B1(new_n296), .B2(new_n304), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n291), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n291), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n256), .A2(G1), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n309), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT25), .A3(new_n302), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT25), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n309), .B2(G107), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n312), .A2(G107), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n283), .A2(new_n289), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n308), .A2(KEYINPUT71), .A3(new_n309), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT71), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(new_n313), .B2(new_n291), .ZN(new_n322));
  INV_X1    g0122(.A(G116), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n311), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n313), .A2(new_n323), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(G20), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n291), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT85), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT85), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n291), .A2(new_n331), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(G20), .B1(G33), .B2(G283), .ZN(new_n334));
  INV_X1    g0134(.A(G97), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(G33), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT20), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n291), .A2(new_n331), .A3(new_n328), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n331), .B1(new_n291), .B2(new_n328), .ZN(new_n339));
  OAI211_X1 g0139(.A(KEYINPUT20), .B(new_n336), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n327), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n272), .A2(G270), .A3(new_n274), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT84), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n272), .A2(KEYINPUT84), .A3(G270), .A4(new_n274), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n278), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n348));
  OAI211_X1 g0148(.A(G257), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n349));
  INV_X1    g0149(.A(G303), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n348), .B(new_n349), .C1(new_n350), .C2(new_n259), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n267), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n281), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n342), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT21), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n347), .A2(G179), .A3(new_n352), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n342), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n342), .A2(new_n353), .A3(KEYINPUT21), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n319), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(G20), .A2(G33), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n362), .ZN(new_n363));
  XOR2_X1   g0163(.A(KEYINPUT8), .B(G58), .Z(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT68), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT8), .B(G58), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT68), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n209), .A2(G33), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n363), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(new_n291), .B1(new_n202), .B2(new_n313), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT69), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n310), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n308), .A2(KEYINPUT69), .A3(new_n309), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n374), .A2(new_n375), .B1(new_n208), .B2(G20), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G50), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT9), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT73), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n259), .A2(G222), .A3(new_n262), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n259), .A2(G223), .A3(G1698), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n382), .B(new_n383), .C1(new_n222), .C2(new_n259), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n267), .ZN(new_n385));
  INV_X1    g0185(.A(G41), .ZN(new_n386));
  AOI21_X1  g0186(.A(G1), .B1(new_n386), .B2(new_n268), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(new_n274), .A3(G274), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n274), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(G226), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n385), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G200), .ZN(new_n395));
  INV_X1    g0195(.A(G190), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(new_n394), .ZN(new_n397));
  INV_X1    g0197(.A(new_n378), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n397), .B1(KEYINPUT9), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n381), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT10), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n395), .B2(KEYINPUT74), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n400), .B(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G179), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n385), .A2(new_n404), .A3(new_n393), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n394), .A2(new_n281), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n378), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n209), .A2(G33), .A3(G77), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n362), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n308), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n411), .A2(KEYINPUT11), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n208), .A2(G20), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n320), .A2(new_n322), .A3(G68), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n313), .A2(new_n220), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT12), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(KEYINPUT11), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n412), .A2(new_n414), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n388), .B1(new_n221), .B2(new_n391), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT75), .ZN(new_n421));
  OR2_X1    g0221(.A1(G226), .A2(G1698), .ZN(new_n422));
  INV_X1    g0222(.A(G232), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G1698), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n422), .B(new_n424), .C1(new_n263), .C2(new_n264), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G97), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n421), .B1(new_n427), .B2(new_n267), .ZN(new_n428));
  AOI211_X1 g0228(.A(KEYINPUT75), .B(new_n274), .C1(new_n425), .C2(new_n426), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n420), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT13), .ZN(new_n431));
  INV_X1    g0231(.A(new_n426), .ZN(new_n432));
  NOR2_X1   g0232(.A1(G226), .A2(G1698), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n423), .B2(G1698), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n432), .B1(new_n434), .B2(new_n259), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT75), .B1(new_n435), .B2(new_n274), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n427), .A2(new_n421), .A3(new_n267), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT13), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n439), .A3(new_n420), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n431), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT14), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(G169), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n441), .B2(new_n404), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n442), .B1(new_n441), .B2(G169), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n418), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n439), .B1(new_n438), .B2(new_n420), .ZN(new_n447));
  AOI211_X1 g0247(.A(KEYINPUT13), .B(new_n419), .C1(new_n436), .C2(new_n437), .ZN(new_n448));
  OAI21_X1  g0248(.A(G200), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n449), .A2(KEYINPUT76), .B1(new_n450), .B2(G190), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n431), .A2(new_n440), .A3(KEYINPUT76), .A4(G190), .ZN(new_n452));
  INV_X1    g0252(.A(new_n418), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n451), .A2(KEYINPUT77), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT77), .ZN(new_n456));
  INV_X1    g0256(.A(new_n454), .ZN(new_n457));
  INV_X1    g0257(.A(G200), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n431), .B2(new_n440), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT76), .ZN(new_n460));
  OAI22_X1  g0260(.A1(new_n459), .A2(new_n460), .B1(new_n441), .B2(new_n396), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n456), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n446), .B1(new_n455), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n313), .B1(new_n365), .B2(new_n368), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT69), .B1(new_n308), .B2(new_n309), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n313), .A2(new_n291), .A3(new_n373), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n413), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n369), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G58), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n220), .ZN(new_n471));
  OAI21_X1  g0271(.A(G20), .B1(new_n471), .B2(new_n201), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n362), .A2(G159), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n257), .A2(new_n209), .A3(new_n258), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT7), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n258), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n474), .B1(new_n479), .B2(G68), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n308), .B1(new_n480), .B2(KEYINPUT16), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT16), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n220), .B1(new_n477), .B2(new_n478), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(new_n474), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n469), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n274), .A2(G232), .A3(new_n390), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n388), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(G223), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n488));
  OAI211_X1 g0288(.A(G226), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G87), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n487), .B1(new_n267), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n492), .A2(G179), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(new_n281), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT18), .B1(new_n485), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n263), .A2(new_n264), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT7), .B1(new_n497), .B2(new_n209), .ZN(new_n498));
  INV_X1    g0298(.A(new_n478), .ZN(new_n499));
  OAI21_X1  g0299(.A(G68), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n474), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(KEYINPUT16), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n484), .A2(new_n502), .A3(new_n291), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n491), .A2(new_n267), .ZN(new_n504));
  INV_X1    g0304(.A(new_n487), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n396), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(G200), .B2(new_n492), .ZN(new_n507));
  INV_X1    g0307(.A(new_n464), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n376), .B2(new_n369), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n503), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT17), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n503), .A2(new_n509), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT18), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n492), .A2(G179), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n281), .B2(new_n492), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n503), .A2(new_n507), .A3(new_n509), .A4(KEYINPUT17), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n496), .A2(new_n512), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n423), .A2(new_n262), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n221), .A2(G1698), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n497), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n267), .B1(new_n259), .B2(G107), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n388), .B1(new_n223), .B2(new_n391), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n281), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT70), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n362), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n364), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g0332(.A(KEYINPUT15), .B(G87), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n533), .A2(new_n370), .B1(new_n209), .B2(new_n222), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n291), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n320), .A2(new_n322), .A3(G77), .A4(new_n413), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n313), .A2(new_n222), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n528), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n526), .A2(new_n404), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n528), .A2(KEYINPUT72), .A3(new_n538), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n527), .A2(G200), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n535), .A2(new_n537), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n526), .A2(G190), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(new_n536), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NOR4_X1   g0349(.A1(new_n408), .A2(new_n463), .A3(new_n519), .A4(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n309), .A2(G97), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n312), .B2(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n479), .A2(G107), .ZN(new_n553));
  AND2_X1   g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n554), .A2(new_n205), .B1(KEYINPUT78), .B2(KEYINPUT6), .ZN(new_n555));
  NOR2_X1   g0355(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(KEYINPUT6), .B2(new_n335), .ZN(new_n557));
  XNOR2_X1  g0357(.A(G97), .B(G107), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n555), .B(G20), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n362), .A2(G77), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n553), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT79), .B1(new_n561), .B2(new_n291), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n560), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n302), .B1(new_n477), .B2(new_n478), .ZN(new_n564));
  OAI211_X1 g0364(.A(KEYINPUT79), .B(new_n291), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n552), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G250), .A2(G1698), .ZN(new_n568));
  NAND2_X1  g0368(.A1(KEYINPUT4), .A2(G244), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(G1698), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n259), .A2(new_n570), .B1(G33), .B2(G283), .ZN(new_n571));
  OAI211_X1 g0371(.A(G244), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT80), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT80), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n571), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n267), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n272), .A2(G257), .A3(new_n274), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n279), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n281), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n274), .B1(new_n575), .B2(KEYINPUT80), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n581), .B1(new_n585), .B2(new_n578), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n404), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n567), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n579), .A2(new_n396), .A3(new_n582), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(G200), .B2(new_n586), .ZN(new_n590));
  INV_X1    g0390(.A(new_n552), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n291), .B1(new_n563), .B2(new_n564), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT79), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n591), .B1(new_n594), .B2(new_n565), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n286), .A2(G190), .ZN(new_n597));
  AOI21_X1  g0397(.A(G200), .B1(new_n276), .B2(new_n279), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n307), .B(new_n317), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n588), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n342), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n345), .A2(new_n346), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n602), .A2(new_n352), .A3(new_n279), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G190), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n601), .B(new_n604), .C1(new_n458), .C2(new_n603), .ZN(new_n605));
  OAI211_X1 g0405(.A(G244), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT83), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT83), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n259), .A2(new_n608), .A3(G244), .A4(G1698), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n259), .A2(G238), .A3(new_n262), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n607), .A2(new_n609), .A3(new_n298), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n267), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT81), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n268), .B2(G1), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n208), .A2(KEYINPUT81), .A3(G45), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n274), .A2(new_n614), .A3(G250), .A4(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n274), .A2(G274), .A3(new_n269), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT82), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT82), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n616), .A2(new_n620), .A3(new_n617), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n612), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G200), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n612), .A2(new_n622), .A3(G190), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n259), .A2(new_n209), .A3(G68), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT19), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n209), .B1(new_n426), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(G87), .B2(new_n206), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n370), .B2(new_n335), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n626), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n291), .B1(new_n313), .B2(new_n533), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n312), .A2(G87), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n624), .A2(new_n625), .A3(new_n634), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n267), .A2(new_n611), .B1(new_n619), .B2(new_n621), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n404), .ZN(new_n637));
  INV_X1    g0437(.A(new_n533), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n312), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n637), .B(new_n640), .C1(G169), .C2(new_n636), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n605), .A2(new_n635), .A3(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n361), .A2(new_n550), .A3(new_n600), .A4(new_n642), .ZN(G372));
  NAND2_X1  g0443(.A1(new_n359), .A2(new_n358), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT21), .B1(new_n342), .B2(new_n353), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT90), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT90), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n356), .A2(new_n647), .A3(new_n358), .A4(new_n359), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n318), .B1(new_n282), .B2(new_n280), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT89), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n588), .A2(new_n596), .A3(new_n599), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n624), .A2(KEYINPUT88), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT88), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n623), .A2(new_n655), .A3(G200), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n654), .A2(new_n625), .A3(new_n634), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n641), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n652), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n594), .A2(new_n565), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(new_n552), .B1(new_n404), .B2(new_n586), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n661), .A2(new_n584), .B1(new_n595), .B2(new_n590), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n640), .B1(new_n636), .B2(G169), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n623), .A2(G179), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n634), .A2(new_n625), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n655), .B1(new_n623), .B2(G200), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n665), .B1(new_n668), .B2(new_n656), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n662), .A2(new_n669), .A3(KEYINPUT89), .A4(new_n599), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n651), .A2(new_n659), .A3(new_n670), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n567), .A2(new_n584), .A3(new_n587), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n641), .A2(new_n635), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT26), .B1(new_n588), .B2(new_n675), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n674), .A2(new_n641), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n550), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n407), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT77), .B1(new_n451), .B2(new_n454), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n457), .A2(new_n461), .A3(new_n456), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n544), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(new_n446), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n512), .A2(new_n518), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n496), .B(new_n517), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n680), .B1(new_n688), .B2(new_n403), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n679), .A2(new_n689), .ZN(G369));
  INV_X1    g0490(.A(new_n360), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G343), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT91), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n601), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n605), .B1(new_n691), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n649), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n319), .A2(new_n698), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n283), .A2(new_n289), .A3(new_n318), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n318), .A2(new_n698), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n599), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n702), .A2(G330), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n360), .A2(new_n699), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n706), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n650), .A2(new_n698), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n708), .A2(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n212), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n208), .ZN(new_n716));
  INV_X1    g0516(.A(G87), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n205), .A2(new_n717), .A3(new_n323), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT92), .Z(new_n719));
  INV_X1    g0519(.A(new_n219), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n716), .A2(new_n719), .B1(new_n720), .B2(new_n715), .ZN(new_n721));
  XNOR2_X1  g0521(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G330), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n586), .A2(new_n276), .A3(new_n636), .ZN(new_n726));
  INV_X1    g0526(.A(new_n357), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n603), .A2(new_n636), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(new_n404), .A3(new_n286), .A4(new_n583), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n636), .A2(new_n276), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n357), .A3(KEYINPUT30), .A4(new_n586), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n728), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n733), .B2(new_n698), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n600), .A2(new_n361), .A3(new_n642), .A4(new_n699), .ZN(new_n737));
  AOI211_X1 g0537(.A(KEYINPUT94), .B(new_n724), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT94), .ZN(new_n739));
  INV_X1    g0539(.A(new_n735), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n737), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n739), .B1(new_n742), .B2(G330), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT95), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n678), .B2(new_n699), .ZN(new_n747));
  AOI211_X1 g0547(.A(KEYINPUT95), .B(new_n698), .C1(new_n671), .C2(new_n677), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(KEYINPUT26), .B1(new_n658), .B2(new_n588), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n672), .A2(new_n673), .A3(new_n635), .A4(new_n641), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(new_n641), .A3(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n361), .A2(new_n653), .A3(new_n658), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n699), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(new_n745), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n744), .B1(new_n749), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n723), .B1(new_n756), .B2(G1), .ZN(G364));
  AND2_X1   g0557(.A1(new_n209), .A2(G13), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G45), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n759), .A2(KEYINPUT96), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(KEYINPUT96), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n760), .A2(G1), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n715), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n215), .B1(G20), .B2(new_n281), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n209), .A2(new_n404), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n396), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(KEYINPUT98), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n769), .A2(KEYINPUT98), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G50), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n768), .A2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n209), .A2(G179), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n776), .A2(new_n220), .B1(new_n778), .B2(new_n717), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n396), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n209), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n777), .A2(new_n396), .A3(G200), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n335), .B1(new_n782), .B2(new_n302), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n777), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G159), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT32), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n767), .A2(G190), .A3(new_n458), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n259), .B1(new_n790), .B2(new_n470), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n767), .A2(new_n785), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n791), .B1(G77), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n774), .A2(new_n784), .A3(new_n789), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n773), .A2(G326), .ZN(new_n796));
  INV_X1    g0596(.A(G322), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n790), .A2(new_n797), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n786), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n259), .B(new_n799), .C1(G329), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n781), .ZN(new_n802));
  INV_X1    g0602(.A(new_n778), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n802), .A2(G294), .B1(new_n803), .B2(G303), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT33), .B(G317), .ZN(new_n805));
  INV_X1    g0605(.A(new_n782), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n775), .A2(new_n805), .B1(new_n806), .B2(G283), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n796), .A2(new_n801), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n766), .B1(new_n795), .B2(new_n808), .ZN(new_n809));
  OR3_X1    g0609(.A1(KEYINPUT97), .A2(G13), .A3(G33), .ZN(new_n810));
  OAI21_X1  g0610(.A(KEYINPUT97), .B1(G13), .B2(G33), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(G20), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n765), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n714), .A2(new_n497), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n816), .A2(G355), .B1(new_n323), .B2(new_n714), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n714), .A2(new_n259), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(G45), .B2(new_n219), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n252), .A2(new_n268), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n764), .B(new_n809), .C1(new_n815), .C2(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT99), .Z(new_n823));
  INV_X1    g0623(.A(new_n814), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n702), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n763), .B1(new_n702), .B2(G330), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(G330), .B2(new_n702), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NAND2_X1  g0629(.A1(new_n698), .A2(new_n538), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n548), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n544), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT103), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT103), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n544), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n833), .B(new_n835), .C1(new_n544), .C2(new_n830), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n747), .B2(new_n748), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n833), .A2(new_n835), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n678), .A2(new_n699), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n744), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n763), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n813), .A2(new_n766), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n763), .B1(G77), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n773), .A2(G137), .B1(G150), .B2(new_n775), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT101), .ZN(new_n848));
  XNOR2_X1  g0648(.A(KEYINPUT102), .B(G143), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n787), .B2(new_n792), .C1(new_n790), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT34), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n782), .A2(new_n220), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n497), .B(new_n852), .C1(G132), .C2(new_n800), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n802), .A2(G58), .B1(new_n803), .B2(G50), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n775), .A2(G283), .B1(new_n793), .B2(G116), .ZN(new_n856));
  INV_X1    g0656(.A(new_n773), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n350), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT100), .ZN(new_n859));
  INV_X1    g0659(.A(G294), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n497), .B1(new_n790), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G311), .B2(new_n800), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n802), .A2(G97), .B1(new_n806), .B2(G87), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n862), .B(new_n863), .C1(new_n302), .C2(new_n778), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n855), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n846), .B1(new_n865), .B2(new_n765), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n813), .B2(new_n836), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n844), .A2(new_n867), .ZN(G384));
  NOR2_X1   g0668(.A1(new_n217), .A2(new_n323), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT35), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n871), .B2(new_n870), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT36), .ZN(new_n874));
  OR3_X1    g0674(.A1(new_n219), .A2(new_n222), .A3(new_n471), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n208), .B(G13), .C1(new_n875), .C2(new_n248), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT105), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT104), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n483), .B2(new_n474), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n500), .A2(KEYINPUT104), .A3(new_n501), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(new_n482), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n469), .B1(new_n882), .B2(new_n481), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n510), .B1(new_n883), .B2(new_n495), .ZN(new_n884));
  INV_X1    g0684(.A(new_n695), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n513), .A2(new_n516), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n513), .A2(new_n695), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .A4(new_n510), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n519), .A2(new_n886), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n892), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n698), .A2(new_n418), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n463), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n446), .B(new_n899), .C1(new_n455), .C2(new_n462), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI221_X4 g0703(.A(new_n698), .B1(new_n833), .B2(new_n835), .C1(new_n671), .C2(new_n677), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n544), .A2(new_n698), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n898), .B(new_n903), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n496), .A2(new_n517), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n885), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n878), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n446), .A2(new_n698), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT106), .Z(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n892), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n892), .B2(new_n893), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT39), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n510), .B1(new_n485), .B2(new_n495), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n485), .A2(new_n885), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT37), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n891), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n519), .A2(new_n917), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n895), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n922), .A2(KEYINPUT107), .A3(new_n923), .A4(new_n897), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n915), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT39), .B1(new_n921), .B2(new_n895), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT107), .B1(new_n926), .B2(new_n897), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT108), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n897), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT107), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT108), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(new_n932), .A3(new_n924), .A4(new_n915), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n912), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n909), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n906), .A2(new_n878), .A3(new_n908), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n749), .A2(new_n550), .A3(new_n755), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n689), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n938), .B(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n902), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n899), .B1(new_n683), .B2(new_n446), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n742), .B(new_n836), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n922), .A2(new_n897), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT40), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n913), .A2(new_n914), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n948), .B1(new_n944), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n903), .A2(new_n898), .A3(new_n742), .A4(new_n836), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT109), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n953), .A3(new_n948), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n947), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n955), .A2(new_n550), .A3(new_n742), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n955), .B1(new_n550), .B2(new_n742), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n956), .A2(new_n957), .A3(new_n724), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n941), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT110), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n960), .B1(new_n208), .B2(new_n758), .C1(new_n941), .C2(new_n958), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n959), .A2(KEYINPUT110), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n877), .B1(new_n961), .B2(new_n962), .ZN(G367));
  INV_X1    g0763(.A(new_n818), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n238), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n815), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n714), .B2(new_n638), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n764), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n658), .B1(new_n634), .B2(new_n699), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n699), .A2(new_n634), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n641), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n849), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n773), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(G137), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n792), .A2(new_n202), .B1(new_n786), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n790), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n497), .B(new_n977), .C1(G150), .C2(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n775), .A2(G159), .B1(new_n806), .B2(G77), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n802), .A2(G68), .B1(new_n803), .B2(G58), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n975), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n782), .A2(new_n335), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G107), .B2(new_n802), .ZN(new_n984));
  XNOR2_X1  g0784(.A(KEYINPUT111), .B(G311), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n984), .B1(new_n860), .B2(new_n776), .C1(new_n857), .C2(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G283), .A2(new_n793), .B1(new_n800), .B2(G317), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n259), .B1(new_n978), .B2(G303), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT46), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n778), .B2(new_n323), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n803), .A2(KEYINPUT46), .A3(G116), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n987), .A2(new_n988), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n982), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT47), .Z(new_n994));
  OAI221_X1 g0794(.A(new_n968), .B1(new_n973), .B2(new_n824), .C1(new_n766), .C2(new_n994), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n588), .B(new_n596), .C1(new_n595), .C2(new_n699), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(new_n704), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n698), .B1(new_n997), .B2(new_n588), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n672), .A2(new_n698), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n710), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n998), .B1(new_n1001), .B2(KEYINPUT42), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(KEYINPUT42), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1002), .A2(new_n1003), .B1(KEYINPUT43), .B2(new_n973), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1000), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n708), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1006), .B(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n712), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1011), .B1(new_n1012), .B2(new_n1007), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n712), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(KEYINPUT44), .A3(new_n1007), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT44), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n712), .B2(new_n1000), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n708), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1015), .A2(new_n708), .A3(new_n1019), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n702), .A2(G330), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n703), .A2(new_n709), .A3(new_n706), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n706), .B2(new_n709), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1025), .B(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n756), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n715), .B(KEYINPUT41), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n762), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n995), .B1(new_n1010), .B2(new_n1031), .ZN(G387));
  INV_X1    g0832(.A(new_n1028), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n818), .B1(new_n242), .B2(new_n268), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n816), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n719), .B2(new_n1035), .ZN(new_n1036));
  OR3_X1    g0836(.A1(new_n366), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1037));
  OAI21_X1  g0837(.A(KEYINPUT50), .B1(new_n366), .B2(G50), .ZN(new_n1038));
  AOI21_X1  g0838(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n719), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1036), .A2(new_n1040), .B1(new_n302), .B2(new_n714), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n763), .B1(new_n1041), .B2(new_n966), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n978), .A2(G317), .B1(new_n793), .B2(G303), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n776), .B2(new_n985), .C1(new_n857), .C2(new_n797), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n802), .A2(G283), .B1(new_n803), .B2(G294), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n782), .A2(new_n323), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n259), .B(new_n1053), .C1(G326), .C2(new_n800), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n857), .A2(new_n787), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n790), .A2(new_n202), .B1(new_n792), .B2(new_n220), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n497), .B(new_n1057), .C1(G150), .C2(new_n800), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n778), .A2(new_n222), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n983), .B(new_n1059), .C1(new_n638), .C2(new_n802), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n468), .A2(new_n775), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1055), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1042), .B1(new_n1063), .B2(new_n765), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n703), .A2(new_n706), .A3(new_n814), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1033), .A2(new_n762), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n749), .A2(new_n755), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n842), .A3(new_n1033), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n715), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n756), .A2(new_n1033), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(G393));
  OR2_X1    g0871(.A1(new_n1068), .A2(new_n1024), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1068), .A2(new_n1024), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1072), .A2(new_n715), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1022), .A2(new_n762), .A3(new_n1023), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n815), .B1(new_n335), .B2(new_n212), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n964), .A2(new_n246), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n763), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n773), .A2(G150), .B1(G159), .B2(new_n978), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT51), .Z(new_n1080));
  AOI21_X1  g0880(.A(new_n497), .B1(new_n800), .B2(new_n974), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n220), .B2(new_n778), .C1(new_n717), .C2(new_n782), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT112), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n792), .A2(new_n366), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n781), .A2(new_n222), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(G50), .C2(new_n775), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1080), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1087), .A2(KEYINPUT113), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n773), .A2(G317), .B1(G311), .B2(new_n978), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n497), .B1(new_n786), .B2(new_n797), .C1(new_n860), .C2(new_n792), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n776), .A2(new_n350), .B1(new_n302), .B2(new_n782), .ZN(new_n1092));
  INV_X1    g0892(.A(G283), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n781), .A2(new_n323), .B1(new_n778), .B2(new_n1093), .ZN(new_n1094));
  OR4_X1    g0894(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1087), .A2(KEYINPUT113), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1088), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1078), .B1(new_n1097), .B2(new_n765), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n824), .B2(new_n1000), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1074), .A2(new_n1075), .A3(new_n1099), .ZN(G390));
  INV_X1    g0900(.A(new_n905), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n754), .B2(new_n837), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n903), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n912), .A2(new_n1103), .A3(new_n945), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n928), .A2(new_n933), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n840), .A2(new_n1101), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n911), .B1(new_n1106), .B2(new_n903), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1104), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n903), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n742), .A2(G330), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n837), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1111), .A2(KEYINPUT114), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n743), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n724), .B1(new_n736), .B2(new_n737), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n739), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1114), .A2(new_n1116), .A3(new_n836), .A4(new_n903), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1110), .A2(KEYINPUT114), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1104), .B1(new_n1117), .B2(new_n1118), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n762), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n763), .B1(new_n468), .B2(new_n845), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n802), .A2(G159), .B1(new_n793), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n976), .B2(new_n776), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT115), .Z(new_n1128));
  NAND2_X1  g0928(.A1(new_n773), .A2(G128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n806), .A2(G50), .ZN(new_n1130));
  INV_X1    g0930(.A(G132), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n790), .A2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n497), .B(new_n1132), .C1(G125), .C2(new_n800), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1129), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n803), .A2(G150), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1128), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1137), .A2(KEYINPUT116), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(KEYINPUT116), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n497), .B1(new_n778), .B2(new_n717), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n773), .A2(G283), .B1(KEYINPUT117), .B2(new_n1140), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n790), .A2(new_n323), .B1(new_n786), .B2(new_n860), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G97), .B2(new_n793), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n852), .B(new_n1085), .C1(G107), .C2(new_n775), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1140), .A2(KEYINPUT117), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1138), .A2(new_n1139), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1123), .B1(new_n1147), .B2(new_n765), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n1105), .B2(new_n813), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n550), .A2(new_n1115), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n939), .A2(new_n689), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1115), .A2(new_n836), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1102), .B1(new_n1109), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1117), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1114), .A2(new_n1116), .A3(new_n836), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1111), .B1(new_n1155), .B2(new_n1109), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1106), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1154), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1151), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n715), .B1(new_n1121), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1113), .A2(new_n1119), .A3(new_n1151), .A4(new_n1158), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1122), .B(new_n1149), .C1(new_n1161), .C2(new_n1163), .ZN(G378));
  INV_X1    g0964(.A(new_n947), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n954), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n953), .B1(new_n952), .B2(new_n948), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1165), .B(G330), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n398), .A2(new_n885), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n408), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n403), .B(new_n407), .C1(new_n398), .C2(new_n885), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1168), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n955), .B2(G330), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n938), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1168), .A2(new_n1177), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n955), .A2(G330), .A3(new_n1179), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1182), .A2(new_n1183), .A3(new_n937), .A4(new_n935), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1177), .A2(new_n812), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n763), .B1(G50), .B2(new_n845), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(G33), .A2(G41), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G50), .B(new_n1188), .C1(new_n497), .C2(new_n386), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n773), .A2(G116), .B1(G68), .B2(new_n802), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT118), .Z(new_n1191));
  OAI22_X1  g0991(.A1(new_n790), .A2(new_n302), .B1(new_n786), .B2(new_n1093), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n386), .B(new_n497), .C1(new_n792), .C2(new_n533), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1059), .B1(G97), .B2(new_n775), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n470), .B2(new_n782), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1189), .B1(new_n1196), .B2(KEYINPUT58), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n802), .A2(G150), .B1(new_n793), .B2(G137), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1131), .B2(new_n776), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G128), .A2(new_n978), .B1(new_n803), .B2(new_n1125), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT119), .Z(new_n1201));
  AOI211_X1 g1001(.A(new_n1199), .B(new_n1201), .C1(G125), .C2(new_n773), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT59), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1205));
  INV_X1    g1005(.A(G124), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1188), .B1(new_n786), .B2(new_n1206), .C1(new_n787), .C2(new_n782), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT120), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1204), .A2(new_n1205), .A3(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1197), .B(new_n1209), .C1(KEYINPUT58), .C2(new_n1196), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1187), .B1(new_n1210), .B2(new_n765), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1185), .A2(new_n762), .B1(new_n1186), .B2(new_n1211), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1181), .A2(new_n1184), .B1(new_n1162), .B2(new_n1151), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n715), .B1(new_n1213), .B2(KEYINPUT57), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1162), .A2(new_n1151), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1185), .A2(KEYINPUT57), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1212), .B1(new_n1214), .B2(new_n1216), .ZN(G375));
  XOR2_X1   g1017(.A(new_n762), .B(KEYINPUT121), .Z(new_n1218));
  NAND2_X1  g1018(.A1(new_n1109), .A2(new_n812), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n763), .B1(G68), .B2(new_n845), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n773), .A2(G132), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT123), .Z(new_n1222));
  AOI22_X1  g1022(.A1(new_n802), .A2(G50), .B1(new_n803), .B2(G159), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n775), .A2(new_n1125), .B1(new_n806), .B2(G58), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n497), .B1(new_n978), .B2(G137), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G150), .A2(new_n793), .B1(new_n800), .B2(G128), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n497), .B1(new_n782), .B2(new_n222), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT122), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n773), .A2(G294), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n790), .A2(new_n1093), .B1(new_n792), .B2(new_n302), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G303), .B2(new_n800), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n803), .A2(G97), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n638), .A2(new_n802), .B1(new_n775), .B2(G116), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1230), .A2(new_n1232), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n1222), .A2(new_n1227), .B1(new_n1229), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1220), .B1(new_n1236), .B2(new_n765), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1158), .A2(new_n1218), .B1(new_n1219), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1159), .A2(new_n1030), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1151), .A2(new_n1158), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(G381));
  AND3_X1   g1041(.A1(new_n1074), .A2(new_n1075), .A3(new_n1099), .ZN(new_n1242));
  INV_X1    g1042(.A(G384), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  OR4_X1    g1044(.A1(G396), .A2(new_n1244), .A3(G393), .A4(G381), .ZN(new_n1245));
  OR4_X1    g1045(.A1(G387), .A2(new_n1245), .A3(G375), .A4(G378), .ZN(G407));
  INV_X1    g1046(.A(G343), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(G213), .ZN(new_n1248));
  OR3_X1    g1048(.A1(G375), .A2(G378), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(G213), .A3(new_n1249), .ZN(G409));
  OAI211_X1 g1050(.A(G390), .B(new_n995), .C1(new_n1031), .C2(new_n1010), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1242), .A2(G387), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G393), .B(new_n828), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1251), .A2(new_n1252), .A3(new_n1254), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1256), .A2(KEYINPUT126), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT126), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G378), .B(new_n1212), .C1(new_n1214), .C2(new_n1216), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n762), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1149), .B1(new_n1120), .B2(new_n1262), .ZN(new_n1263));
  AOI211_X1 g1063(.A(G41), .B(new_n714), .C1(new_n1120), .C2(new_n1159), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n1162), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1213), .A2(new_n1030), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1185), .A2(new_n1218), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1186), .A2(new_n1211), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1265), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1261), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT124), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1151), .B2(new_n1158), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n939), .A2(new_n689), .A3(new_n1150), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n903), .B1(new_n744), .B2(new_n836), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1106), .B1(new_n1276), .B2(new_n1111), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1275), .A2(new_n1277), .A3(KEYINPUT60), .A4(new_n1154), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1274), .A2(new_n715), .A3(new_n1159), .A4(new_n1278), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1279), .A2(G384), .A3(new_n1238), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G384), .B1(new_n1279), .B2(new_n1238), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1272), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(new_n1238), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1243), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1279), .A2(G384), .A3(new_n1238), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(KEYINPUT124), .A3(new_n1285), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1282), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1271), .A2(new_n1287), .A3(new_n1288), .A4(new_n1248), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1261), .A2(new_n1270), .B1(G213), .B2(new_n1247), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1247), .A2(G213), .A3(G2897), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1282), .A2(new_n1286), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1294), .B1(new_n1295), .B2(new_n1293), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1289), .B(new_n1290), .C1(new_n1291), .C2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1288), .B1(new_n1291), .B2(new_n1287), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1260), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1256), .A2(new_n1257), .A3(new_n1290), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT125), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1300), .B(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1291), .A2(new_n1287), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OR2_X1    g1105(.A1(new_n1296), .A2(new_n1291), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1291), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1302), .A2(new_n1305), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1299), .A2(new_n1308), .ZN(G405));
  NAND2_X1  g1109(.A1(G375), .A2(new_n1265), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT127), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n1311), .A3(new_n1261), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(G375), .A2(KEYINPUT127), .A3(new_n1265), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1312), .A2(new_n1295), .A3(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1292), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1314), .A2(new_n1315), .A3(new_n1260), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1292), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1261), .A2(new_n1311), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1185), .A2(new_n1215), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT57), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1213), .A2(KEYINPUT57), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(new_n715), .A3(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(G378), .B1(new_n1324), .B2(new_n1212), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1319), .A2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1313), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1318), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1312), .A2(new_n1295), .A3(new_n1313), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1317), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1316), .A2(new_n1330), .ZN(G402));
endmodule


