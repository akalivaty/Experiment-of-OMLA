

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774;

  AND2_X2 U371 ( .A1(n380), .A2(n416), .ZN(n687) );
  XNOR2_X1 U372 ( .A(n585), .B(KEYINPUT0), .ZN(n620) );
  NAND2_X1 U373 ( .A1(n584), .A2(n419), .ZN(n585) );
  NOR2_X1 U374 ( .A1(G953), .A2(G237), .ZN(n469) );
  XNOR2_X1 U375 ( .A(KEYINPUT74), .B(G110), .ZN(n762) );
  XNOR2_X1 U376 ( .A(n349), .B(n761), .ZN(n642) );
  XNOR2_X1 U377 ( .A(n451), .B(n450), .ZN(n349) );
  NAND2_X2 U378 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X2 U379 ( .A(n508), .B(n397), .ZN(n666) );
  INV_X1 U380 ( .A(G953), .ZN(n446) );
  NOR2_X1 U381 ( .A1(n721), .A2(n587), .ZN(n350) );
  NOR2_X2 U382 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X2 U383 ( .A(n616), .B(KEYINPUT6), .ZN(n587) );
  OR2_X1 U384 ( .A1(n588), .A2(n721), .ZN(n590) );
  NOR2_X1 U385 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U386 ( .A1(n646), .A2(n696), .ZN(n647) );
  NAND2_X1 U387 ( .A1(n377), .A2(n657), .ZN(n637) );
  AND2_X1 U388 ( .A1(n387), .A2(n386), .ZN(n385) );
  AND2_X1 U389 ( .A1(n392), .A2(n594), .ZN(n708) );
  XNOR2_X1 U390 ( .A(n512), .B(n511), .ZN(n586) );
  OR2_X1 U391 ( .A1(n552), .A2(n528), .ZN(n540) );
  XNOR2_X1 U392 ( .A(n673), .B(n672), .ZN(n674) );
  OR2_X1 U393 ( .A1(n479), .A2(n487), .ZN(n480) );
  OR2_X1 U394 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U395 ( .A(n455), .B(n454), .ZN(n472) );
  XNOR2_X1 U396 ( .A(KEYINPUT3), .B(G119), .ZN(n454) );
  XNOR2_X1 U397 ( .A(G113), .B(G101), .ZN(n455) );
  XNOR2_X2 U398 ( .A(n351), .B(n485), .ZN(n602) );
  NAND2_X1 U399 ( .A1(n688), .A2(n573), .ZN(n351) );
  NAND2_X1 U400 ( .A1(n353), .A2(n352), .ZN(n688) );
  NAND2_X1 U401 ( .A1(n396), .A2(n654), .ZN(n352) );
  NAND2_X1 U402 ( .A1(n370), .A2(n371), .ZN(n353) );
  XNOR2_X2 U403 ( .A(n655), .B(G146), .ZN(n508) );
  XNOR2_X2 U404 ( .A(n468), .B(n467), .ZN(n655) );
  XNOR2_X2 U405 ( .A(n443), .B(KEYINPUT4), .ZN(n468) );
  BUF_X1 U406 ( .A(n549), .Z(n354) );
  BUF_X1 U407 ( .A(n666), .Z(n355) );
  XNOR2_X2 U408 ( .A(n463), .B(KEYINPUT38), .ZN(n737) );
  XNOR2_X1 U409 ( .A(n394), .B(n393), .ZN(n774) );
  OR2_X1 U410 ( .A1(n753), .A2(n536), .ZN(n394) );
  NOR2_X2 U411 ( .A1(n666), .A2(G902), .ZN(n357) );
  INV_X1 U412 ( .A(n603), .ZN(n356) );
  XNOR2_X2 U413 ( .A(n357), .B(n358), .ZN(n515) );
  XOR2_X1 U414 ( .A(KEYINPUT92), .B(G472), .Z(n358) );
  NAND2_X1 U415 ( .A1(n402), .A2(n377), .ZN(n401) );
  XNOR2_X1 U416 ( .A(n570), .B(KEYINPUT81), .ZN(n402) );
  BUF_X1 U417 ( .A(n586), .Z(n722) );
  XNOR2_X2 U418 ( .A(G143), .B(G128), .ZN(n443) );
  INV_X1 U419 ( .A(n716), .ZN(n391) );
  NAND2_X1 U420 ( .A1(n708), .A2(n389), .ZN(n386) );
  NAND2_X1 U421 ( .A1(n607), .A2(n664), .ZN(n375) );
  NAND2_X1 U422 ( .A1(n409), .A2(G234), .ZN(n408) );
  INV_X1 U423 ( .A(G953), .ZN(n409) );
  XNOR2_X1 U424 ( .A(KEYINPUT96), .B(KEYINPUT12), .ZN(n420) );
  NAND2_X1 U425 ( .A1(G234), .A2(G237), .ZN(n490) );
  XNOR2_X1 U426 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n444) );
  XNOR2_X1 U427 ( .A(n762), .B(KEYINPUT70), .ZN(n505) );
  XNOR2_X1 U428 ( .A(n457), .B(n458), .ZN(n761) );
  XOR2_X1 U429 ( .A(KEYINPUT73), .B(KEYINPUT16), .Z(n456) );
  NAND2_X1 U430 ( .A1(n366), .A2(n417), .ZN(n414) );
  INV_X1 U431 ( .A(KEYINPUT75), .ZN(n376) );
  NAND2_X1 U432 ( .A1(n350), .A2(n356), .ZN(n378) );
  INV_X1 U433 ( .A(KEYINPUT19), .ZN(n535) );
  INV_X1 U434 ( .A(KEYINPUT68), .ZN(n389) );
  XOR2_X1 U435 ( .A(n525), .B(KEYINPUT46), .Z(n526) );
  XNOR2_X1 U436 ( .A(KEYINPUT83), .B(KEYINPUT48), .ZN(n556) );
  INV_X1 U437 ( .A(G221), .ZN(n487) );
  XNOR2_X1 U438 ( .A(n482), .B(KEYINPUT20), .ZN(n486) );
  XNOR2_X1 U439 ( .A(KEYINPUT91), .B(KEYINPUT5), .ZN(n471) );
  NAND2_X1 U440 ( .A1(n407), .A2(G234), .ZN(n410) );
  NAND2_X1 U441 ( .A1(n408), .A2(KEYINPUT8), .ZN(n411) );
  NOR2_X1 U442 ( .A1(KEYINPUT8), .A2(G953), .ZN(n407) );
  XOR2_X1 U443 ( .A(G140), .B(KEYINPUT95), .Z(n427) );
  XNOR2_X1 U444 ( .A(G113), .B(KEYINPUT94), .ZN(n426) );
  XNOR2_X1 U445 ( .A(G131), .B(G143), .ZN(n421) );
  XNOR2_X1 U446 ( .A(G131), .B(G134), .ZN(n467) );
  XNOR2_X1 U447 ( .A(n473), .B(G140), .ZN(n500) );
  XOR2_X1 U448 ( .A(G122), .B(G104), .Z(n452) );
  XOR2_X1 U449 ( .A(G116), .B(G107), .Z(n453) );
  INV_X1 U450 ( .A(G237), .ZN(n460) );
  INV_X1 U451 ( .A(G902), .ZN(n573) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n470), .B(n471), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n472), .B(n360), .ZN(n399) );
  XOR2_X1 U455 ( .A(KEYINPUT78), .B(G104), .Z(n499) );
  XNOR2_X1 U456 ( .A(G101), .B(G107), .ZN(n498) );
  NAND2_X1 U457 ( .A1(n412), .A2(n366), .ZN(n416) );
  INV_X1 U458 ( .A(n637), .ZN(n373) );
  NOR2_X1 U459 ( .A1(n740), .A2(n741), .ZN(n466) );
  XNOR2_X1 U460 ( .A(n433), .B(n432), .ZN(n552) );
  XNOR2_X1 U461 ( .A(n431), .B(G475), .ZN(n432) );
  XNOR2_X1 U462 ( .A(n679), .B(n678), .ZN(n680) );
  AND2_X1 U463 ( .A1(n414), .A2(G210), .ZN(n413) );
  NAND2_X1 U464 ( .A1(n637), .A2(n366), .ZN(n415) );
  INV_X1 U465 ( .A(KEYINPUT42), .ZN(n393) );
  AND2_X1 U466 ( .A1(n587), .A2(n543), .ZN(n544) );
  NAND2_X1 U467 ( .A1(n359), .A2(n594), .ZN(n596) );
  XNOR2_X1 U468 ( .A(n379), .B(n367), .ZN(n664) );
  XNOR2_X1 U469 ( .A(KEYINPUT53), .B(KEYINPUT117), .ZN(n403) );
  NAND2_X1 U470 ( .A1(n760), .A2(n405), .ZN(n404) );
  AND2_X1 U471 ( .A1(n759), .A2(n446), .ZN(n405) );
  XOR2_X1 U472 ( .A(n593), .B(KEYINPUT34), .Z(n359) );
  XOR2_X1 U473 ( .A(G137), .B(G116), .Z(n360) );
  XOR2_X1 U474 ( .A(KEYINPUT93), .B(KEYINPUT11), .Z(n361) );
  AND2_X1 U475 ( .A1(n709), .A2(n541), .ZN(n362) );
  NOR2_X1 U476 ( .A1(n740), .A2(n599), .ZN(n363) );
  AND2_X1 U477 ( .A1(n415), .A2(n413), .ZN(n364) );
  XOR2_X1 U478 ( .A(KEYINPUT71), .B(KEYINPUT39), .Z(n365) );
  NAND2_X1 U479 ( .A1(n639), .A2(KEYINPUT2), .ZN(n366) );
  XOR2_X1 U480 ( .A(n604), .B(KEYINPUT32), .Z(n367) );
  INV_X1 U481 ( .A(n418), .ZN(n417) );
  BUF_X1 U482 ( .A(n686), .Z(n368) );
  XNOR2_X1 U483 ( .A(n395), .B(n524), .ZN(n686) );
  BUF_X1 U484 ( .A(n515), .Z(n728) );
  BUF_X1 U485 ( .A(n687), .Z(n369) );
  INV_X1 U486 ( .A(n638), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n726), .B(KEYINPUT90), .ZN(n599) );
  INV_X1 U488 ( .A(n396), .ZN(n370) );
  INV_X1 U489 ( .A(n654), .ZN(n371) );
  XNOR2_X1 U490 ( .A(n474), .B(n500), .ZN(n654) );
  BUF_X1 U491 ( .A(n523), .Z(n372) );
  OR2_X2 U492 ( .A1(n510), .A2(n547), .ZN(n536) );
  OR2_X2 U493 ( .A1(n742), .A2(n704), .ZN(n538) );
  XNOR2_X1 U494 ( .A(n522), .B(n521), .ZN(n549) );
  NAND2_X1 U495 ( .A1(n373), .A2(n418), .ZN(n412) );
  XNOR2_X2 U496 ( .A(n374), .B(n534), .ZN(n542) );
  NAND2_X1 U497 ( .A1(n533), .A2(n736), .ZN(n374) );
  INV_X1 U498 ( .A(n375), .ZN(n611) );
  NAND2_X1 U499 ( .A1(n608), .A2(n375), .ZN(n613) );
  XNOR2_X1 U500 ( .A(n404), .B(n403), .ZN(G75) );
  OR2_X1 U501 ( .A1(n719), .A2(n637), .ZN(n759) );
  INV_X1 U502 ( .A(n380), .ZN(n719) );
  XNOR2_X2 U503 ( .A(n401), .B(n376), .ZN(n380) );
  NAND2_X1 U504 ( .A1(n549), .A2(n737), .ZN(n400) );
  NAND2_X1 U505 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X2 U506 ( .A(n590), .B(n589), .ZN(n752) );
  NAND2_X1 U507 ( .A1(n377), .A2(n446), .ZN(n765) );
  XNOR2_X2 U508 ( .A(n635), .B(KEYINPUT45), .ZN(n377) );
  OR2_X1 U509 ( .A1(n626), .A2(n603), .ZN(n606) );
  NOR2_X1 U510 ( .A1(n626), .A2(n378), .ZN(n379) );
  NAND2_X1 U511 ( .A1(n364), .A2(n380), .ZN(n644) );
  NAND2_X1 U512 ( .A1(n390), .A2(n716), .ZN(n388) );
  XNOR2_X2 U513 ( .A(n538), .B(n537), .ZN(n390) );
  NAND2_X1 U514 ( .A1(n384), .A2(n381), .ZN(n383) );
  NOR2_X1 U515 ( .A1(n382), .A2(n708), .ZN(n381) );
  INV_X1 U516 ( .A(n390), .ZN(n382) );
  NAND2_X1 U517 ( .A1(n385), .A2(n383), .ZN(n554) );
  NOR2_X1 U518 ( .A1(n391), .A2(n389), .ZN(n384) );
  NAND2_X1 U519 ( .A1(n388), .A2(n389), .ZN(n387) );
  XNOR2_X1 U520 ( .A(n550), .B(KEYINPUT105), .ZN(n392) );
  XNOR2_X1 U521 ( .A(n466), .B(n465), .ZN(n753) );
  NOR2_X2 U522 ( .A1(n686), .A2(n774), .ZN(n527) );
  NAND2_X1 U523 ( .A1(n523), .A2(n531), .ZN(n395) );
  XNOR2_X2 U524 ( .A(n400), .B(n365), .ZN(n523) );
  XNOR2_X1 U525 ( .A(n481), .B(n480), .ZN(n396) );
  INV_X1 U526 ( .A(n372), .ZN(n568) );
  OR2_X1 U527 ( .A1(n719), .A2(n718), .ZN(n758) );
  XNOR2_X1 U528 ( .A(n406), .B(G128), .ZN(n477) );
  XNOR2_X2 U529 ( .A(G110), .B(KEYINPUT23), .ZN(n406) );
  NAND2_X1 U530 ( .A1(n411), .A2(n410), .ZN(n479) );
  XNOR2_X1 U531 ( .A(n514), .B(n513), .ZN(n520) );
  INV_X1 U532 ( .A(n542), .ZN(n543) );
  XNOR2_X2 U533 ( .A(G146), .B(G125), .ZN(n445) );
  XNOR2_X2 U534 ( .A(G119), .B(KEYINPUT24), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n583), .A2(n582), .ZN(n419) );
  BUF_X1 U536 ( .A(n688), .Z(n689) );
  XNOR2_X1 U537 ( .A(n542), .B(n535), .ZN(n571) );
  OR2_X1 U538 ( .A1(n548), .A2(n721), .ZN(n716) );
  XNOR2_X1 U539 ( .A(n361), .B(n420), .ZN(n424) );
  NAND2_X1 U540 ( .A1(n469), .A2(G214), .ZN(n422) );
  XNOR2_X1 U541 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U542 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U543 ( .A(n445), .B(KEYINPUT10), .ZN(n474) );
  XNOR2_X1 U544 ( .A(n425), .B(n474), .ZN(n430) );
  XNOR2_X1 U545 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U546 ( .A(n452), .B(n428), .ZN(n429) );
  XNOR2_X1 U547 ( .A(n430), .B(n429), .ZN(n679) );
  NOR2_X1 U548 ( .A1(G902), .A2(n679), .ZN(n433) );
  XNOR2_X1 U549 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n431) );
  XOR2_X1 U550 ( .A(n453), .B(G122), .Z(n435) );
  XOR2_X1 U551 ( .A(n443), .B(G134), .Z(n434) );
  XNOR2_X1 U552 ( .A(n435), .B(n434), .ZN(n440) );
  XOR2_X1 U553 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n438) );
  INV_X1 U554 ( .A(G217), .ZN(n436) );
  NOR2_X1 U555 ( .A1(n479), .A2(n436), .ZN(n437) );
  XOR2_X1 U556 ( .A(n438), .B(n437), .Z(n439) );
  XNOR2_X1 U557 ( .A(n440), .B(n439), .ZN(n693) );
  NOR2_X1 U558 ( .A1(G902), .A2(n693), .ZN(n442) );
  INV_X1 U559 ( .A(G478), .ZN(n441) );
  XNOR2_X1 U560 ( .A(n442), .B(n441), .ZN(n528) );
  INV_X1 U561 ( .A(n528), .ZN(n551) );
  NAND2_X1 U562 ( .A1(n552), .A2(n551), .ZN(n740) );
  XNOR2_X1 U563 ( .A(n468), .B(n505), .ZN(n451) );
  XNOR2_X1 U564 ( .A(n445), .B(n444), .ZN(n449) );
  NAND2_X1 U565 ( .A1(n446), .A2(G224), .ZN(n447) );
  XNOR2_X1 U566 ( .A(n447), .B(KEYINPUT87), .ZN(n448) );
  XNOR2_X1 U567 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U568 ( .A(n453), .B(n452), .ZN(n458) );
  XNOR2_X1 U569 ( .A(n472), .B(n456), .ZN(n457) );
  XNOR2_X2 U570 ( .A(G902), .B(KEYINPUT15), .ZN(n638) );
  NAND2_X1 U571 ( .A1(n642), .A2(n638), .ZN(n462) );
  NAND2_X1 U572 ( .A1(n573), .A2(n460), .ZN(n464) );
  AND2_X1 U573 ( .A1(n464), .A2(G210), .ZN(n461) );
  XNOR2_X2 U574 ( .A(n462), .B(n461), .ZN(n533) );
  INV_X1 U575 ( .A(n533), .ZN(n463) );
  NAND2_X1 U576 ( .A1(n464), .A2(G214), .ZN(n736) );
  NAND2_X1 U577 ( .A1(n737), .A2(n736), .ZN(n741) );
  XNOR2_X1 U578 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n465) );
  NAND2_X1 U579 ( .A1(n469), .A2(G210), .ZN(n470) );
  INV_X1 U580 ( .A(G137), .ZN(n473) );
  XNOR2_X2 U581 ( .A(KEYINPUT69), .B(KEYINPUT89), .ZN(n475) );
  XNOR2_X1 U582 ( .A(n476), .B(n475), .ZN(n478) );
  XNOR2_X1 U583 ( .A(n478), .B(n477), .ZN(n481) );
  NAND2_X1 U584 ( .A1(n638), .A2(G234), .ZN(n482) );
  AND2_X1 U585 ( .A1(n486), .A2(G217), .ZN(n484) );
  XNOR2_X1 U586 ( .A(KEYINPUT77), .B(KEYINPUT25), .ZN(n483) );
  XNOR2_X1 U587 ( .A(n484), .B(n483), .ZN(n485) );
  INV_X1 U588 ( .A(n486), .ZN(n488) );
  XNOR2_X2 U589 ( .A(n489), .B(KEYINPUT21), .ZN(n726) );
  INV_X1 U590 ( .A(n726), .ZN(n495) );
  XNOR2_X1 U591 ( .A(KEYINPUT14), .B(n490), .ZN(n720) );
  NOR2_X1 U592 ( .A1(n446), .A2(G900), .ZN(n491) );
  NAND2_X1 U593 ( .A1(n491), .A2(G902), .ZN(n492) );
  NAND2_X1 U594 ( .A1(n446), .A2(G952), .ZN(n579) );
  NAND2_X1 U595 ( .A1(n492), .A2(n579), .ZN(n493) );
  NAND2_X1 U596 ( .A1(n720), .A2(n493), .ZN(n517) );
  INV_X1 U597 ( .A(n517), .ZN(n494) );
  AND2_X1 U598 ( .A1(n495), .A2(n494), .ZN(n496) );
  AND2_X1 U599 ( .A1(n602), .A2(n496), .ZN(n541) );
  NAND2_X1 U600 ( .A1(n515), .A2(n541), .ZN(n497) );
  XNOR2_X1 U601 ( .A(n497), .B(KEYINPUT28), .ZN(n510) );
  XNOR2_X1 U602 ( .A(n499), .B(n498), .ZN(n504) );
  INV_X1 U603 ( .A(n500), .ZN(n502) );
  NAND2_X1 U604 ( .A1(n446), .A2(G227), .ZN(n501) );
  XNOR2_X1 U605 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U606 ( .A(n504), .B(n503), .ZN(n506) );
  XNOR2_X1 U607 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U608 ( .A(n508), .B(n507), .ZN(n673) );
  OR2_X1 U609 ( .A1(n673), .A2(G902), .ZN(n509) );
  XNOR2_X1 U610 ( .A(n509), .B(G469), .ZN(n617) );
  INV_X1 U611 ( .A(n617), .ZN(n547) );
  NOR2_X2 U612 ( .A1(n602), .A2(n599), .ZN(n512) );
  INV_X1 U613 ( .A(KEYINPUT67), .ZN(n511) );
  NAND2_X1 U614 ( .A1(n586), .A2(n617), .ZN(n514) );
  INV_X1 U615 ( .A(KEYINPUT104), .ZN(n513) );
  NAND2_X1 U616 ( .A1(n515), .A2(n736), .ZN(n516) );
  XNOR2_X1 U617 ( .A(n516), .B(KEYINPUT30), .ZN(n518) );
  INV_X1 U618 ( .A(KEYINPUT76), .ZN(n521) );
  INV_X1 U619 ( .A(KEYINPUT40), .ZN(n524) );
  INV_X1 U620 ( .A(KEYINPUT64), .ZN(n525) );
  XNOR2_X1 U621 ( .A(n527), .B(n526), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n552), .A2(n528), .ZN(n530) );
  INV_X1 U623 ( .A(KEYINPUT98), .ZN(n529) );
  XNOR2_X1 U624 ( .A(n530), .B(n529), .ZN(n567) );
  INV_X1 U625 ( .A(n540), .ZN(n531) );
  OR2_X1 U626 ( .A1(n567), .A2(n531), .ZN(n532) );
  XNOR2_X1 U627 ( .A(n532), .B(KEYINPUT99), .ZN(n742) );
  INV_X1 U628 ( .A(KEYINPUT85), .ZN(n534) );
  OR2_X1 U629 ( .A1(n571), .A2(n536), .ZN(n704) );
  INV_X1 U630 ( .A(KEYINPUT47), .ZN(n537) );
  INV_X1 U631 ( .A(KEYINPUT102), .ZN(n539) );
  XNOR2_X1 U632 ( .A(n540), .B(n539), .ZN(n709) );
  INV_X1 U633 ( .A(n515), .ZN(n616) );
  NAND2_X1 U634 ( .A1(n362), .A2(n544), .ZN(n545) );
  XNOR2_X1 U635 ( .A(n545), .B(KEYINPUT36), .ZN(n548) );
  XNOR2_X1 U636 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n546) );
  XNOR2_X2 U637 ( .A(n547), .B(n546), .ZN(n721) );
  NAND2_X1 U638 ( .A1(n354), .A2(n533), .ZN(n550) );
  OR2_X1 U639 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U640 ( .A(n553), .B(KEYINPUT101), .ZN(n594) );
  NAND2_X1 U641 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X1 U642 ( .A(n557), .B(n556), .ZN(n564) );
  NAND2_X1 U643 ( .A1(n362), .A2(n736), .ZN(n559) );
  INV_X1 U644 ( .A(n587), .ZN(n558) );
  NOR2_X1 U645 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U646 ( .A1(n560), .A2(n721), .ZN(n562) );
  XNOR2_X1 U647 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n561) );
  XNOR2_X1 U648 ( .A(n562), .B(n561), .ZN(n563) );
  OR2_X1 U649 ( .A1(n563), .A2(n533), .ZN(n651) );
  NAND2_X1 U650 ( .A1(n564), .A2(n651), .ZN(n566) );
  INV_X1 U651 ( .A(KEYINPUT82), .ZN(n565) );
  XNOR2_X1 U652 ( .A(n566), .B(n565), .ZN(n636) );
  INV_X1 U653 ( .A(n567), .ZN(n703) );
  OR2_X1 U654 ( .A1(n568), .A2(n703), .ZN(n653) );
  AND2_X1 U655 ( .A1(n653), .A2(KEYINPUT2), .ZN(n569) );
  NAND2_X1 U656 ( .A1(n636), .A2(n569), .ZN(n570) );
  INV_X1 U657 ( .A(n571), .ZN(n584) );
  INV_X1 U658 ( .A(G898), .ZN(n572) );
  NAND2_X1 U659 ( .A1(n572), .A2(G953), .ZN(n577) );
  NOR2_X1 U660 ( .A1(n577), .A2(n573), .ZN(n574) );
  NAND2_X1 U661 ( .A1(n720), .A2(n574), .ZN(n576) );
  INV_X1 U662 ( .A(KEYINPUT88), .ZN(n575) );
  NAND2_X1 U663 ( .A1(n576), .A2(n575), .ZN(n583) );
  INV_X1 U664 ( .A(n577), .ZN(n763) );
  AND2_X1 U665 ( .A1(G902), .A2(KEYINPUT88), .ZN(n578) );
  NAND2_X1 U666 ( .A1(n763), .A2(n578), .ZN(n580) );
  NAND2_X1 U667 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U668 ( .A1(n720), .A2(n581), .ZN(n582) );
  INV_X1 U669 ( .A(n620), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n587), .A2(n722), .ZN(n588) );
  INV_X1 U671 ( .A(KEYINPUT33), .ZN(n589) );
  INV_X1 U672 ( .A(n752), .ZN(n591) );
  NAND2_X1 U673 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U674 ( .A(KEYINPUT35), .ZN(n595) );
  XNOR2_X2 U675 ( .A(n596), .B(n595), .ZN(n773) );
  INV_X1 U676 ( .A(KEYINPUT84), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n773), .A2(n597), .ZN(n598) );
  INV_X1 U678 ( .A(KEYINPUT44), .ZN(n630) );
  AND2_X1 U679 ( .A1(n598), .A2(n630), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n592), .A2(n363), .ZN(n601) );
  XNOR2_X1 U681 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n601), .B(n600), .ZN(n626) );
  INV_X1 U683 ( .A(n602), .ZN(n603) );
  INV_X1 U684 ( .A(KEYINPUT65), .ZN(n604) );
  NAND2_X1 U685 ( .A1(n721), .A2(n616), .ZN(n605) );
  NOR2_X1 U686 ( .A1(n606), .A2(n605), .ZN(n702) );
  INV_X1 U687 ( .A(n702), .ZN(n607) );
  AND2_X1 U688 ( .A1(n630), .A2(KEYINPUT84), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n773), .A2(n609), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n634) );
  NAND2_X1 U692 ( .A1(n722), .A2(n728), .ZN(n614) );
  OR2_X1 U693 ( .A1(n721), .A2(n614), .ZN(n732) );
  OR2_X1 U694 ( .A1(n620), .A2(n732), .ZN(n615) );
  XNOR2_X1 U695 ( .A(n615), .B(KEYINPUT31), .ZN(n712) );
  AND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n618), .A2(n722), .ZN(n619) );
  OR2_X1 U698 ( .A1(n712), .A2(n621), .ZN(n623) );
  INV_X1 U699 ( .A(n742), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n587), .A2(n602), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n624), .A2(n721), .ZN(n625) );
  OR2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n652) );
  NAND2_X1 U704 ( .A1(n627), .A2(n652), .ZN(n629) );
  INV_X1 U705 ( .A(KEYINPUT100), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n629), .B(n628), .ZN(n632) );
  OR2_X1 U707 ( .A1(n773), .A2(n630), .ZN(n631) );
  AND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n633) );
  AND2_X1 U709 ( .A1(n636), .A2(n653), .ZN(n657) );
  XOR2_X1 U710 ( .A(KEYINPUT80), .B(n638), .Z(n639) );
  XNOR2_X1 U711 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n640), .B(KEYINPUT118), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(n646) );
  INV_X1 U715 ( .A(G952), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n645), .A2(G953), .ZN(n682) );
  INV_X1 U717 ( .A(n682), .ZN(n696) );
  XNOR2_X1 U718 ( .A(n647), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U719 ( .A(n709), .ZN(n648) );
  NOR2_X1 U720 ( .A1(n704), .A2(n648), .ZN(n650) );
  XNOR2_X1 U721 ( .A(G146), .B(KEYINPUT109), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n650), .B(n649), .ZN(G48) );
  XNOR2_X1 U723 ( .A(n651), .B(G140), .ZN(G42) );
  XNOR2_X1 U724 ( .A(n652), .B(G101), .ZN(G3) );
  XNOR2_X1 U725 ( .A(n653), .B(G134), .ZN(G36) );
  XOR2_X1 U726 ( .A(n655), .B(n654), .Z(n659) );
  XNOR2_X1 U727 ( .A(n659), .B(KEYINPUT126), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n658), .A2(n446), .ZN(n663) );
  XOR2_X1 U730 ( .A(G227), .B(n659), .Z(n660) );
  NAND2_X1 U731 ( .A1(n660), .A2(G900), .ZN(n661) );
  NAND2_X1 U732 ( .A1(n661), .A2(G953), .ZN(n662) );
  NAND2_X1 U733 ( .A1(n663), .A2(n662), .ZN(G72) );
  XNOR2_X1 U734 ( .A(n664), .B(G119), .ZN(G21) );
  NAND2_X1 U735 ( .A1(n687), .A2(G472), .ZN(n668) );
  XNOR2_X1 U736 ( .A(KEYINPUT107), .B(KEYINPUT62), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n355), .B(n665), .ZN(n667) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n669), .A2(n682), .ZN(n671) );
  XNOR2_X1 U740 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(G57) );
  NAND2_X1 U742 ( .A1(n687), .A2(G469), .ZN(n675) );
  XNOR2_X1 U743 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U745 ( .A1(n676), .A2(n682), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(KEYINPUT119), .ZN(G54) );
  NAND2_X1 U747 ( .A1(n687), .A2(G475), .ZN(n681) );
  XNOR2_X1 U748 ( .A(KEYINPUT120), .B(KEYINPUT59), .ZN(n678) );
  XNOR2_X1 U749 ( .A(n681), .B(n680), .ZN(n683) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n685) );
  XNOR2_X1 U751 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n685), .B(n684), .ZN(G60) );
  XOR2_X1 U753 ( .A(n368), .B(G131), .Z(G33) );
  NAND2_X1 U754 ( .A1(n369), .A2(G217), .ZN(n691) );
  XNOR2_X1 U755 ( .A(n689), .B(KEYINPUT123), .ZN(n690) );
  XNOR2_X1 U756 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U757 ( .A1(n692), .A2(n696), .ZN(G66) );
  NAND2_X1 U758 ( .A1(n369), .A2(G478), .ZN(n695) );
  XNOR2_X1 U759 ( .A(n693), .B(KEYINPUT122), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n695), .B(n694), .ZN(n697) );
  NOR2_X1 U761 ( .A1(n697), .A2(n696), .ZN(G63) );
  NAND2_X1 U762 ( .A1(n621), .A2(n709), .ZN(n698) );
  XNOR2_X1 U763 ( .A(n698), .B(G104), .ZN(G6) );
  XOR2_X1 U764 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n700) );
  NAND2_X1 U765 ( .A1(n621), .A2(n567), .ZN(n699) );
  XNOR2_X1 U766 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U767 ( .A(G107), .B(n701), .ZN(G9) );
  XOR2_X1 U768 ( .A(n702), .B(G110), .Z(G12) );
  NOR2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n706) );
  XNOR2_X1 U770 ( .A(KEYINPUT108), .B(KEYINPUT29), .ZN(n705) );
  XNOR2_X1 U771 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U772 ( .A(G128), .B(n707), .ZN(G30) );
  XOR2_X1 U773 ( .A(G143), .B(n708), .Z(G45) );
  NAND2_X1 U774 ( .A1(n709), .A2(n712), .ZN(n710) );
  XNOR2_X1 U775 ( .A(n710), .B(KEYINPUT110), .ZN(n711) );
  XNOR2_X1 U776 ( .A(G113), .B(n711), .ZN(G15) );
  XOR2_X1 U777 ( .A(G116), .B(KEYINPUT111), .Z(n714) );
  NAND2_X1 U778 ( .A1(n712), .A2(n567), .ZN(n713) );
  XNOR2_X1 U779 ( .A(n714), .B(n713), .ZN(G18) );
  XOR2_X1 U780 ( .A(KEYINPUT37), .B(KEYINPUT112), .Z(n715) );
  XNOR2_X1 U781 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U782 ( .A(G125), .B(n717), .ZN(G27) );
  XNOR2_X1 U783 ( .A(KEYINPUT79), .B(KEYINPUT2), .ZN(n718) );
  NAND2_X1 U784 ( .A1(G952), .A2(n720), .ZN(n751) );
  XOR2_X1 U785 ( .A(KEYINPUT113), .B(KEYINPUT50), .Z(n725) );
  INV_X1 U786 ( .A(n721), .ZN(n723) );
  NOR2_X1 U787 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U788 ( .A(n725), .B(n724), .Z(n731) );
  NAND2_X1 U789 ( .A1(n356), .A2(n726), .ZN(n727) );
  XNOR2_X1 U790 ( .A(n727), .B(KEYINPUT49), .ZN(n729) );
  NOR2_X1 U791 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U792 ( .A1(n731), .A2(n730), .ZN(n733) );
  AND2_X1 U793 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U794 ( .A(KEYINPUT51), .B(n734), .Z(n735) );
  NOR2_X1 U795 ( .A1(n753), .A2(n735), .ZN(n748) );
  NOR2_X1 U796 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U797 ( .A(n738), .B(KEYINPUT114), .ZN(n739) );
  NOR2_X1 U798 ( .A1(n740), .A2(n739), .ZN(n745) );
  NOR2_X1 U799 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U800 ( .A(KEYINPUT115), .B(n743), .Z(n744) );
  NOR2_X1 U801 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U802 ( .A1(n746), .A2(n752), .ZN(n747) );
  NOR2_X1 U803 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U804 ( .A(n749), .B(KEYINPUT52), .ZN(n750) );
  NOR2_X1 U805 ( .A1(n751), .A2(n750), .ZN(n755) );
  NOR2_X1 U806 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U807 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U808 ( .A(n756), .B(KEYINPUT116), .ZN(n757) );
  AND2_X1 U809 ( .A1(n758), .A2(n757), .ZN(n760) );
  XNOR2_X1 U810 ( .A(n762), .B(n761), .ZN(n764) );
  NOR2_X1 U811 ( .A1(n764), .A2(n763), .ZN(n771) );
  XNOR2_X1 U812 ( .A(n765), .B(KEYINPUT124), .ZN(n769) );
  NAND2_X1 U813 ( .A1(G953), .A2(G224), .ZN(n766) );
  XNOR2_X1 U814 ( .A(KEYINPUT61), .B(n766), .ZN(n767) );
  NAND2_X1 U815 ( .A1(n767), .A2(G898), .ZN(n768) );
  NAND2_X1 U816 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U817 ( .A(n771), .B(n770), .ZN(n772) );
  XOR2_X1 U818 ( .A(KEYINPUT125), .B(n772), .Z(G69) );
  XNOR2_X1 U819 ( .A(n773), .B(G122), .ZN(G24) );
  XOR2_X1 U820 ( .A(n774), .B(G137), .Z(G39) );
endmodule

