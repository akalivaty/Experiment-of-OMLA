//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT66), .B(G77), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G58), .A2(G232), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT67), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT68), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n207), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n227), .B(new_n230), .C1(new_n218), .C2(new_n219), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n221), .A2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  INV_X1    g0042(.A(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT70), .B(G50), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  AND2_X1   g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(G274), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G222), .A2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G223), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n253), .B1(new_n209), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n262), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G169), .ZN(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(new_n274), .ZN(new_n277));
  INV_X1    g0077(.A(G13), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n278), .A2(new_n225), .A3(G1), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n224), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n258), .A2(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G50), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G50), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n282), .A2(new_n285), .B1(new_n286), .B2(new_n279), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n225), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n225), .A2(new_n268), .A3(KEYINPUT71), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT71), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(G20), .B2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n289), .A2(new_n291), .B1(new_n295), .B2(G150), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n203), .A2(G20), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n281), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n287), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n277), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n300), .B(KEYINPUT9), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT72), .B1(new_n274), .B2(G190), .ZN(new_n304));
  INV_X1    g0104(.A(G200), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n303), .B(new_n304), .C1(new_n305), .C2(new_n274), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT18), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT16), .ZN(new_n311));
  INV_X1    g0111(.A(G68), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT7), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(G20), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT75), .B1(new_n268), .B2(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n269), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n271), .A2(KEYINPUT75), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n313), .B1(new_n263), .B2(G20), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n312), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n295), .A2(G159), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n243), .A2(new_n312), .ZN(new_n322));
  OAI21_X1  g0122(.A(G20), .B1(new_n322), .B2(new_n202), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n311), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n263), .A2(new_n313), .A3(G20), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT7), .B1(new_n272), .B2(new_n225), .ZN(new_n327));
  OAI21_X1  g0127(.A(G68), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n324), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT16), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n325), .A2(new_n281), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n288), .B1(new_n258), .B2(G20), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(new_n282), .B1(new_n279), .B2(new_n288), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  OR2_X1    g0135(.A1(G223), .A2(G1698), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n261), .A2(G1698), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n269), .A2(new_n336), .A3(new_n271), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G87), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n253), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n253), .A2(G232), .A3(new_n259), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n257), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n335), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n253), .B1(new_n338), .B2(new_n339), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n257), .A2(new_n343), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n346), .A2(new_n347), .A3(new_n276), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n310), .B1(new_n334), .B2(new_n350), .ZN(new_n351));
  AOI211_X1 g0151(.A(KEYINPUT18), .B(new_n349), .C1(new_n331), .C2(new_n333), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT76), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n333), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n312), .B1(new_n319), .B2(new_n355), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n356), .A2(new_n324), .A3(new_n311), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n299), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n354), .B1(new_n358), .B2(new_n325), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT18), .B1(new_n359), .B2(new_n349), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT76), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n334), .A2(new_n310), .A3(new_n350), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n353), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n342), .A2(new_n344), .ZN(new_n365));
  INV_X1    g0165(.A(G190), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n365), .B2(G200), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n359), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT17), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n286), .B1(new_n292), .B2(new_n294), .ZN(new_n372));
  INV_X1    g0172(.A(G77), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n290), .A2(new_n373), .B1(new_n225), .B2(G68), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n281), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT11), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(KEYINPUT11), .B(new_n281), .C1(new_n372), .C2(new_n374), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT73), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT73), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n377), .A2(new_n381), .A3(new_n378), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n278), .A2(G1), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n225), .A2(G68), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT12), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n383), .B(new_n384), .C1(KEYINPUT74), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n386), .B(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n282), .A2(G68), .A3(new_n283), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n380), .A2(new_n382), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT14), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT13), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n261), .A2(new_n265), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n265), .A2(G232), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n263), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n341), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n256), .B1(new_n251), .B2(new_n252), .ZN(new_n399));
  INV_X1    g0199(.A(G274), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n251), .B2(new_n252), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n399), .A2(G238), .B1(new_n401), .B2(new_n256), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n392), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n253), .B1(new_n395), .B2(new_n396), .ZN(new_n404));
  INV_X1    g0204(.A(G238), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n257), .B1(new_n260), .B2(new_n405), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n404), .A2(new_n406), .A3(KEYINPUT13), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n391), .B(G169), .C1(new_n403), .C2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n398), .A2(new_n392), .A3(new_n402), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT13), .B1(new_n404), .B2(new_n406), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(G179), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n410), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n391), .B1(new_n413), .B2(G169), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n390), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(G200), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n388), .A2(new_n389), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n379), .B2(KEYINPUT73), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n409), .A2(G190), .A3(new_n410), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n416), .A2(new_n418), .A3(new_n382), .A4(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n257), .B1(new_n260), .B2(new_n210), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n263), .A2(G238), .A3(G1698), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n263), .A2(G232), .A3(new_n265), .ZN(new_n423));
  INV_X1    g0223(.A(G107), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n422), .B(new_n423), .C1(new_n424), .C2(new_n263), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n421), .B1(new_n425), .B2(new_n341), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n291), .B1(new_n208), .B2(G20), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n289), .A2(new_n295), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n299), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n282), .A2(G77), .A3(new_n283), .ZN(new_n432));
  INV_X1    g0232(.A(new_n279), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n208), .B2(new_n433), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n426), .A2(G169), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n426), .A2(new_n276), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n426), .A2(G190), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n431), .A2(new_n434), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(new_n305), .C2(new_n426), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n415), .A2(new_n420), .A3(new_n438), .A4(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n309), .A2(new_n371), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT19), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n225), .B1(new_n396), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G87), .ZN(new_n446));
  INV_X1    g0246(.A(G97), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n424), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n269), .A2(new_n271), .A3(new_n225), .A4(G68), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n444), .B1(new_n290), .B2(new_n447), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(new_n281), .B1(new_n279), .B2(new_n427), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT83), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT78), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n258), .B2(G33), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n268), .A2(KEYINPUT78), .A3(G1), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n282), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n454), .B1(new_n459), .B2(new_n427), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n282), .A2(new_n458), .A3(KEYINPUT83), .A4(new_n428), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n453), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n258), .A2(G45), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n401), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n253), .A2(G250), .A3(new_n463), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n269), .A2(new_n271), .A3(G238), .A4(new_n265), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n269), .A2(new_n271), .A3(G244), .A4(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G116), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n467), .B1(new_n341), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n276), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n341), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n463), .A2(G250), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n253), .A2(new_n475), .B1(new_n401), .B2(new_n464), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n335), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n462), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n282), .A2(new_n458), .A3(G87), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n453), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n474), .A2(G190), .A3(new_n476), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n472), .B2(new_n305), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n269), .A2(new_n271), .A3(G244), .A4(new_n265), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT79), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n263), .A2(KEYINPUT79), .A3(G244), .A4(new_n265), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(KEYINPUT4), .A2(G244), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n269), .A2(new_n271), .A3(new_n492), .A4(new_n265), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT80), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n263), .A2(KEYINPUT80), .A3(new_n265), .A4(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n269), .A2(new_n271), .A3(G250), .A4(G1698), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n491), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n341), .ZN(new_n503));
  OR2_X1    g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  NAND2_X1  g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n463), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n401), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT5), .B(G41), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n464), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n253), .ZN(new_n510));
  INV_X1    g0310(.A(G257), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n503), .A2(KEYINPUT81), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT81), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n500), .B1(new_n495), .B2(new_n496), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n253), .B1(new_n516), .B2(new_n491), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n517), .B2(new_n512), .ZN(new_n518));
  AOI21_X1  g0318(.A(G169), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n295), .A2(G77), .ZN(new_n520));
  XNOR2_X1  g0320(.A(G97), .B(G107), .ZN(new_n521));
  NOR2_X1   g0321(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n522), .B1(KEYINPUT6), .B2(new_n447), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n520), .B1(new_n526), .B2(new_n225), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n424), .B1(new_n318), .B2(new_n319), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n281), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n433), .A2(G97), .ZN(new_n530));
  INV_X1    g0330(.A(new_n459), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(G97), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n503), .A2(new_n513), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(G179), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT82), .B1(new_n519), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT81), .B1(new_n503), .B2(new_n513), .ZN(new_n537));
  AOI211_X1 g0337(.A(new_n515), .B(new_n512), .C1(new_n502), .C2(new_n341), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n335), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT82), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n517), .A2(new_n512), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(new_n276), .B1(new_n529), .B2(new_n532), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n533), .B1(G200), .B2(new_n534), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n514), .A2(new_n518), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n366), .B2(new_n545), .ZN(new_n546));
  AND4_X1   g0346(.A1(new_n485), .A2(new_n536), .A3(new_n543), .A4(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n506), .A2(new_n341), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(G270), .B1(new_n401), .B2(new_n506), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n269), .A2(new_n271), .A3(G264), .A4(G1698), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n269), .A2(new_n271), .A3(G257), .A4(new_n265), .ZN(new_n551));
  INV_X1    g0351(.A(G303), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n550), .B(new_n551), .C1(new_n552), .C2(new_n263), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n341), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n335), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n282), .A2(new_n458), .A3(G116), .ZN(new_n556));
  INV_X1    g0356(.A(G116), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n279), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n280), .A2(new_n224), .B1(G20), .B2(new_n557), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n499), .B(new_n225), .C1(G33), .C2(new_n447), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n559), .A2(KEYINPUT20), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT20), .B1(new_n559), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n556), .B(new_n558), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n555), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n549), .A2(new_n554), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n567), .B2(G200), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n549), .A2(new_n554), .A3(G190), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n563), .A2(G179), .A3(new_n554), .A4(new_n549), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n567), .A2(new_n563), .A3(KEYINPUT21), .A4(G169), .ZN(new_n572));
  AND4_X1   g0372(.A1(new_n566), .A2(new_n570), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n531), .A2(G107), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n279), .A2(new_n424), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT25), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n269), .A2(new_n271), .A3(new_n225), .A4(G87), .ZN(new_n580));
  XNOR2_X1  g0380(.A(KEYINPUT84), .B(KEYINPUT22), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT22), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(KEYINPUT84), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n263), .A2(new_n225), .A3(G87), .A4(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n470), .A2(G20), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT23), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n225), .B2(G107), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n424), .A2(KEYINPUT23), .A3(G20), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n582), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n591), .B(KEYINPUT24), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n579), .B1(new_n592), .B2(new_n281), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n269), .A2(new_n271), .A3(G250), .A4(new_n265), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT85), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT85), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n263), .A2(new_n597), .A3(G250), .A4(new_n265), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G294), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n263), .A2(G257), .A3(G1698), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n596), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n341), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n548), .A2(G264), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n507), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT86), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(G169), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n601), .A2(new_n341), .B1(G264), .B2(new_n548), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(G179), .A3(new_n507), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n605), .B1(new_n604), .B2(G169), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n594), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n604), .A2(G200), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n607), .A2(G190), .A3(new_n507), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n593), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n574), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n443), .A2(new_n547), .A3(new_n616), .ZN(G372));
  NOR2_X1   g0417(.A1(new_n351), .A2(new_n352), .ZN(new_n618));
  INV_X1    g0418(.A(new_n415), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n420), .B2(new_n437), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT17), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n369), .B(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n618), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT90), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n307), .A2(new_n308), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n623), .B2(KEYINPUT90), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n301), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT87), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n453), .B2(new_n480), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n453), .A2(new_n628), .A3(new_n480), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n483), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n462), .A2(new_n473), .A3(new_n478), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT88), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n477), .A2(G200), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n453), .A2(new_n628), .A3(new_n480), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n635), .B(new_n482), .C1(new_n636), .C2(new_n629), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT88), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n479), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n615), .B1(new_n634), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT89), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n572), .A2(new_n571), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT21), .B1(new_n555), .B2(new_n563), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n566), .A2(KEYINPUT89), .A3(new_n571), .A4(new_n572), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n640), .B1(new_n646), .B2(new_n612), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n536), .A2(new_n543), .A3(new_n546), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n479), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n634), .A2(new_n639), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n519), .A2(new_n535), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT26), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n484), .B1(new_n536), .B2(new_n543), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(KEYINPUT26), .B2(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n443), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n627), .A2(new_n656), .ZN(G369));
  NAND2_X1  g0457(.A1(new_n383), .A2(new_n225), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n563), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n646), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n574), .A2(KEYINPUT91), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(new_n664), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n574), .A2(KEYINPUT91), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n593), .A2(new_n613), .A3(new_n614), .ZN(new_n672));
  INV_X1    g0472(.A(new_n663), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n611), .B(new_n672), .C1(new_n593), .C2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n611), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n566), .A2(new_n571), .A3(new_n572), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n673), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT92), .Z(new_n679));
  XOR2_X1   g0479(.A(new_n663), .B(KEYINPUT93), .Z(new_n680));
  AOI22_X1  g0480(.A1(new_n679), .A2(new_n675), .B1(new_n612), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n676), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n228), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n448), .A2(G116), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G1), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n222), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n650), .A2(KEYINPUT26), .A3(new_n651), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n653), .B2(KEYINPUT26), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n640), .B1(new_n612), .B2(new_n677), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n479), .B1(new_n693), .B2(new_n648), .ZN(new_n694));
  OAI211_X1 g0494(.A(KEYINPUT29), .B(new_n673), .C1(new_n692), .C2(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n655), .A2(new_n680), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(KEYINPUT29), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n537), .A2(new_n538), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n602), .A2(new_n603), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n549), .A2(new_n554), .A3(G179), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n701), .A2(new_n702), .A3(new_n477), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT30), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n472), .A2(G179), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n534), .A2(new_n604), .A3(new_n567), .A4(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n702), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(KEYINPUT30), .A3(new_n472), .A4(new_n607), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n706), .B1(new_n545), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n699), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n703), .A2(new_n518), .A3(new_n514), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n703), .A2(KEYINPUT30), .A3(new_n518), .A4(new_n514), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n713), .A2(KEYINPUT94), .A3(new_n714), .A4(new_n706), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n710), .A2(new_n663), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  AND4_X1   g0517(.A1(new_n611), .A2(new_n573), .A3(new_n672), .A4(new_n680), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n716), .A2(new_n717), .B1(new_n547), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n680), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT31), .B(new_n720), .C1(new_n704), .C2(new_n709), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n698), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n697), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n689), .B1(new_n725), .B2(G1), .ZN(G364));
  NOR2_X1   g0526(.A1(new_n669), .A2(G330), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n278), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n258), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n684), .A2(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n671), .A2(new_n727), .A3(new_n731), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT95), .Z(new_n733));
  INV_X1    g0533(.A(new_n731), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n224), .B1(G20), .B2(new_n335), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n225), .A2(new_n276), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n366), .A3(new_n305), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n225), .A2(G190), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G179), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n739), .A2(G311), .B1(new_n743), .B2(G329), .ZN(new_n744));
  INV_X1    g0544(.A(G322), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n225), .A2(new_n366), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(G179), .A3(new_n305), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n744), .B(new_n272), .C1(new_n745), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n737), .A2(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n366), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G326), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n225), .B1(new_n741), .B2(G190), .ZN(new_n753));
  INV_X1    g0553(.A(G294), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n751), .A2(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n748), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n749), .A2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT33), .B(G317), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(new_n759), .B2(KEYINPUT99), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(KEYINPUT99), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n305), .A2(G179), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT97), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n746), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n760), .A2(new_n761), .B1(new_n765), .B2(G303), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n763), .A2(new_n740), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT98), .Z(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n756), .B(new_n766), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n768), .A2(G107), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n753), .A2(new_n447), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n263), .B1(new_n747), .B2(new_n243), .C1(new_n209), .C2(new_n738), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n773), .B(new_n774), .C1(G68), .C2(new_n757), .ZN(new_n775));
  INV_X1    g0575(.A(G159), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n742), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n777), .B(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G50), .B2(new_n750), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n765), .A2(G87), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n772), .A2(new_n775), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n736), .B1(new_n771), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n735), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n683), .A2(new_n272), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G355), .A2(new_n788), .B1(new_n557), .B2(new_n683), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n246), .A2(G45), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n683), .A2(new_n263), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(G45), .B2(new_n222), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n789), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n734), .B(new_n783), .C1(new_n787), .C2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n786), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n669), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n733), .A2(new_n796), .ZN(G396));
  NAND2_X1  g0597(.A1(new_n655), .A2(new_n680), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n441), .B1(new_n440), .B2(new_n673), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n438), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n438), .A2(new_n663), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT101), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n680), .B(new_n803), .C1(new_n649), .C2(new_n654), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n798), .A2(KEYINPUT101), .A3(new_n804), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n722), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT102), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n812), .B(new_n734), .C1(new_n722), .C2(new_n810), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n735), .A2(new_n784), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n263), .B1(new_n753), .B2(new_n243), .C1(new_n816), .C2(new_n742), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n769), .A2(new_n312), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(G50), .C2(new_n765), .ZN(new_n819));
  INV_X1    g0619(.A(new_n747), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G143), .A2(new_n820), .B1(new_n739), .B2(G159), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  INV_X1    g0622(.A(G150), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n821), .B1(new_n822), .B2(new_n751), .C1(new_n823), .C2(new_n758), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n768), .A2(G87), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n773), .B1(new_n750), .B2(G303), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n770), .B2(new_n758), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n263), .B1(new_n743), .B2(G311), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n829), .B1(new_n557), .B2(new_n738), .C1(new_n754), .C2(new_n747), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n828), .B(new_n830), .C1(G107), .C2(new_n765), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n819), .A2(new_n825), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n731), .B1(G77), .B2(new_n815), .C1(new_n832), .C2(new_n736), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n784), .B2(new_n804), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT100), .Z(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n813), .A2(new_n836), .ZN(G384));
  NOR2_X1   g0637(.A1(new_n728), .A2(new_n258), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT107), .ZN(new_n839));
  INV_X1    g0639(.A(new_n661), .ZN(new_n840));
  INV_X1    g0640(.A(new_n618), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n334), .B(new_n840), .C1(new_n622), .C2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n334), .A2(new_n840), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(KEYINPUT106), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n334), .A2(new_n350), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n369), .A2(new_n846), .A3(new_n844), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n845), .B(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT38), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n311), .B1(new_n356), .B2(new_n324), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n850), .A2(KEYINPUT104), .A3(new_n281), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT104), .B1(new_n850), .B2(new_n281), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n851), .A2(new_n852), .A3(new_n357), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT105), .B1(new_n853), .B2(new_n354), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT104), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT16), .B1(new_n328), .B2(new_n329), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(new_n299), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n850), .A2(KEYINPUT104), .A3(new_n281), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n330), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT105), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n859), .A2(new_n860), .A3(new_n333), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n854), .A2(new_n840), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n364), .B2(new_n370), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n854), .A2(new_n350), .A3(new_n861), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n864), .A3(new_n369), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n369), .A2(new_n846), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(new_n843), .A3(new_n844), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n863), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n849), .B1(new_n869), .B2(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n716), .A2(new_n717), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n547), .A2(new_n718), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n710), .A2(new_n715), .A3(KEYINPUT31), .A4(new_n663), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n415), .A2(KEYINPUT103), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT103), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n876), .B(new_n390), .C1(new_n412), .C2(new_n414), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n390), .A2(new_n663), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n420), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n390), .B(new_n663), .C1(new_n412), .C2(new_n414), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n803), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n874), .A2(KEYINPUT40), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n839), .B1(new_n870), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n863), .ZN(new_n887));
  INV_X1    g0687(.A(new_n369), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n850), .A2(new_n281), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n357), .B1(new_n889), .B2(new_n855), .ZN(new_n890));
  AOI211_X1 g0690(.A(KEYINPUT105), .B(new_n354), .C1(new_n890), .C2(new_n858), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n860), .B1(new_n859), .B2(new_n333), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n888), .B1(new_n893), .B2(new_n350), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n843), .B1(new_n894), .B2(new_n862), .ZN(new_n895));
  INV_X1    g0695(.A(new_n868), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n887), .B(KEYINPUT38), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n849), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n900), .B(new_n883), .C1(new_n719), .C2(new_n873), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(new_n901), .A3(KEYINPUT107), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n886), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n883), .B1(new_n719), .B2(new_n873), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n866), .A2(new_n868), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT38), .B1(new_n905), .B2(new_n887), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n896), .B1(new_n865), .B2(KEYINPUT37), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n907), .A2(new_n908), .A3(new_n863), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n904), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n903), .B1(new_n900), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n443), .A2(new_n874), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n698), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n443), .B(new_n695), .C1(new_n696), .C2(KEYINPUT29), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n627), .ZN(new_n916));
  INV_X1    g0716(.A(new_n882), .ZN(new_n917));
  INV_X1    g0717(.A(new_n802), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n807), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n908), .B1(new_n907), .B2(new_n863), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n897), .A2(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n919), .A2(new_n921), .B1(new_n841), .B2(new_n661), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n909), .B2(new_n849), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n875), .A2(new_n877), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n673), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n897), .A2(new_n920), .A3(KEYINPUT39), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n916), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n838), .B1(new_n914), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n914), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT35), .ZN(new_n934));
  OAI211_X1 g0734(.A(G116), .B(new_n226), .C1(new_n526), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n934), .B2(new_n526), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT36), .Z(new_n937));
  NOR3_X1   g0737(.A1(new_n209), .A2(new_n222), .A3(new_n322), .ZN(new_n938));
  INV_X1    g0738(.A(new_n201), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n312), .ZN(new_n940));
  OAI211_X1 g0740(.A(G1), .B(new_n278), .C1(new_n938), .C2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n933), .A2(new_n937), .A3(new_n941), .ZN(G367));
  INV_X1    g0742(.A(new_n648), .ZN(new_n943));
  INV_X1    g0743(.A(new_n533), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n680), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n651), .A2(new_n720), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n681), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n681), .A2(new_n947), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT45), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n949), .A2(new_n676), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n676), .B1(new_n949), .B2(new_n952), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n679), .A2(new_n675), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n679), .A2(new_n675), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n671), .A2(KEYINPUT112), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT112), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n670), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n959), .B2(new_n962), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n724), .B1(new_n955), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n684), .B(KEYINPUT41), .Z(new_n966));
  OAI21_X1  g0766(.A(new_n729), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n636), .A2(new_n629), .A3(new_n673), .ZN(new_n968));
  MUX2_X1   g0768(.A(new_n650), .B(new_n633), .S(new_n968), .Z(new_n969));
  XNOR2_X1  g0769(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(KEYINPUT43), .B2(new_n969), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT109), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n947), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT109), .B1(new_n945), .B2(new_n946), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n612), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n536), .A2(new_n543), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n720), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n957), .A2(KEYINPUT42), .A3(new_n947), .ZN(new_n980));
  AOI21_X1  g0780(.A(KEYINPUT42), .B1(new_n957), .B2(new_n947), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n972), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT111), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n982), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n947), .B(new_n973), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n977), .B1(new_n987), .B2(new_n612), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n986), .B(new_n971), .C1(new_n988), .C2(new_n720), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT110), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n979), .A2(new_n982), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT110), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(new_n992), .A3(new_n971), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n987), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n985), .A2(new_n994), .B1(new_n676), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n983), .B(KEYINPUT111), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n995), .A2(new_n676), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n997), .A2(new_n998), .A3(new_n990), .A4(new_n993), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n967), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n240), .A2(new_n791), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1001), .B(new_n787), .C1(new_n228), .C2(new_n427), .ZN(new_n1002));
  INV_X1    g0802(.A(G311), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n758), .A2(new_n754), .B1(new_n751), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n753), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1004), .B1(G107), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n272), .B1(new_n747), .B2(new_n552), .ZN(new_n1007));
  INV_X1    g0807(.A(G317), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n738), .A2(new_n770), .B1(new_n742), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n767), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1007), .B(new_n1009), .C1(new_n1010), .C2(G97), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n765), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT46), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n764), .B2(new_n557), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1006), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1005), .A2(G68), .ZN(new_n1016));
  INV_X1    g0816(.A(G143), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n823), .B2(new_n747), .C1(new_n751), .C2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT113), .Z(new_n1019));
  AOI22_X1  g0819(.A1(G159), .A2(new_n757), .B1(new_n739), .B2(new_n939), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT114), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n263), .B1(new_n742), .B2(new_n822), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n1010), .B2(new_n208), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(new_n243), .C2(new_n764), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1015), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT47), .Z(new_n1026));
  OAI211_X1 g0826(.A(new_n731), .B(new_n1002), .C1(new_n1026), .C2(new_n736), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT115), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n969), .B2(new_n795), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1000), .A2(new_n1029), .ZN(G387));
  NAND2_X1  g0830(.A1(new_n964), .A2(new_n730), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n686), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n788), .A2(new_n1032), .B1(new_n424), .B2(new_n683), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT116), .ZN(new_n1034));
  AOI211_X1 g0834(.A(G45), .B(new_n1032), .C1(G68), .C2(G77), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n288), .A2(G50), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n683), .B(new_n263), .C1(new_n1035), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n237), .A2(G45), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1034), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n787), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n731), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1005), .A2(new_n428), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n751), .B2(new_n776), .C1(new_n288), .C2(new_n758), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n764), .A2(new_n209), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n820), .A2(G50), .B1(new_n743), .B2(G150), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1047), .B(new_n263), .C1(new_n312), .C2(new_n738), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n769), .B2(new_n447), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n764), .A2(new_n754), .B1(new_n770), .B2(new_n753), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G303), .A2(new_n739), .B1(new_n820), .B2(G317), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n1003), .B2(new_n758), .C1(new_n745), .C2(new_n751), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT48), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n1054), .B2(new_n1053), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT49), .Z(new_n1057));
  OAI221_X1 g0857(.A(new_n272), .B1(new_n752), .B2(new_n742), .C1(new_n767), .C2(new_n557), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1050), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1043), .B1(new_n1059), .B2(new_n735), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n675), .B2(new_n795), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n964), .A2(new_n725), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n684), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n964), .A2(new_n725), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1031), .B(new_n1061), .C1(new_n1063), .C2(new_n1064), .ZN(G393));
  OAI21_X1  g0865(.A(new_n1062), .B1(new_n953), .B2(new_n954), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n955), .A2(new_n725), .A3(new_n964), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n1067), .A3(new_n684), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n955), .A2(new_n730), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1042), .B1(G97), .B2(new_n683), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n249), .A2(new_n791), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n734), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n263), .B1(new_n742), .B2(new_n1017), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n758), .A2(new_n201), .B1(new_n753), .B2(new_n373), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(new_n289), .C2(new_n739), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n765), .A2(G68), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n751), .A2(new_n823), .B1(new_n776), .B2(new_n747), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT51), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1075), .A2(new_n826), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n272), .B1(new_n742), .B2(new_n745), .C1(new_n738), .C2(new_n754), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n758), .A2(new_n552), .B1(new_n753), .B2(new_n557), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(G283), .C2(new_n765), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n751), .A2(new_n1008), .B1(new_n1003), .B2(new_n747), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n772), .A3(new_n1084), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1079), .A2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1072), .B1(new_n736), .B2(new_n1086), .C1(new_n987), .C2(new_n795), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1069), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1068), .A2(new_n1088), .ZN(G390));
  AOI21_X1  g0889(.A(new_n698), .B1(new_n719), .B2(new_n873), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n443), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n915), .A2(new_n627), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n807), .A2(new_n918), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n882), .B1(new_n722), .B2(new_n803), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT119), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1090), .A2(new_n884), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1093), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n871), .A2(new_n872), .A3(new_n721), .ZN(new_n1100));
  AND4_X1   g0900(.A1(G330), .A2(new_n1100), .A3(new_n803), .A4(new_n882), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT88), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n638), .B1(new_n637), .B2(new_n479), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n672), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n610), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n608), .A3(new_n606), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n677), .B1(new_n1106), .B2(new_n594), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n633), .B1(new_n1108), .B2(new_n943), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n663), .B(new_n801), .C1(new_n1109), .C2(new_n691), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1101), .A2(new_n802), .A3(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1090), .A2(new_n803), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n882), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1092), .B1(new_n1099), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1093), .A2(new_n882), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1116), .A2(new_n926), .B1(new_n924), .B2(new_n928), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n899), .A2(new_n926), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n673), .B(new_n800), .C1(new_n692), .C2(new_n694), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n917), .B1(new_n1119), .B2(new_n918), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n884), .B(new_n1090), .C1(new_n1117), .C2(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n897), .A2(new_n920), .A3(KEYINPUT39), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT39), .B1(new_n897), .B2(new_n898), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1123), .A2(new_n1124), .B1(new_n919), .B2(new_n927), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n882), .B1(new_n1110), .B2(new_n802), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n927), .B1(new_n897), .B2(new_n898), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1101), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1125), .A2(new_n1128), .A3(KEYINPUT118), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT118), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1122), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n685), .B1(new_n1115), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1131), .B2(new_n1115), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n731), .B1(new_n289), .B2(new_n815), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n785), .B1(new_n924), .B2(new_n928), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n272), .B1(new_n742), .B2(new_n754), .C1(new_n747), .C2(new_n557), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n751), .A2(new_n770), .B1(new_n753), .B2(new_n373), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1136), .B(new_n1137), .C1(G87), .C2(new_n765), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n758), .A2(new_n424), .B1(new_n738), .B2(new_n447), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT120), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1138), .B(new_n1140), .C1(new_n312), .C2(new_n769), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1141), .A2(KEYINPUT121), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n764), .A2(new_n823), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT53), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n272), .B1(new_n743), .B2(G125), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT54), .B(G143), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1145), .B1(new_n816), .B2(new_n747), .C1(new_n738), .C2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n939), .B2(new_n1010), .ZN(new_n1148));
  INV_X1    g0948(.A(G128), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n751), .A2(new_n1149), .B1(new_n753), .B2(new_n776), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G137), .B2(new_n757), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1144), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1141), .A2(KEYINPUT121), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1142), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1134), .B(new_n1135), .C1(new_n735), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1097), .B1(new_n1125), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT118), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1101), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1117), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1125), .A2(new_n1128), .A3(KEYINPUT118), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1157), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1155), .B1(new_n1163), .B2(new_n730), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1133), .A2(new_n1164), .ZN(G378));
  NAND2_X1  g0965(.A1(new_n886), .A2(new_n902), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n698), .B1(new_n910), .B2(new_n900), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n309), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n300), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1168), .B1(new_n1169), .B2(new_n661), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n309), .A2(new_n300), .A3(new_n840), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1166), .A2(new_n1167), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1177), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1178), .A2(new_n1179), .A3(new_n930), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n930), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1177), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n874), .A2(new_n884), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n897), .B2(new_n920), .ZN(new_n1184));
  OAI21_X1  g0984(.A(G330), .B1(new_n1184), .B2(KEYINPUT40), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1182), .B1(new_n903), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1166), .A2(new_n1167), .A3(new_n1177), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1181), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(KEYINPUT57), .B1(new_n1180), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1092), .B1(new_n1163), .B2(new_n1114), .ZN(new_n1190));
  OAI21_X1  g0990(.A(KEYINPUT123), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT57), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1180), .A2(new_n1188), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n1190), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1092), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1099), .A2(new_n1113), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1195), .B1(new_n1131), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT123), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n930), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1186), .A2(new_n1181), .A3(new_n1187), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1198), .A2(new_n1199), .A3(KEYINPUT57), .A4(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1191), .A2(new_n1194), .A3(new_n684), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1182), .A2(new_n784), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n731), .B1(new_n939), .B2(new_n815), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1016), .B1(new_n751), .B2(new_n557), .C1(new_n447), .C2(new_n758), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G107), .A2(new_n820), .B1(new_n739), .B2(new_n428), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n263), .A2(G41), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n770), .C2(new_n742), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n767), .A2(new_n243), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(new_n1207), .A2(new_n1210), .A3(new_n1046), .A4(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT122), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1213), .A2(KEYINPUT58), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(KEYINPUT58), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(G33), .A2(G41), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1209), .A2(G50), .A3(new_n1216), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n747), .A2(new_n1149), .B1(new_n738), .B2(new_n822), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G132), .B2(new_n757), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n750), .A2(G125), .B1(G150), .B2(new_n1005), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n764), .C2(new_n1146), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n743), .A2(G124), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1216), .B(new_n1223), .C1(new_n767), .C2(new_n776), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1221), .B2(KEYINPUT59), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1217), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1214), .A2(new_n1215), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1206), .B1(new_n1227), .B2(new_n735), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1202), .A2(new_n730), .B1(new_n1205), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1204), .A2(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n1197), .A2(new_n1092), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n966), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1115), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n917), .A2(new_n784), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n731), .B1(G68), .B2(new_n815), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT124), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1044), .B1(new_n751), .B2(new_n754), .C1(new_n557), .C2(new_n758), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n272), .B1(new_n742), .B2(new_n552), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n747), .A2(new_n770), .B1(new_n738), .B2(new_n424), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(new_n765), .C2(G97), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1238), .B(new_n1241), .C1(new_n769), .C2(new_n373), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n750), .A2(G132), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT125), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1211), .B1(G159), .B2(new_n765), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n738), .A2(new_n823), .B1(new_n742), .B2(new_n1149), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n272), .B(new_n1246), .C1(G137), .C2(new_n820), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1146), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n757), .A2(new_n1248), .B1(G50), .B2(new_n1005), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1245), .A2(new_n1247), .A3(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1242), .B1(new_n1244), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1236), .B1(new_n1251), .B2(new_n735), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1196), .A2(new_n730), .B1(new_n1234), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1233), .A2(new_n1253), .ZN(G381));
  OR4_X1    g1054(.A1(G396), .A2(G384), .A3(G393), .A4(G390), .ZN(new_n1255));
  INV_X1    g1055(.A(G378), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1204), .A2(new_n1256), .A3(new_n1229), .ZN(new_n1257));
  OR4_X1    g1057(.A1(G387), .A2(new_n1255), .A3(G381), .A4(new_n1257), .ZN(G407));
  OAI211_X1 g1058(.A(G407), .B(G213), .C1(G343), .C2(new_n1257), .ZN(G409));
  NAND3_X1  g1059(.A1(new_n1000), .A2(new_n1029), .A3(G390), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT127), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(G393), .B(G396), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G387), .A2(new_n1068), .A3(new_n1088), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1260), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1265), .A2(new_n1263), .A3(KEYINPUT127), .A4(new_n1260), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1204), .A2(G378), .A3(new_n1229), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1198), .A2(new_n1232), .A3(new_n1202), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1229), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1256), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n662), .A2(G213), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1099), .A2(KEYINPUT60), .A3(new_n1092), .A4(new_n1113), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n684), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1115), .A2(KEYINPUT60), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1278), .B2(new_n1231), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(G384), .A2(new_n1280), .A3(new_n1253), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1253), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n813), .B(new_n836), .C1(new_n1279), .C2(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1274), .A2(new_n1275), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT126), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1270), .A2(new_n1273), .B1(G213), .B2(new_n662), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1288), .A3(new_n1284), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT62), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n662), .A2(G213), .A3(G2897), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1281), .A2(new_n1283), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT61), .B1(new_n1291), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1285), .A2(KEYINPUT62), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1269), .B1(new_n1290), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1286), .A2(new_n1300), .A3(new_n1289), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1287), .A2(KEYINPUT63), .A3(new_n1284), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .A4(new_n1296), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1299), .A2(new_n1304), .ZN(G405));
  NAND2_X1  g1105(.A1(G375), .A2(new_n1256), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1270), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1269), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1303), .A2(new_n1270), .A3(new_n1306), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1308), .A2(new_n1284), .A3(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1284), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(G402));
endmodule


