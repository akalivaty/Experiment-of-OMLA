//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT4), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT79), .B1(new_n189), .B2(G104), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT79), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G107), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n189), .A3(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n188), .B(G101), .C1(new_n194), .C2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT80), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n190), .A2(new_n193), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n195), .A3(new_n197), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n203), .A2(KEYINPUT80), .A3(new_n188), .A4(G101), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n202), .A2(new_n205), .A3(new_n195), .A4(new_n197), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n206), .A2(KEYINPUT4), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(G101), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n201), .A2(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n210));
  INV_X1    g024(.A(G113), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT67), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(KEYINPUT2), .B2(G113), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT2), .A2(G113), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G116), .B(G119), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT68), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G116), .ZN(new_n221));
  INV_X1    g035(.A(G116), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G119), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n221), .A2(new_n223), .A3(KEYINPUT68), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n217), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n226));
  AND4_X1   g040(.A1(new_n226), .A2(new_n215), .A3(new_n216), .A4(new_n218), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n212), .A2(new_n214), .B1(KEYINPUT2), .B2(G113), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n228), .B2(new_n218), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT70), .B(new_n225), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT69), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n226), .A3(new_n218), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT70), .B1(new_n235), .B2(new_n225), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n209), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT82), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n192), .A2(G107), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n189), .A2(G104), .ZN(new_n240));
  OAI21_X1  g054(.A(G101), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n206), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT5), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n219), .A2(new_n224), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n220), .A3(G116), .ZN(new_n245));
  OR2_X1    g059(.A1(new_n245), .A2(KEYINPUT83), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(KEYINPUT83), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(G113), .A3(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n235), .B(new_n242), .C1(new_n244), .C2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n230), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT82), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n209), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n238), .A2(new_n249), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G110), .B(G122), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT84), .ZN(new_n258));
  OR2_X1    g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n262), .A2(KEYINPUT64), .A3(G146), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT64), .B1(new_n262), .B2(G146), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT0), .ZN(new_n266));
  INV_X1    g080(.A(G128), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n267), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n262), .A2(G146), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n268), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G125), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n267), .A2(KEYINPUT1), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(new_n261), .A3(new_n272), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT64), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n260), .B2(G143), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n262), .A2(KEYINPUT64), .A3(G146), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n281), .A2(new_n282), .B1(G143), .B2(new_n260), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n267), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n279), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n277), .B1(new_n276), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G224), .ZN(new_n287));
  OR3_X1    g101(.A1(new_n287), .A2(KEYINPUT87), .A3(G953), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT87), .B1(new_n287), .B2(G953), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n289), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n235), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n248), .B1(KEYINPUT5), .B2(new_n218), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n242), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  XOR2_X1   g108(.A(new_n258), .B(KEYINPUT8), .Z(new_n295));
  OAI21_X1  g109(.A(new_n235), .B1(new_n244), .B2(new_n248), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n294), .B(new_n295), .C1(new_n296), .C2(new_n242), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n286), .A2(new_n290), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(KEYINPUT88), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n259), .A2(new_n291), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT6), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n256), .A2(new_n258), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n256), .B2(new_n258), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n256), .A2(new_n258), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n288), .A2(new_n289), .ZN(new_n308));
  XOR2_X1   g122(.A(new_n308), .B(KEYINPUT86), .Z(new_n309));
  XNOR2_X1  g123(.A(new_n286), .B(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n187), .B(new_n300), .C1(new_n307), .C2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G210), .B1(G237), .B2(G902), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(KEYINPUT89), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n256), .A2(new_n258), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n302), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n256), .A2(new_n258), .A3(new_n303), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n259), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(G902), .B1(new_n319), .B2(new_n310), .ZN(new_n320));
  INV_X1    g134(.A(new_n314), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(new_n300), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(G475), .ZN(new_n325));
  XNOR2_X1  g139(.A(G113), .B(G122), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(new_n192), .ZN(new_n327));
  XNOR2_X1  g141(.A(G125), .B(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT16), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n276), .A2(KEYINPUT16), .A3(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(G146), .A3(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(new_n328), .B(KEYINPUT19), .Z(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(G146), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT91), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G237), .ZN(new_n336));
  INV_X1    g150(.A(G953), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G214), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(G143), .ZN(new_n339));
  INV_X1    g153(.A(G131), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT91), .B(new_n331), .C1(new_n332), .C2(G146), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n335), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n328), .A2(new_n260), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT76), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n260), .B2(new_n328), .ZN(new_n346));
  AND4_X1   g160(.A1(KEYINPUT90), .A2(new_n339), .A3(KEYINPUT18), .A4(G131), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n339), .A2(KEYINPUT90), .B1(KEYINPUT18), .B2(G131), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n327), .B1(new_n343), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n329), .A2(new_n330), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(G146), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n339), .A2(new_n340), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT17), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n352), .B(new_n354), .C1(new_n341), .C2(KEYINPUT17), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n355), .A2(new_n349), .A3(new_n327), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n325), .B(new_n187), .C1(new_n350), .C2(new_n356), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n357), .A2(KEYINPUT92), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(KEYINPUT92), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(KEYINPUT20), .A3(new_n359), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n359), .A2(KEYINPUT20), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n327), .B1(new_n355), .B2(new_n349), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n187), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G475), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n360), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G952), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(G953), .ZN(new_n367));
  NAND2_X1  g181(.A1(G234), .A2(G237), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  XOR2_X1   g184(.A(KEYINPUT21), .B(G898), .Z(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(G902), .A3(G953), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT94), .B(KEYINPUT13), .Z(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(G128), .A3(new_n262), .ZN(new_n377));
  XNOR2_X1  g191(.A(G128), .B(G143), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n377), .B(G134), .C1(new_n379), .C2(new_n376), .ZN(new_n380));
  INV_X1    g194(.A(G134), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G122), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G116), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT93), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n222), .A2(G122), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(new_n189), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n385), .A2(new_n189), .A3(new_n386), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n380), .B(new_n382), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n385), .B1(KEYINPUT14), .B2(new_n386), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n386), .A2(KEYINPUT14), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(KEYINPUT95), .ZN(new_n393));
  OAI21_X1  g207(.A(G107), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n389), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n378), .B(new_n381), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(KEYINPUT9), .B(G234), .Z(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(G217), .A3(new_n337), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n398), .B(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n187), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT15), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G478), .ZN(new_n404));
  INV_X1    g218(.A(G478), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n401), .B(new_n187), .C1(KEYINPUT15), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n365), .A2(new_n375), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n323), .A2(new_n324), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G469), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n283), .A2(new_n268), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n411), .A2(new_n270), .B1(new_n273), .B2(new_n268), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n209), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT11), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n381), .B2(G137), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n381), .A2(G137), .ZN(new_n416));
  INV_X1    g230(.A(G137), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT11), .A3(G134), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G131), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT66), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT66), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n422), .A3(G131), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n417), .A2(KEYINPUT11), .A3(G134), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT11), .B1(new_n417), .B2(G134), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n340), .A4(new_n416), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n415), .A2(new_n418), .A3(new_n340), .A4(new_n416), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT65), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n421), .A2(new_n423), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n279), .B1(new_n273), .B2(new_n284), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n242), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT10), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n242), .A2(KEYINPUT10), .A3(new_n285), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n413), .A2(new_n431), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G140), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n337), .A2(G227), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n433), .B1(new_n285), .B2(new_n242), .ZN(new_n442));
  INV_X1    g256(.A(new_n431), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n442), .A2(KEYINPUT12), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT12), .B1(new_n442), .B2(new_n443), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n413), .A2(new_n435), .A3(new_n436), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n443), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n440), .B1(new_n449), .B2(new_n437), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n410), .B(new_n187), .C1(new_n447), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(G469), .A2(G902), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n437), .B1(new_n444), .B2(new_n445), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n440), .B(KEYINPUT78), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n437), .A3(new_n440), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n451), .B(new_n452), .C1(new_n410), .C2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G221), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n399), .B2(new_n187), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n458), .A2(KEYINPUT81), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT81), .B1(new_n458), .B2(new_n461), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n409), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G217), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n466), .B1(G234), .B2(new_n187), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT23), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n220), .B2(G128), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n267), .A2(KEYINPUT23), .A3(G119), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n470), .B(new_n471), .C1(G119), .C2(new_n267), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G110), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT75), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  XOR2_X1   g289(.A(KEYINPUT24), .B(G110), .Z(new_n476));
  XNOR2_X1  g290(.A(G119), .B(G128), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n479), .A2(new_n352), .ZN(new_n480));
  OAI22_X1  g294(.A1(new_n472), .A2(G110), .B1(new_n477), .B2(new_n476), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n345), .A2(new_n331), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT22), .B(G137), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n337), .A2(G221), .A3(G234), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n484), .B(new_n485), .Z(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n486), .B(new_n482), .C1(new_n479), .C2(new_n352), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n187), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT77), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT25), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n486), .B1(new_n480), .B2(new_n482), .ZN(new_n494));
  INV_X1    g308(.A(new_n489), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n492), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n187), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n468), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n467), .A2(G902), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G472), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT31), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n505));
  INV_X1    g319(.A(new_n416), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n381), .A2(G137), .ZN(new_n507));
  OAI21_X1  g321(.A(G131), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n429), .A2(KEYINPUT65), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n429), .A2(KEYINPUT65), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n285), .B(new_n508), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n505), .B(new_n511), .C1(new_n431), .C2(new_n275), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n419), .A2(new_n422), .A3(G131), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n422), .B1(new_n419), .B2(G131), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n429), .B(new_n427), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n412), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n505), .B1(new_n518), .B2(new_n511), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n253), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n252), .A2(new_n518), .A3(new_n230), .A4(new_n511), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n336), .A2(new_n337), .A3(G210), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(new_n205), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n520), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT71), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n511), .B1(new_n431), .B2(new_n275), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n253), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n421), .A2(new_n423), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n428), .A2(new_n430), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n275), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n511), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT30), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n512), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n530), .B1(new_n536), .B2(new_n253), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT71), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n526), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n504), .B1(new_n528), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n504), .A3(new_n526), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT28), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n253), .A2(new_n529), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n521), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n530), .A2(KEYINPUT28), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n525), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n503), .B(new_n187), .C1(new_n540), .C2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT32), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n538), .B1(new_n537), .B2(new_n526), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n535), .A2(new_n512), .B1(new_n252), .B2(new_n230), .ZN(new_n553));
  NOR4_X1   g367(.A1(new_n553), .A2(new_n530), .A3(KEYINPUT71), .A4(new_n525), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT31), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n541), .A2(new_n546), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n557), .A2(KEYINPUT32), .A3(new_n503), .A4(new_n187), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n550), .A2(new_n551), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n548), .A2(KEYINPUT72), .A3(new_n549), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n544), .A2(new_n545), .A3(new_n525), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT29), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n187), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT74), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT29), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT73), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n537), .A2(new_n526), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(KEYINPUT73), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n566), .B(new_n568), .C1(new_n570), .C2(new_n562), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT74), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n563), .A2(new_n572), .A3(new_n187), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n565), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G472), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n502), .B1(new_n561), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n465), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G101), .ZN(G3));
  OAI21_X1  g392(.A(new_n187), .B1(new_n540), .B2(new_n547), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n557), .A2(KEYINPUT96), .A3(new_n187), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(G472), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n583), .B2(new_n548), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n464), .A2(new_n502), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n324), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT98), .B1(new_n320), .B2(new_n300), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(new_n313), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n312), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n313), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n320), .A2(KEYINPUT98), .A3(new_n300), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT99), .B(G478), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n402), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n401), .A2(KEYINPUT33), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n401), .A2(KEYINPUT33), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n187), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n600), .B1(new_n603), .B2(new_n405), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n365), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n375), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n589), .A2(new_n598), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G104), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT100), .B(KEYINPUT34), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  XNOR2_X1  g424(.A(new_n375), .B(KEYINPUT101), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n365), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n407), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n589), .A2(new_n598), .A3(new_n612), .A4(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NAND2_X1  g432(.A1(new_n493), .A2(new_n498), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n467), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n480), .A2(new_n621), .A3(new_n482), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n480), .B2(new_n482), .ZN(new_n624));
  OAI22_X1  g438(.A1(new_n623), .A2(new_n624), .B1(KEYINPUT36), .B2(new_n487), .ZN(new_n625));
  INV_X1    g439(.A(new_n624), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n487), .A2(KEYINPUT36), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n622), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n625), .A2(new_n628), .A3(new_n500), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n620), .A2(KEYINPUT103), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n631));
  INV_X1    g445(.A(new_n629), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n631), .B1(new_n499), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n587), .A2(new_n465), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT37), .B(G110), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  AOI21_X1  g452(.A(new_n464), .B1(new_n561), .B2(new_n575), .ZN(new_n639));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n374), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n369), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n614), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n639), .A2(new_n598), .A3(new_n635), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  XNOR2_X1  g460(.A(new_n323), .B(KEYINPUT38), .ZN(new_n647));
  INV_X1    g461(.A(new_n407), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n613), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n649), .A2(new_n324), .A3(new_n634), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n552), .A2(new_n554), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n543), .A2(new_n521), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n652), .B2(new_n525), .ZN(new_n653));
  OAI21_X1  g467(.A(G472), .B1(new_n653), .B2(G902), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n561), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n647), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(KEYINPUT104), .ZN(new_n657));
  INV_X1    g471(.A(new_n464), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n642), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(KEYINPUT40), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n656), .A2(KEYINPUT104), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n657), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  NOR2_X1   g479(.A1(new_n605), .A2(new_n643), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n639), .A2(new_n598), .A3(new_n635), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G146), .ZN(G48));
  OR2_X1    g482(.A1(new_n447), .A2(new_n450), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(G469), .B1(new_n670), .B2(G902), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n451), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n460), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n592), .A2(new_n597), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n576), .A2(new_n674), .A3(new_n606), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NOR3_X1   g491(.A1(new_n365), .A2(new_n648), .A3(new_n611), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n576), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G116), .ZN(G18));
  NAND2_X1  g494(.A1(new_n561), .A2(new_n575), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n674), .A2(new_n681), .A3(new_n408), .A4(new_n635), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G119), .ZN(G21));
  AOI21_X1  g497(.A(KEYINPUT106), .B1(new_n579), .B2(G472), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n548), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n557), .A2(KEYINPUT106), .A3(new_n503), .A4(new_n187), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n502), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n674), .A2(new_n612), .A3(new_n649), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G122), .ZN(G24));
  AOI21_X1  g503(.A(new_n634), .B1(new_n685), .B2(new_n686), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n674), .A2(new_n666), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT107), .B(G125), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G27));
  NAND3_X1  g507(.A1(new_n575), .A2(new_n550), .A3(new_n558), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n452), .B(KEYINPUT108), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n451), .B(new_n695), .C1(new_n410), .C2(new_n457), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n696), .A2(new_n461), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n694), .A2(KEYINPUT42), .A3(new_n501), .A4(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n315), .A2(new_n324), .A3(new_n322), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n666), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n576), .A2(new_n666), .A3(new_n697), .A4(new_n700), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n340), .ZN(G33));
  AND4_X1   g520(.A1(new_n576), .A2(new_n644), .A3(new_n697), .A4(new_n700), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n381), .ZN(G36));
  NAND2_X1  g522(.A1(new_n613), .A2(new_n604), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT43), .Z(new_n710));
  OAI211_X1 g524(.A(new_n710), .B(new_n635), .C1(new_n586), .C2(new_n585), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n699), .B1(new_n712), .B2(KEYINPUT44), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n457), .B(KEYINPUT45), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G469), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n695), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n715), .A2(KEYINPUT46), .A3(new_n695), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n451), .A3(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n720), .A2(new_n461), .A3(new_n660), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n713), .B(new_n721), .C1(KEYINPUT44), .C2(new_n712), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT109), .B(G137), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G39));
  NAND2_X1  g538(.A1(new_n720), .A2(new_n461), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n701), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n725), .A2(new_n729), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n681), .A2(new_n501), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  OR3_X1    g550(.A1(new_n734), .A2(KEYINPUT111), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT111), .B1(new_n734), .B2(new_n736), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G140), .ZN(G42));
  AND3_X1   g554(.A1(new_n592), .A2(new_n597), .A3(new_n649), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n499), .A2(new_n632), .A3(new_n643), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n655), .A3(new_n697), .A4(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n645), .A2(new_n667), .A3(new_n743), .A4(new_n691), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n559), .A2(new_n560), .B1(G472), .B2(new_n574), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n464), .A3(new_n634), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n748), .B(new_n598), .C1(new_n644), .C2(new_n666), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(KEYINPUT52), .A3(new_n691), .A4(new_n743), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n323), .A2(new_n324), .A3(new_n678), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT113), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n323), .A2(new_n754), .A3(new_n678), .A4(new_n324), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n587), .A2(new_n753), .A3(new_n588), .A4(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n636), .A3(new_n688), .A4(new_n682), .ZN(new_n757));
  INV_X1    g571(.A(new_n605), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n323), .A2(new_n324), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n587), .A2(new_n588), .A3(new_n612), .A4(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(new_n675), .A3(new_n679), .A4(new_n577), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n705), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n747), .A2(new_n502), .A3(new_n699), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n644), .A3(new_n697), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n690), .A2(new_n666), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n634), .A2(new_n407), .A3(new_n365), .A4(new_n643), .ZN(new_n768));
  AOI22_X1  g582(.A1(new_n767), .A2(new_n697), .B1(new_n639), .B2(new_n768), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n764), .B(new_n766), .C1(new_n769), .C2(new_n699), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n681), .A2(new_n768), .A3(new_n658), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n690), .A2(new_n666), .A3(new_n697), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n699), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT114), .B1(new_n773), .B2(new_n707), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n762), .A2(new_n763), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n751), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n773), .A2(new_n707), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n705), .B1(new_n778), .B2(new_n764), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(KEYINPUT115), .A3(new_n762), .A4(new_n774), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT53), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n746), .A2(new_n750), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT53), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n775), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n781), .A2(KEYINPUT54), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n757), .ZN(new_n786));
  AND4_X1   g600(.A1(new_n577), .A2(new_n760), .A3(new_n675), .A4(new_n679), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n787), .A3(new_n774), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n770), .A2(new_n763), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n776), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n780), .A3(new_n782), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT116), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n777), .A2(new_n795), .A3(KEYINPUT53), .A4(new_n780), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n785), .B1(new_n797), .B2(KEYINPUT54), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n710), .A2(new_n370), .A3(new_n687), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n674), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n699), .A2(new_n460), .A3(new_n369), .A4(new_n672), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n710), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n694), .A2(new_n501), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT48), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(KEYINPUT118), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(KEYINPUT118), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n806), .A2(KEYINPUT118), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n803), .A2(new_n804), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n655), .A2(new_n502), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(new_n802), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n758), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n807), .A2(new_n367), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n604), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n812), .A2(new_n613), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n647), .A2(new_n324), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n800), .A2(new_n673), .A3(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n819));
  AOI21_X1  g633(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n803), .A2(new_n690), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n818), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n731), .A2(new_n733), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n672), .B(KEYINPUT112), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n461), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n700), .B(new_n800), .C1(new_n823), .C2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT51), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT51), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n814), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n798), .A2(new_n801), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n366), .A2(new_n337), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n798), .A2(KEYINPUT119), .A3(new_n830), .A4(new_n801), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n824), .A2(KEYINPUT49), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n824), .A2(KEYINPUT49), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n837), .A2(new_n838), .A3(new_n647), .A4(new_n709), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(new_n461), .A3(new_n324), .A4(new_n811), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n840), .ZN(G75));
  AOI21_X1  g655(.A(new_n784), .B1(new_n791), .B2(new_n792), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n187), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(G210), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n319), .B(new_n311), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT55), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n847), .B1(new_n844), .B2(new_n845), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n337), .A2(G952), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(G51));
  INV_X1    g665(.A(new_n850), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT120), .B1(new_n842), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n842), .A2(new_n853), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n856), .B(KEYINPUT54), .C1(new_n781), .C2(new_n784), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n695), .B(KEYINPUT57), .Z(new_n859));
  AOI21_X1  g673(.A(new_n670), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n842), .A2(new_n187), .A3(new_n715), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n852), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g678(.A(KEYINPUT121), .B(new_n852), .C1(new_n860), .C2(new_n861), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(G54));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n843), .A2(KEYINPUT58), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(G475), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n350), .A2(new_n356), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n867), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n871), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n868), .A2(KEYINPUT122), .A3(G475), .A4(new_n870), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n852), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(G60));
  NOR2_X1   g689(.A1(new_n601), .A2(new_n602), .ZN(new_n876));
  NAND2_X1  g690(.A1(G478), .A2(G902), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT59), .Z(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n798), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n852), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n876), .A2(new_n878), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n858), .B2(new_n881), .ZN(G63));
  INV_X1    g696(.A(new_n842), .ZN(new_n883));
  XNOR2_X1  g697(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n466), .A2(new_n187), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n883), .A2(new_n628), .A3(new_n625), .A4(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n883), .A2(new_n886), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n852), .B(new_n887), .C1(new_n888), .C2(new_n496), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g706(.A(G953), .B1(new_n372), .B2(new_n287), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n762), .B2(G953), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n307), .B1(G898), .B2(new_n337), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT125), .Z(new_n896));
  XNOR2_X1  g710(.A(new_n894), .B(new_n896), .ZN(G69));
  AOI21_X1  g711(.A(new_n337), .B1(G227), .B2(G900), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n721), .A2(new_n804), .A3(new_n741), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n739), .A2(new_n722), .A3(new_n766), .A4(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n749), .A2(new_n691), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n763), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n901), .A2(G953), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n640), .A2(new_n337), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n536), .B(new_n332), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n906), .B(KEYINPUT126), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n664), .A2(new_n902), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT62), .Z(new_n912));
  INV_X1    g726(.A(new_n661), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n765), .B(new_n913), .C1(new_n758), .C2(new_n615), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n912), .A2(new_n722), .A3(new_n739), .A4(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n910), .B1(new_n915), .B2(new_n337), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT127), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n908), .A2(new_n916), .A3(KEYINPUT127), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n899), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n919), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n898), .A3(new_n917), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(G72));
  NAND2_X1  g737(.A1(G472), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT63), .Z(new_n925));
  INV_X1    g739(.A(new_n762), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n915), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n927), .B(new_n526), .C1(new_n530), .C2(new_n553), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n901), .A2(new_n926), .A3(new_n903), .ZN(new_n929));
  INV_X1    g743(.A(new_n925), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n525), .B(new_n537), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n797), .B(new_n925), .C1(new_n569), .C2(new_n651), .ZN(new_n932));
  AND4_X1   g746(.A1(new_n852), .A2(new_n928), .A3(new_n931), .A4(new_n932), .ZN(G57));
endmodule


