//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT66), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n469), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n470));
  OR2_X1    g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n466), .A2(new_n472), .A3(G2105), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n468), .A2(new_n471), .A3(new_n473), .ZN(G160));
  AND3_X1   g049(.A1(new_n461), .A2(new_n463), .A3(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G136), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n469), .A2(new_n478), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n476), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT67), .Z(G162));
  NAND4_X1  g058(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n478), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT69), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n469), .A2(new_n486), .A3(G138), .A4(new_n478), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n485), .A2(new_n487), .A3(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(new_n478), .B2(G114), .ZN(new_n490));
  NOR2_X1   g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n491), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n493), .A2(new_n495), .A3(KEYINPUT68), .A4(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n484), .A2(KEYINPUT69), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n469), .A2(G126), .A3(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n488), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(G543), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n510), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n519), .B(new_n521), .C1(new_n512), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n515), .A2(KEYINPUT70), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n511), .A2(new_n525), .A3(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n523), .B1(G51), .B2(new_n527), .ZN(G168));
  AND3_X1   g103(.A1(new_n507), .A2(G90), .A3(new_n511), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n526), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n525), .B1(new_n511), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n504), .A2(new_n506), .A3(G64), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n509), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT71), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n534), .B1(new_n524), .B2(new_n526), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n529), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n542));
  INV_X1    g117(.A(new_n538), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n539), .A2(new_n544), .ZN(G171));
  AND3_X1   g120(.A1(new_n507), .A2(G81), .A3(new_n511), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n504), .A2(new_n506), .A3(G56), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n509), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n547), .B(new_n551), .C1(new_n533), .C2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n546), .B1(new_n527), .B2(G43), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n556), .A2(KEYINPUT72), .A3(new_n551), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT73), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G188));
  NOR2_X1   g140(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n515), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n569), .B2(new_n512), .ZN(new_n570));
  AND2_X1   g145(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n571));
  NOR4_X1   g146(.A1(new_n515), .A2(new_n567), .A3(new_n571), .A4(new_n566), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n504), .A2(new_n506), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(KEYINPUT75), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(KEYINPUT75), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(G651), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n573), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  INV_X1    g157(.A(G168), .ZN(G286));
  INV_X1    g158(.A(new_n512), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G87), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n511), .A2(G49), .A3(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(new_n507), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n593));
  INV_X1    g168(.A(G48), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n515), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n511), .A2(KEYINPUT76), .A3(G48), .A4(G543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n584), .A2(G86), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n592), .A2(new_n597), .A3(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n509), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT77), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n527), .A2(G47), .B1(G85), .B2(new_n584), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n575), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n527), .A2(G54), .B1(G651), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n584), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n512), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT79), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT78), .B1(new_n615), .B2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NOR2_X1   g192(.A1(G171), .A2(new_n617), .ZN(new_n618));
  MUX2_X1   g193(.A(new_n616), .B(KEYINPUT78), .S(new_n618), .Z(G284));
  MUX2_X1   g194(.A(new_n616), .B(KEYINPUT78), .S(new_n618), .Z(G321));
  NAND2_X1  g195(.A1(G299), .A2(new_n617), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n617), .B2(G168), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(new_n617), .B2(G168), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n615), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n615), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g204(.A1(new_n464), .A2(G2105), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G2104), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT80), .B(KEYINPUT13), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n630), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n475), .A2(G123), .ZN(new_n637));
  NOR2_X1   g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(new_n478), .B2(G111), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT81), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n635), .A2(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2435), .ZN(new_n645));
  XOR2_X1   g220(.A(G2427), .B(G2438), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT14), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G1341), .B(G1348), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G14), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n658), .B1(new_n662), .B2(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2096), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  AOI21_X1  g242(.A(KEYINPUT18), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n665), .B(new_n668), .Z(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT82), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n679), .A2(new_n671), .A3(new_n674), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n677), .B(new_n680), .C1(new_n671), .C2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT22), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  MUX2_X1   g264(.A(G6), .B(G305), .S(G16), .Z(new_n690));
  XOR2_X1   g265(.A(KEYINPUT32), .B(G1981), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G22), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G166), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G1971), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(G1971), .ZN(new_n697));
  NOR2_X1   g272(.A1(G16), .A2(G23), .ZN(new_n698));
  INV_X1    g273(.A(G288), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G16), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT33), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n692), .A2(new_n696), .A3(new_n697), .A4(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT34), .Z(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G25), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n630), .A2(G131), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n475), .A2(G119), .ZN(new_n708));
  OR2_X1    g283(.A1(G95), .A2(G2105), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n709), .B(G2104), .C1(G107), .C2(new_n478), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(new_n705), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G290), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(new_n693), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n693), .B2(G24), .ZN(new_n718));
  INV_X1    g293(.A(G1986), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n715), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n719), .B2(new_n718), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n704), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(KEYINPUT83), .A2(KEYINPUT36), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n722), .B(new_n723), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n705), .A2(G32), .ZN(new_n725));
  NAND2_X1  g300(.A1(G105), .A2(G2104), .ZN(new_n726));
  INV_X1    g301(.A(G141), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n464), .B2(new_n727), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n728), .A2(new_n478), .B1(G129), .B2(new_n475), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT26), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n725), .B1(new_n733), .B2(new_n705), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT27), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1996), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n693), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n693), .ZN(new_n738));
  INV_X1    g313(.A(G1966), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n693), .A2(G4), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n615), .B2(new_n693), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1348), .ZN(new_n743));
  NOR2_X1   g318(.A1(G29), .A2(G35), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G162), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT29), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n743), .B1(G2090), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n705), .A2(G27), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n705), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT88), .B(G2078), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G19), .ZN(new_n752));
  OAI21_X1  g327(.A(KEYINPUT84), .B1(new_n752), .B2(G16), .ZN(new_n753));
  OR3_X1    g328(.A1(new_n752), .A2(KEYINPUT84), .A3(G16), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n753), .B(new_n754), .C1(new_n558), .C2(new_n693), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1341), .ZN(new_n756));
  NOR2_X1   g331(.A1(G5), .A2(G16), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G171), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1961), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n630), .A2(G139), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n761), .B(new_n762), .C1(new_n478), .C2(new_n763), .ZN(new_n764));
  MUX2_X1   g339(.A(G33), .B(new_n764), .S(G29), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2072), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n756), .A2(new_n759), .A3(new_n766), .ZN(new_n767));
  AND4_X1   g342(.A1(new_n740), .A2(new_n747), .A3(new_n751), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n641), .A2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT85), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G28), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT86), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n774), .B(new_n705), .C1(new_n772), .C2(G28), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n769), .A2(new_n771), .A3(new_n775), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT87), .Z(new_n777));
  NOR2_X1   g352(.A1(new_n746), .A2(G2090), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n705), .A2(G26), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n630), .A2(G140), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n475), .A2(G128), .ZN(new_n783));
  NOR2_X1   g358(.A1(G104), .A2(G2105), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(new_n478), .B2(G116), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n781), .B1(new_n786), .B2(G29), .ZN(new_n787));
  MUX2_X1   g362(.A(new_n781), .B(new_n787), .S(KEYINPUT28), .Z(new_n788));
  INV_X1    g363(.A(G2067), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G34), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(KEYINPUT24), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(KEYINPUT24), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n705), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G160), .B2(new_n705), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2084), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n780), .A2(new_n790), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n724), .A2(new_n736), .A3(new_n768), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n778), .A2(new_n779), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(G299), .A2(G16), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n693), .A2(KEYINPUT23), .A3(G20), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT23), .ZN(new_n803));
  INV_X1    g378(.A(G20), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G16), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1956), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n798), .A2(new_n800), .A3(new_n807), .ZN(G311));
  AND3_X1   g383(.A1(new_n724), .A2(new_n768), .A3(new_n797), .ZN(new_n809));
  INV_X1    g384(.A(new_n807), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n809), .A2(new_n799), .A3(new_n810), .A4(new_n736), .ZN(G150));
  NAND2_X1  g386(.A1(G80), .A2(G543), .ZN(new_n812));
  INV_X1    g387(.A(G67), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n575), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G651), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n527), .A2(G55), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT90), .B(G93), .Z(new_n817));
  AND3_X1   g392(.A1(new_n507), .A2(new_n817), .A3(new_n511), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(KEYINPUT91), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n524), .B2(new_n526), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n822), .A2(new_n823), .A3(new_n818), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n815), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n615), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT39), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT92), .B(KEYINPUT38), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n553), .B(new_n815), .C1(new_n820), .C2(new_n824), .ZN(new_n832));
  AOI21_X1  g407(.A(KEYINPUT72), .B1(new_n556), .B2(new_n551), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n552), .B1(new_n524), .B2(new_n526), .ZN(new_n834));
  NOR4_X1   g409(.A1(new_n834), .A2(new_n546), .A3(new_n554), .A4(new_n550), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n816), .A2(KEYINPUT91), .A3(new_n819), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n823), .B1(new_n822), .B2(new_n818), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n837), .A2(new_n838), .B1(G651), .B2(new_n814), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n832), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n831), .B(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n827), .B1(new_n842), .B2(G860), .ZN(G145));
  INV_X1    g418(.A(KEYINPUT93), .ZN(new_n844));
  XNOR2_X1  g419(.A(G162), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n641), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G160), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n630), .A2(KEYINPUT95), .A3(G142), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n849));
  INV_X1    g424(.A(G142), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n481), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n475), .A2(G130), .ZN(new_n852));
  OR2_X1    g427(.A1(G106), .A2(G2105), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(G2104), .C1(G118), .C2(new_n478), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n848), .A2(new_n851), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n711), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT96), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n632), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT97), .Z(new_n859));
  XOR2_X1   g434(.A(new_n732), .B(new_n786), .Z(new_n860));
  INV_X1    g435(.A(KEYINPUT94), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n488), .B2(new_n501), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n492), .A2(new_n496), .B1(new_n475), .B2(G126), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n485), .A2(new_n487), .A3(KEYINPUT4), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT94), .A4(new_n499), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n860), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n764), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n859), .A2(new_n868), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n847), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n847), .B(KEYINPUT98), .ZN(new_n873));
  INV_X1    g448(.A(new_n868), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n858), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT40), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT40), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n872), .A2(new_n876), .A3(new_n880), .A4(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(G395));
  XNOR2_X1  g457(.A(G303), .B(G288), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n883), .A2(G305), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(G305), .ZN(new_n885));
  OAI21_X1  g460(.A(G290), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n883), .A2(G305), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(G305), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n716), .A3(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT100), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT42), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n841), .B(new_n626), .ZN(new_n893));
  NAND2_X1  g468(.A1(G299), .A2(new_n614), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n573), .A2(new_n580), .A3(new_n608), .A4(new_n613), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n896), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT41), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n893), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n898), .B(KEYINPUT99), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n892), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n891), .B(KEYINPUT42), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n902), .B2(new_n900), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(G868), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT101), .B1(new_n825), .B2(new_n617), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(new_n907), .ZN(G295));
  AOI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n907), .ZN(G331));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n913));
  XNOR2_X1  g488(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n542), .B1(new_n541), .B2(new_n543), .ZN(new_n916));
  NOR4_X1   g491(.A1(new_n540), .A2(new_n529), .A3(KEYINPUT71), .A4(new_n538), .ZN(new_n917));
  OAI21_X1  g492(.A(G286), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n539), .A2(new_n544), .A3(G168), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n840), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n558), .A2(new_n825), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n922), .A2(new_n832), .A3(new_n919), .A4(new_n918), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(KEYINPUT103), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n899), .A2(new_n897), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n918), .A2(new_n919), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n841), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n886), .A2(new_n889), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n921), .A2(new_n923), .A3(new_n894), .A4(new_n896), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n932), .A2(new_n877), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n929), .A2(new_n931), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n890), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n915), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n877), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n924), .A2(new_n928), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n898), .A2(KEYINPUT104), .A3(KEYINPUT41), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n921), .B2(new_n923), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n899), .A2(KEYINPUT104), .A3(new_n897), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n939), .A2(new_n901), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n938), .B1(new_n943), .B2(new_n930), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n942), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n901), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n924), .B2(new_n928), .ZN(new_n948));
  OAI211_X1 g523(.A(KEYINPUT105), .B(new_n890), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n937), .B1(new_n944), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n936), .B1(new_n950), .B2(new_n915), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n913), .B1(new_n951), .B2(KEYINPUT44), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n953));
  AOI211_X1 g528(.A(new_n914), .B(new_n937), .C1(new_n944), .C2(new_n949), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT106), .B(new_n953), .C1(new_n954), .C2(new_n936), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n944), .A2(new_n949), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n933), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n950), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(KEYINPUT43), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n933), .A2(new_n935), .A3(new_n915), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(KEYINPUT44), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n956), .A2(new_n964), .ZN(G397));
  XNOR2_X1  g540(.A(KEYINPUT108), .B(G1384), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n862), .B2(new_n865), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n968));
  AND4_X1   g543(.A1(G40), .A2(new_n468), .A3(new_n471), .A4(new_n473), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n786), .B(new_n789), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n732), .A2(G1996), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n732), .A2(G1996), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n711), .B(new_n714), .Z(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(G290), .B(G1986), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n971), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT109), .Z(new_n981));
  NAND2_X1  g556(.A1(G286), .A2(G8), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT51), .B1(new_n982), .B2(KEYINPUT120), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n488), .B2(new_n501), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n863), .A2(new_n864), .A3(new_n499), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n989), .A3(new_n985), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n987), .A2(new_n969), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G2084), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n986), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n988), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(new_n969), .A3(new_n995), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n991), .A2(new_n992), .B1(new_n996), .B2(new_n739), .ZN(new_n997));
  INV_X1    g572(.A(G8), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n982), .B(new_n984), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n994), .A2(new_n969), .A3(new_n995), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n987), .A2(new_n969), .A3(new_n990), .ZN(new_n1001));
  OAI22_X1  g576(.A1(new_n1000), .A2(G1966), .B1(G2084), .B2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(G8), .B(new_n983), .C1(new_n1002), .C2(G286), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(G8), .A3(G286), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n999), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1005), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT125), .B1(new_n1005), .B2(KEYINPUT62), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OR2_X1    g583(.A1(G305), .A2(G1981), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT114), .B(G86), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n507), .A2(new_n511), .A3(new_n1010), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n597), .A2(KEYINPUT115), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT115), .B1(new_n597), .B2(new_n1011), .ZN(new_n1013));
  INV_X1    g588(.A(new_n592), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1981), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT49), .B(new_n1009), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT116), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1009), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n986), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n998), .B1(new_n969), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n597), .A2(new_n1011), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n597), .A2(KEYINPUT115), .A3(new_n1011), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n592), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G1981), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1029), .A2(new_n1030), .A3(KEYINPUT49), .A4(new_n1009), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1018), .A2(new_n1021), .A3(new_n1023), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1976), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G288), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(new_n1023), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT113), .B1(new_n699), .B2(G1976), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1023), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1023), .B(new_n1037), .C1(KEYINPUT52), .C2(new_n1035), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1032), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n970), .B1(new_n994), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n994), .A2(new_n1043), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n1047));
  INV_X1    g622(.A(new_n966), .ZN(new_n1048));
  AND4_X1   g623(.A1(new_n1047), .A2(new_n866), .A3(KEYINPUT45), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1047), .B1(new_n967), .B2(KEYINPUT45), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1044), .B(new_n1046), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1971), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1001), .A2(G2090), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n998), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(G166), .B2(new_n998), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1042), .B1(new_n1056), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1063), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1001), .A2(KEYINPUT118), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n1067));
  AOI21_X1  g642(.A(G2090), .B1(new_n991), .B2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1051), .A2(new_n1052), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1065), .B1(new_n1069), .B2(new_n998), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n991), .A2(G1961), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT94), .B1(new_n1072), .B2(new_n864), .ZN(new_n1073));
  AND4_X1   g648(.A1(KEYINPUT94), .A2(new_n863), .A3(new_n864), .A4(new_n499), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT45), .B(new_n1048), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT111), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n967), .A2(new_n1047), .A3(KEYINPUT45), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G2078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1071), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1000), .A2(KEYINPUT53), .A3(new_n1079), .ZN(new_n1083));
  AOI21_X1  g658(.A(G301), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n999), .A2(new_n1003), .A3(new_n1085), .A4(new_n1004), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1064), .A2(new_n1070), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT126), .B1(new_n1008), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1045), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1089));
  AOI21_X1  g664(.A(G1971), .B1(new_n1089), .B2(new_n1044), .ZN(new_n1090));
  OAI211_X1 g665(.A(G8), .B(new_n1063), .C1(new_n1090), .C2(new_n1054), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1032), .A2(new_n1041), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1070), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1071), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(new_n1083), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(new_n1086), .A3(G171), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT125), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1005), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1098), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1088), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1091), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1032), .A2(new_n1033), .A3(new_n699), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1009), .ZN(new_n1109));
  XOR2_X1   g684(.A(new_n1023), .B(KEYINPUT117), .Z(new_n1110));
  AOI22_X1  g685(.A1(new_n1107), .A2(new_n1092), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n997), .A2(new_n998), .A3(G286), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1070), .A2(new_n1091), .A3(new_n1092), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT63), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT119), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1117), .A3(new_n1114), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1056), .A2(new_n1063), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1119), .A2(new_n1064), .A3(KEYINPUT63), .A4(new_n1112), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1116), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1106), .A2(new_n1111), .A3(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT56), .B(G2072), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1078), .A2(new_n1044), .A3(new_n1046), .A4(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(G299), .B(KEYINPUT57), .Z(new_n1125));
  OR2_X1    g700(.A1(new_n991), .A2(G1956), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n969), .A2(new_n1022), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n991), .A2(G1348), .B1(G2067), .B2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1127), .A2(new_n615), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1125), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT61), .B1(new_n1132), .B2(new_n1131), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1123), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1126), .B1(new_n1051), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1125), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(new_n1138), .A3(new_n1127), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT58), .B(G1341), .Z(new_n1140));
  NAND2_X1  g715(.A1(new_n1128), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1051), .B2(G1996), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n558), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT59), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1142), .A2(new_n1145), .A3(new_n558), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1133), .A2(new_n1139), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n615), .A2(KEYINPUT60), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(new_n1129), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n615), .A2(KEYINPUT60), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1149), .B(new_n1150), .Z(new_n1151));
  AOI211_X1 g726(.A(new_n1130), .B(new_n1131), .C1(new_n1147), .C2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n1154));
  OAI21_X1  g729(.A(G40), .B1(new_n1154), .B2(G2078), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n478), .B1(new_n466), .B2(KEYINPUT122), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(KEYINPUT122), .B2(new_n466), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n471), .B(KEYINPUT53), .C1(KEYINPUT123), .C2(new_n1079), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1156), .A2(new_n968), .A3(new_n1158), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1155), .B(new_n1159), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1164), .A2(KEYINPUT124), .A3(new_n968), .A4(new_n1158), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1082), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(G171), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1153), .B1(new_n1167), .B2(new_n1084), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(G171), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1082), .A2(G301), .A3(new_n1083), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1169), .A2(new_n1170), .A3(KEYINPUT54), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1093), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1168), .A2(new_n1171), .A3(new_n1172), .A4(new_n1005), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1152), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n981), .B1(new_n1122), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n971), .A2(new_n719), .A3(new_n716), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT48), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1177), .A2(new_n977), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n968), .A2(G1996), .A3(new_n970), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1179), .A2(KEYINPUT46), .ZN(new_n1180));
  INV_X1    g755(.A(new_n972), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n971), .B1(new_n732), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(KEYINPUT46), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1180), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT47), .Z(new_n1185));
  NAND2_X1  g760(.A1(new_n712), .A2(new_n714), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT127), .Z(new_n1187));
  OAI22_X1  g762(.A1(new_n1187), .A2(new_n975), .B1(G2067), .B2(new_n786), .ZN(new_n1188));
  AOI211_X1 g763(.A(new_n1178), .B(new_n1185), .C1(new_n971), .C2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1175), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g765(.A1(G401), .A2(G227), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n878), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g767(.A(new_n936), .ZN(new_n1194));
  OAI21_X1  g768(.A(new_n1194), .B1(new_n958), .B2(new_n914), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n688), .A2(new_n1195), .A3(G319), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n1193), .A2(new_n1196), .ZN(G308));
  AND2_X1   g771(.A1(new_n1195), .A2(G319), .ZN(new_n1198));
  NAND4_X1  g772(.A1(new_n1198), .A2(new_n688), .A3(new_n878), .A4(new_n1192), .ZN(G225));
endmodule


