

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590;

  XNOR2_X1 U326 ( .A(n341), .B(n340), .ZN(n343) );
  XNOR2_X1 U327 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U328 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n394) );
  XNOR2_X1 U329 ( .A(n395), .B(n394), .ZN(n524) );
  NOR2_X1 U330 ( .A1(n514), .A2(n413), .ZN(n576) );
  INV_X1 U331 ( .A(G183GAT), .ZN(n451) );
  XNOR2_X1 U332 ( .A(n449), .B(n448), .ZN(n526) );
  XOR2_X1 U333 ( .A(KEYINPUT28), .B(n459), .Z(n529) );
  XNOR2_X1 U334 ( .A(n451), .B(KEYINPUT124), .ZN(n452) );
  XNOR2_X1 U335 ( .A(n453), .B(n452), .ZN(G1350GAT) );
  XOR2_X1 U336 ( .A(G64GAT), .B(G211GAT), .Z(n295) );
  XNOR2_X1 U337 ( .A(G22GAT), .B(G78GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U339 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n297) );
  XNOR2_X1 U340 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n310) );
  XOR2_X1 U343 ( .A(G57GAT), .B(KEYINPUT13), .Z(n366) );
  XOR2_X1 U344 ( .A(G155GAT), .B(G71GAT), .Z(n301) );
  XNOR2_X1 U345 ( .A(G127GAT), .B(G183GAT), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U347 ( .A(n366), .B(n302), .Z(n304) );
  NAND2_X1 U348 ( .A1(G231GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U350 ( .A(n305), .B(KEYINPUT76), .Z(n308) );
  XNOR2_X1 U351 ( .A(G15GAT), .B(G1GAT), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n306), .B(KEYINPUT67), .ZN(n374) );
  XNOR2_X1 U353 ( .A(n374), .B(KEYINPUT15), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n310), .B(n309), .ZN(n585) );
  XOR2_X1 U356 ( .A(KEYINPUT6), .B(G148GAT), .Z(n312) );
  XNOR2_X1 U357 ( .A(G141GAT), .B(G1GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U359 ( .A(G85GAT), .B(G162GAT), .Z(n314) );
  XNOR2_X1 U360 ( .A(G29GAT), .B(G120GAT), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n334) );
  XOR2_X1 U363 ( .A(G57GAT), .B(KEYINPUT1), .Z(n318) );
  XNOR2_X1 U364 ( .A(KEYINPUT92), .B(KEYINPUT88), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U366 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n320) );
  XNOR2_X1 U367 ( .A(KEYINPUT91), .B(KEYINPUT89), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U369 ( .A(n322), .B(n321), .Z(n332) );
  XOR2_X1 U370 ( .A(KEYINPUT79), .B(G134GAT), .Z(n324) );
  XNOR2_X1 U371 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U373 ( .A(G113GAT), .B(n325), .Z(n436) );
  XOR2_X1 U374 ( .A(G155GAT), .B(KEYINPUT86), .Z(n327) );
  XNOR2_X1 U375 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n327), .B(n326), .ZN(n424) );
  XOR2_X1 U377 ( .A(n424), .B(KEYINPUT4), .Z(n329) );
  NAND2_X1 U378 ( .A1(G225GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n436), .B(n330), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U382 ( .A(n334), .B(n333), .ZN(n514) );
  XOR2_X1 U383 ( .A(G92GAT), .B(G85GAT), .Z(n336) );
  XNOR2_X1 U384 ( .A(G99GAT), .B(G106GAT), .ZN(n335) );
  XNOR2_X1 U385 ( .A(n336), .B(n335), .ZN(n359) );
  INV_X1 U386 ( .A(KEYINPUT11), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n359), .B(n337), .ZN(n341) );
  NAND2_X1 U388 ( .A1(G232GAT), .A2(G233GAT), .ZN(n339) );
  INV_X1 U389 ( .A(KEYINPUT73), .ZN(n338) );
  XOR2_X1 U390 ( .A(G36GAT), .B(G190GAT), .Z(n401) );
  XNOR2_X1 U391 ( .A(n401), .B(KEYINPUT74), .ZN(n342) );
  XNOR2_X1 U392 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U393 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n345) );
  XNOR2_X1 U394 ( .A(G134GAT), .B(KEYINPUT72), .ZN(n344) );
  XNOR2_X1 U395 ( .A(n345), .B(n344), .ZN(n346) );
  OR2_X1 U396 ( .A1(n347), .A2(n346), .ZN(n349) );
  NAND2_X1 U397 ( .A1(n347), .A2(n346), .ZN(n348) );
  NAND2_X1 U398 ( .A1(n349), .A2(n348), .ZN(n355) );
  XOR2_X1 U399 ( .A(G29GAT), .B(G43GAT), .Z(n351) );
  XNOR2_X1 U400 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n350) );
  XNOR2_X1 U401 ( .A(n351), .B(n350), .ZN(n375) );
  XOR2_X1 U402 ( .A(G162GAT), .B(KEYINPUT71), .Z(n353) );
  XNOR2_X1 U403 ( .A(G50GAT), .B(G218GAT), .ZN(n352) );
  XNOR2_X1 U404 ( .A(n353), .B(n352), .ZN(n425) );
  XOR2_X1 U405 ( .A(n375), .B(n425), .Z(n354) );
  XNOR2_X1 U406 ( .A(n355), .B(n354), .ZN(n387) );
  XNOR2_X1 U407 ( .A(n387), .B(KEYINPUT75), .ZN(n570) );
  XNOR2_X1 U408 ( .A(n570), .B(KEYINPUT36), .ZN(n485) );
  NOR2_X1 U409 ( .A1(n485), .A2(n585), .ZN(n356) );
  XNOR2_X1 U410 ( .A(KEYINPUT45), .B(n356), .ZN(n385) );
  XOR2_X1 U411 ( .A(KEYINPUT32), .B(KEYINPUT70), .Z(n358) );
  XNOR2_X1 U412 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n360) );
  XOR2_X1 U414 ( .A(n360), .B(n359), .Z(n362) );
  XOR2_X1 U415 ( .A(G120GAT), .B(G71GAT), .Z(n432) );
  XOR2_X1 U416 ( .A(G148GAT), .B(G78GAT), .Z(n416) );
  XNOR2_X1 U417 ( .A(n432), .B(n416), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n370) );
  XOR2_X1 U419 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n364) );
  NAND2_X1 U420 ( .A1(G230GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U422 ( .A(n365), .B(KEYINPUT68), .Z(n368) );
  XOR2_X1 U423 ( .A(G176GAT), .B(G64GAT), .Z(n396) );
  XNOR2_X1 U424 ( .A(n366), .B(n396), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U426 ( .A(n370), .B(n369), .Z(n581) );
  INV_X1 U427 ( .A(n581), .ZN(n454) );
  XOR2_X1 U428 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n372) );
  NAND2_X1 U429 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U431 ( .A(n373), .B(KEYINPUT30), .Z(n377) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U434 ( .A(G197GAT), .B(G113GAT), .Z(n379) );
  XNOR2_X1 U435 ( .A(G36GAT), .B(G50GAT), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U437 ( .A(n381), .B(n380), .Z(n383) );
  XOR2_X1 U438 ( .A(G141GAT), .B(G22GAT), .Z(n414) );
  XOR2_X1 U439 ( .A(G169GAT), .B(G8GAT), .Z(n397) );
  XNOR2_X1 U440 ( .A(n414), .B(n397), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n577) );
  INV_X1 U442 ( .A(n577), .ZN(n549) );
  NOR2_X1 U443 ( .A1(n454), .A2(n549), .ZN(n384) );
  AND2_X1 U444 ( .A1(n385), .A2(n384), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n386), .B(KEYINPUT112), .ZN(n393) );
  XOR2_X1 U446 ( .A(KEYINPUT41), .B(n581), .Z(n564) );
  INV_X1 U447 ( .A(n564), .ZN(n553) );
  NAND2_X1 U448 ( .A1(n549), .A2(n553), .ZN(n388) );
  XNOR2_X1 U449 ( .A(KEYINPUT46), .B(n388), .ZN(n389) );
  NAND2_X1 U450 ( .A1(n389), .A2(n585), .ZN(n390) );
  NOR2_X1 U451 ( .A1(n387), .A2(n390), .ZN(n391) );
  XOR2_X1 U452 ( .A(KEYINPUT47), .B(n391), .Z(n392) );
  NOR2_X1 U453 ( .A1(n393), .A2(n392), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n411) );
  XOR2_X1 U455 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n399) );
  XNOR2_X1 U456 ( .A(G218GAT), .B(G92GAT), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U458 ( .A(n401), .B(n400), .Z(n403) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n409) );
  XOR2_X1 U461 ( .A(G183GAT), .B(KEYINPUT19), .Z(n405) );
  XNOR2_X1 U462 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n431) );
  XOR2_X1 U464 ( .A(G204GAT), .B(G211GAT), .Z(n407) );
  XNOR2_X1 U465 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(n406), .ZN(n417) );
  XOR2_X1 U467 ( .A(n431), .B(n417), .Z(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n475) );
  NOR2_X1 U470 ( .A1(n524), .A2(n475), .ZN(n412) );
  XOR2_X1 U471 ( .A(KEYINPUT54), .B(n412), .Z(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(G106GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n415), .B(KEYINPUT23), .ZN(n429) );
  XOR2_X1 U474 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U477 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n421) );
  XNOR2_X1 U478 ( .A(KEYINPUT85), .B(KEYINPUT24), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U480 ( .A(n423), .B(n422), .Z(n427) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n459) );
  NAND2_X1 U484 ( .A1(n576), .A2(n459), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n430), .B(KEYINPUT55), .ZN(n450) );
  XOR2_X1 U486 ( .A(n432), .B(n431), .Z(n434) );
  XNOR2_X1 U487 ( .A(G43GAT), .B(G99GAT), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n449) );
  XOR2_X1 U490 ( .A(G176GAT), .B(G190GAT), .Z(n438) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(G15GAT), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U493 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n440) );
  XNOR2_X1 U494 ( .A(KEYINPUT20), .B(KEYINPUT82), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n442), .B(n441), .Z(n447) );
  XOR2_X1 U497 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n444) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U500 ( .A(KEYINPUT65), .B(n445), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n448) );
  NAND2_X1 U502 ( .A1(n450), .A2(n526), .ZN(n571) );
  NOR2_X1 U503 ( .A1(n585), .A2(n571), .ZN(n453) );
  NOR2_X1 U504 ( .A1(n577), .A2(n454), .ZN(n489) );
  XOR2_X1 U505 ( .A(KEYINPUT27), .B(n475), .Z(n461) );
  NAND2_X1 U506 ( .A1(n514), .A2(n461), .ZN(n525) );
  NOR2_X1 U507 ( .A1(n525), .A2(n529), .ZN(n531) );
  XNOR2_X1 U508 ( .A(KEYINPUT95), .B(n531), .ZN(n455) );
  NOR2_X1 U509 ( .A1(n526), .A2(n455), .ZN(n467) );
  INV_X1 U510 ( .A(n526), .ZN(n533) );
  NOR2_X1 U511 ( .A1(n533), .A2(n475), .ZN(n456) );
  XOR2_X1 U512 ( .A(KEYINPUT96), .B(n456), .Z(n457) );
  NAND2_X1 U513 ( .A1(n457), .A2(n459), .ZN(n458) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(n458), .Z(n463) );
  NOR2_X1 U515 ( .A1(n459), .A2(n526), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n460), .B(KEYINPUT26), .ZN(n575) );
  NAND2_X1 U517 ( .A1(n575), .A2(n461), .ZN(n462) );
  NAND2_X1 U518 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U519 ( .A(KEYINPUT97), .B(n464), .ZN(n465) );
  NOR2_X1 U520 ( .A1(n514), .A2(n465), .ZN(n466) );
  NOR2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n486) );
  INV_X1 U522 ( .A(n585), .ZN(n558) );
  NAND2_X1 U523 ( .A1(n570), .A2(n558), .ZN(n468) );
  XNOR2_X1 U524 ( .A(n468), .B(KEYINPUT16), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT78), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n486), .A2(n470), .ZN(n501) );
  AND2_X1 U527 ( .A1(n489), .A2(n501), .ZN(n482) );
  NAND2_X1 U528 ( .A1(n482), .A2(n514), .ZN(n474) );
  XOR2_X1 U529 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n472) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(G1324GAT) );
  INV_X1 U533 ( .A(n475), .ZN(n517) );
  NAND2_X1 U534 ( .A1(n482), .A2(n517), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(KEYINPUT100), .ZN(n477) );
  XNOR2_X1 U536 ( .A(G8GAT), .B(n477), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n479) );
  NAND2_X1 U538 ( .A1(n482), .A2(n526), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(n481) );
  XOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT101), .Z(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  XOR2_X1 U542 ( .A(G22GAT), .B(KEYINPUT103), .Z(n484) );
  NAND2_X1 U543 ( .A1(n482), .A2(n529), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1327GAT) );
  NOR2_X1 U545 ( .A1(n485), .A2(n486), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n585), .A2(n487), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n488), .ZN(n513) );
  NAND2_X1 U548 ( .A1(n489), .A2(n513), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(KEYINPUT38), .ZN(n491) );
  XNOR2_X1 U550 ( .A(KEYINPUT105), .B(n491), .ZN(n499) );
  NAND2_X1 U551 ( .A1(n514), .A2(n499), .ZN(n493) );
  XOR2_X1 U552 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(n494), .ZN(G1328GAT) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(KEYINPUT106), .ZN(n496) );
  NAND2_X1 U556 ( .A1(n517), .A2(n499), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n499), .A2(n526), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U561 ( .A1(n499), .A2(n529), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n503) );
  NOR2_X1 U564 ( .A1(n564), .A2(n549), .ZN(n512) );
  AND2_X1 U565 ( .A1(n512), .A2(n501), .ZN(n508) );
  NAND2_X1 U566 ( .A1(n508), .A2(n514), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n508), .A2(n517), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n505), .B(KEYINPUT108), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n508), .A2(n526), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U575 ( .A1(n508), .A2(n529), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U577 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n516) );
  AND2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n521) );
  NAND2_X1 U580 ( .A1(n514), .A2(n521), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  XOR2_X1 U582 ( .A(G92GAT), .B(KEYINPUT111), .Z(n519) );
  NAND2_X1 U583 ( .A1(n521), .A2(n517), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n526), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n529), .A2(n521), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  XNOR2_X1 U590 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n524), .A2(n525), .ZN(n547) );
  NAND2_X1 U592 ( .A1(n526), .A2(n547), .ZN(n527) );
  NAND2_X1 U593 ( .A1(KEYINPUT113), .A2(n527), .ZN(n528) );
  NOR2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n535) );
  NOR2_X1 U595 ( .A1(n524), .A2(KEYINPUT113), .ZN(n530) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n544) );
  NOR2_X1 U599 ( .A1(n577), .A2(n544), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XNOR2_X1 U602 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n540) );
  NOR2_X1 U603 ( .A1(n564), .A2(n544), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  NOR2_X1 U606 ( .A1(n585), .A2(n544), .ZN(n542) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(n542), .Z(n543) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  NOR2_X1 U609 ( .A1(n544), .A2(n570), .ZN(n546) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n551) );
  NAND2_X1 U613 ( .A1(n575), .A2(n547), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n548), .B(KEYINPUT117), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n561), .A2(n549), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n557) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  NAND2_X1 U620 ( .A1(n561), .A2(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  XOR2_X1 U623 ( .A(G155GAT), .B(KEYINPUT121), .Z(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n387), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U628 ( .A1(n577), .A2(n571), .ZN(n563) );
  XOR2_X1 U629 ( .A(G169GAT), .B(n563), .Z(G1348GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n571), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n566) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(KEYINPUT122), .B(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  INV_X1 U636 ( .A(KEYINPUT58), .ZN(n573) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(n574), .ZN(G1351GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n588) );
  NOR2_X1 U641 ( .A1(n577), .A2(n588), .ZN(n579) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n588), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT61), .B(KEYINPUT125), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n584), .Z(G1353GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n588), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT126), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n485), .A2(n588), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

