//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  AND2_X1   g0012(.A1(KEYINPUT65), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(KEYINPUT65), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT68), .Z(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT67), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G50), .ZN(new_n227));
  INV_X1    g0027(.A(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT66), .B(G77), .ZN(new_n229));
  INV_X1    g0029(.A(G244), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n208), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n212), .B(new_n220), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G226), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT69), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G107), .ZN(new_n246));
  INV_X1    g0046(.A(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n216), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT72), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n255), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n254), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n255), .A2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT12), .ZN(new_n264));
  OAI21_X1  g0064(.A(G68), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n259), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n266), .A2(new_n264), .A3(G68), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(new_n264), .B2(new_n266), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G68), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n269), .A2(G50), .B1(G20), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n215), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n254), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT11), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n265), .A2(new_n268), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n228), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n238), .A2(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G97), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT13), .ZN(new_n289));
  OR2_X1    g0089(.A1(KEYINPUT70), .A2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT70), .A2(G45), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G1), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(G1), .A2(G13), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G41), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G238), .A3(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n288), .A2(new_n289), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n299), .B1(new_n284), .B2(new_n285), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n296), .A2(new_n301), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT13), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(G169), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n303), .A2(G179), .A3(new_n306), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n308), .B1(new_n307), .B2(G169), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n279), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT75), .ZN(new_n314));
  INV_X1    g0114(.A(new_n254), .ZN(new_n315));
  OR2_X1    g0115(.A1(KEYINPUT65), .A2(G20), .ZN(new_n316));
  NAND2_X1  g0116(.A1(KEYINPUT65), .A2(G20), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT15), .B(G87), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n229), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n320), .A2(new_n322), .B1(new_n323), .B2(new_n318), .ZN(new_n324));
  INV_X1    g0124(.A(new_n269), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(KEYINPUT74), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT8), .B(G58), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT74), .B1(G20), .B2(G33), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OR3_X1    g0129(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n315), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n266), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n229), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n260), .A2(G77), .A3(new_n261), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n314), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT73), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n293), .A2(new_n295), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n299), .A2(G244), .A3(new_n300), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G238), .A2(G1698), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n280), .B(new_n341), .C1(new_n238), .C2(G1698), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(new_n287), .C1(G107), .C2(new_n280), .ZN(new_n343));
  INV_X1    g0143(.A(G45), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n291), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n255), .A2(new_n345), .B1(new_n297), .B2(new_n298), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G244), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT73), .A3(new_n296), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n340), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G200), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n272), .A2(new_n321), .B1(new_n229), .B2(new_n215), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n254), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n353), .A2(KEYINPUT75), .A3(new_n333), .A4(new_n334), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n340), .A2(new_n343), .A3(G190), .A4(new_n348), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n336), .A2(new_n350), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n333), .A3(new_n334), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n358), .B(new_n359), .C1(G179), .C2(new_n349), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n307), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G200), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n303), .B2(new_n306), .ZN(new_n365));
  OR3_X1    g0165(.A1(new_n363), .A2(new_n279), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n313), .A2(new_n361), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n260), .A2(G50), .A3(new_n261), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n332), .A2(new_n227), .ZN(new_n369));
  INV_X1    g0169(.A(G150), .ZN(new_n370));
  INV_X1    g0170(.A(G20), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n370), .A2(new_n325), .B1(new_n201), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G58), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n373), .A2(KEYINPUT71), .A3(KEYINPUT8), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT71), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n327), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n372), .B1(new_n376), .B2(new_n320), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n368), .B(new_n369), .C1(new_n377), .C2(new_n315), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G33), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n229), .ZN(new_n383));
  MUX2_X1   g0183(.A(G222), .B(G223), .S(G1698), .Z(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n287), .C1(new_n382), .C2(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n346), .A2(G226), .B1(new_n293), .B2(new_n295), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n357), .ZN(new_n388));
  INV_X1    g0188(.A(G179), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n378), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n376), .A2(new_n320), .ZN(new_n392));
  INV_X1    g0192(.A(new_n372), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n254), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT9), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(new_n396), .A3(new_n368), .A4(new_n369), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n378), .A2(KEYINPUT9), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT10), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n387), .A2(new_n362), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(G200), .B2(new_n387), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n400), .B1(new_n399), .B2(new_n402), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n391), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n367), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT78), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  OR2_X1    g0209(.A1(G223), .A2(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n228), .A2(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n409), .B1(new_n412), .B2(new_n382), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n287), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n346), .A2(G232), .B1(new_n293), .B2(new_n295), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n362), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT77), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT77), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n414), .A2(new_n415), .A3(new_n418), .A4(new_n362), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n414), .A2(new_n415), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n364), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT16), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT76), .B1(new_n319), .B2(KEYINPUT3), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT76), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(new_n380), .A3(G33), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n426), .A3(new_n379), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT7), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n213), .A2(new_n214), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n280), .B2(G20), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n270), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(G58), .B(G68), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G20), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n269), .A2(G159), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n423), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n433), .A2(G20), .B1(G159), .B2(new_n269), .ZN(new_n438));
  AOI21_X1  g0238(.A(G20), .B1(new_n379), .B2(new_n381), .ZN(new_n439));
  OAI21_X1  g0239(.A(G68), .B1(new_n439), .B2(new_n428), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n318), .A2(new_n280), .A3(KEYINPUT7), .ZN(new_n441));
  OAI211_X1 g0241(.A(KEYINPUT16), .B(new_n438), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n437), .A2(new_n254), .A3(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n376), .A2(new_n266), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n263), .B2(new_n376), .ZN(new_n445));
  AND4_X1   g0245(.A1(new_n408), .A2(new_n422), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n444), .ZN(new_n447));
  INV_X1    g0247(.A(new_n376), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n262), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n380), .A2(G33), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n371), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n270), .B1(new_n452), .B2(KEYINPUT7), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n382), .A2(new_n215), .A3(new_n428), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n436), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n315), .B1(new_n455), .B2(KEYINPUT16), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n449), .B1(new_n456), .B2(new_n437), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n408), .B1(new_n457), .B2(new_n422), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n446), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n420), .A2(G169), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n414), .A2(G179), .A3(new_n415), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT18), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n430), .A2(new_n431), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G68), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT16), .B1(new_n465), .B2(new_n438), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n442), .A2(new_n254), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n445), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT18), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n460), .A2(new_n461), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n407), .B1(new_n459), .B2(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n457), .A2(KEYINPUT18), .A3(new_n462), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n469), .B1(new_n468), .B2(new_n470), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n422), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT17), .B1(new_n477), .B2(new_n468), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n457), .A2(new_n408), .A3(new_n422), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n480), .A3(KEYINPUT78), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n406), .A2(new_n473), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n319), .A2(G97), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n316), .A2(new_n483), .A3(new_n317), .A4(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n253), .A2(new_n216), .B1(G20), .B2(new_n247), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT20), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n255), .A2(G33), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n266), .A2(G116), .A3(new_n315), .A4(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n258), .A2(new_n247), .A3(new_n259), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n485), .A2(KEYINPUT85), .A3(new_n486), .A4(new_n488), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT86), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n495), .A2(new_n494), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n499), .A2(KEYINPUT86), .A3(new_n493), .A4(new_n491), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n281), .A2(G257), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G264), .A2(G1698), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n280), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G303), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n382), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n506), .A3(new_n287), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n344), .A2(G1), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G41), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n291), .A2(KEYINPUT5), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(G270), .A3(new_n299), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT5), .B(G41), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n344), .A2(new_n294), .A3(G1), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n515), .A3(new_n299), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n507), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G169), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n501), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT21), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n501), .A2(KEYINPUT21), .A3(new_n519), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n517), .A2(new_n389), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n501), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n517), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G190), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n517), .A2(G200), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n527), .A2(new_n498), .A3(new_n500), .A4(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n522), .A2(new_n523), .A3(new_n525), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n215), .A2(G33), .A3(G97), .ZN(new_n531));
  OR2_X1    g0331(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n532));
  NAND2_X1  g0332(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G87), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n204), .A3(new_n205), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n285), .B1(new_n532), .B2(new_n533), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n318), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n215), .A2(new_n280), .A3(G68), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(new_n254), .B1(new_n332), .B2(new_n321), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n266), .A2(new_n315), .A3(new_n492), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT80), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n260), .A2(KEYINPUT80), .A3(new_n492), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(G87), .A3(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G238), .A2(G1698), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n230), .A2(G1698), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n550), .A2(new_n379), .A3(new_n381), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G116), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n299), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G250), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n255), .B2(G45), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n299), .B1(new_n515), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT82), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT82), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n549), .B1(new_n230), .B2(G1698), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n280), .B1(G33), .B2(G116), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n560), .B(new_n557), .C1(new_n562), .C2(new_n299), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n362), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n559), .A2(new_n563), .A3(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n548), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n542), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n545), .A2(new_n322), .A3(new_n546), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT84), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n260), .A2(KEYINPUT80), .A3(new_n492), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT80), .B1(new_n260), .B2(new_n492), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT84), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n574), .A3(new_n322), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n568), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n559), .A2(new_n563), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n389), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(G169), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n567), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n316), .A2(new_n379), .A3(new_n381), .A4(new_n317), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT22), .B1(new_n581), .B2(new_n536), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT22), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n215), .A2(new_n280), .A3(new_n583), .A4(G87), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  NAND2_X1  g0386(.A1(KEYINPUT23), .A2(G107), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(G20), .ZN(new_n589));
  NOR2_X1   g0389(.A1(KEYINPUT23), .A2(G107), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n318), .A2(KEYINPUT87), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n213), .B2(new_n214), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n589), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n585), .A2(new_n586), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n586), .B1(new_n585), .B2(new_n595), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n254), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n258), .A2(new_n205), .A3(new_n259), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n599), .B(KEYINPUT25), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n573), .B2(G107), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(G257), .A2(G1698), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n379), .A2(new_n381), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT88), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G294), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n379), .A2(new_n381), .A3(G250), .A4(new_n281), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT88), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n379), .A2(new_n381), .A3(new_n603), .A4(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT89), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n607), .A2(new_n606), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT89), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n605), .A4(new_n609), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n614), .A3(new_n287), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n287), .B1(new_n514), .B2(new_n508), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G264), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n516), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n357), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n299), .B1(new_n610), .B2(KEYINPUT89), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n618), .B1(new_n622), .B2(new_n614), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n389), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n602), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(G200), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n615), .A2(G190), .A3(new_n619), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n626), .A2(new_n598), .A3(new_n601), .A4(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n512), .A2(G257), .A3(new_n299), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n230), .A2(G1698), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(new_n379), .A3(new_n381), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT4), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT81), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n630), .A2(new_n379), .A3(new_n381), .A4(new_n633), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n635), .A2(new_n636), .A3(new_n484), .A4(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n629), .B1(new_n638), .B2(new_n287), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n516), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n357), .ZN(new_n641));
  INV_X1    g0441(.A(new_n516), .ZN(new_n642));
  AOI211_X1 g0442(.A(new_n642), .B(new_n629), .C1(new_n638), .C2(new_n287), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n389), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n205), .B1(new_n430), .B2(new_n431), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n205), .A2(G97), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT6), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(KEYINPUT79), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT79), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(KEYINPUT6), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n646), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(KEYINPUT6), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(KEYINPUT79), .ZN(new_n653));
  NAND2_X1  g0453(.A1(G97), .A2(G107), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n206), .A2(new_n652), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n651), .A2(new_n655), .A3(new_n318), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n269), .A2(G77), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n254), .B1(new_n645), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n545), .A2(G97), .A3(new_n546), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n332), .A2(new_n204), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n641), .A2(new_n644), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n638), .A2(new_n287), .ZN(new_n664));
  INV_X1    g0464(.A(new_n629), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n664), .A2(new_n362), .A3(new_n516), .A4(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n643), .B2(G200), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n659), .A2(new_n661), .A3(new_n660), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n625), .A2(new_n628), .A3(new_n663), .A4(new_n669), .ZN(new_n670));
  NOR4_X1   g0470(.A1(new_n482), .A2(new_n530), .A3(new_n580), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT90), .ZN(G372));
  INV_X1    g0472(.A(new_n391), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n360), .A2(KEYINPUT91), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n360), .A2(KEYINPUT91), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n366), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n313), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT92), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT92), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n676), .A2(new_n679), .A3(new_n313), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n678), .A2(new_n480), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n476), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n403), .A2(new_n404), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n673), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n482), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n574), .B1(new_n573), .B2(new_n322), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n569), .A2(KEYINPUT84), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n542), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n554), .A2(new_n558), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n577), .A2(new_n389), .B1(new_n690), .B2(new_n357), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n520), .A2(new_n521), .B1(new_n501), .B2(new_n524), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n625), .A3(new_n523), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n689), .A2(new_n364), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n564), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n548), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n628), .A2(new_n663), .A3(new_n669), .A4(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n692), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT26), .ZN(new_n701));
  INV_X1    g0501(.A(new_n691), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n698), .B1(new_n576), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n703), .B2(new_n663), .ZN(new_n704));
  INV_X1    g0504(.A(new_n579), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n688), .ZN(new_n706));
  INV_X1    g0506(.A(new_n663), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(KEYINPUT26), .A3(new_n567), .A4(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n685), .B1(new_n700), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n684), .A2(new_n710), .ZN(G369));
  XOR2_X1   g0511(.A(KEYINPUT94), .B(G330), .Z(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n693), .A2(new_n523), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n215), .A2(new_n255), .A3(G13), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n715), .A2(KEYINPUT27), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(KEYINPUT27), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G213), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G343), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n501), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n714), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT93), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n530), .A2(new_n721), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n722), .A2(KEYINPUT93), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n713), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n627), .B1(new_n364), .B2(new_n623), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n602), .ZN(new_n729));
  INV_X1    g0529(.A(new_n720), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n598), .B2(new_n601), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n625), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n602), .A2(new_n621), .A3(new_n624), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n730), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n727), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n714), .A2(new_n730), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n736), .A2(new_n739), .ZN(G399));
  INV_X1    g0540(.A(new_n209), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G41), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n255), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n537), .A2(G116), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n743), .A2(new_n744), .B1(new_n219), .B2(new_n742), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT28), .Z(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n524), .A2(new_n577), .A3(new_n639), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n748), .B2(new_n620), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n526), .A2(new_n639), .A3(G179), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(KEYINPUT30), .A3(new_n577), .A4(new_n623), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n526), .A2(G179), .A3(new_n689), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(new_n620), .A3(new_n640), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n749), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n754), .A2(KEYINPUT31), .A3(new_n720), .ZN(new_n755));
  AOI21_X1  g0555(.A(KEYINPUT31), .B1(new_n754), .B2(new_n720), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n669), .B(new_n663), .C1(new_n728), .C2(new_n602), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n733), .ZN(new_n759));
  INV_X1    g0559(.A(new_n530), .ZN(new_n760));
  INV_X1    g0560(.A(new_n580), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(new_n730), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n712), .B1(new_n757), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n730), .B1(new_n700), .B2(new_n709), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT29), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n692), .A2(new_n707), .A3(KEYINPUT26), .A4(new_n698), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT95), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n542), .A2(new_n547), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n770), .A2(new_n564), .A3(new_n696), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n688), .B2(new_n691), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n772), .A2(KEYINPUT95), .A3(KEYINPUT26), .A4(new_n707), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n701), .B1(new_n580), .B2(new_n663), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n769), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n692), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n758), .A2(new_n771), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(new_n777), .B2(new_n694), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(KEYINPUT29), .A3(new_n730), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n763), .B1(new_n766), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n746), .B1(new_n781), .B2(G1), .ZN(G364));
  INV_X1    g0582(.A(G13), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n318), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G45), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n743), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n727), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n725), .A2(new_n726), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n713), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n216), .B1(G20), .B2(new_n357), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n251), .A2(G45), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT97), .Z(new_n796));
  NOR2_X1   g0596(.A1(new_n741), .A2(new_n280), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n290), .A2(new_n292), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n218), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n741), .A2(new_n382), .ZN(new_n801));
  NAND2_X1  g0601(.A1(G355), .A2(KEYINPUT96), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G355), .A2(KEYINPUT96), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n803), .A2(new_n804), .B1(G116), .B2(new_n209), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n794), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n786), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n215), .A2(new_n389), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n809), .A2(new_n362), .A3(new_n364), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT98), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n809), .A2(G190), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(G200), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n815), .A2(new_n323), .B1(G58), .B2(new_n817), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(KEYINPUT99), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(KEYINPUT99), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G179), .A2(G200), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n318), .A2(new_n362), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G159), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT32), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n362), .A2(G179), .A3(G200), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n215), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n204), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n364), .A2(G179), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n829), .A2(G20), .A3(G190), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n280), .B1(new_n830), .B2(new_n536), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n389), .A2(new_n364), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n318), .A2(new_n362), .A3(new_n833), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n318), .A2(new_n362), .A3(new_n829), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n832), .B1(new_n270), .B2(new_n834), .C1(new_n205), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n816), .A2(new_n364), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n825), .B(new_n837), .C1(G50), .C2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n819), .A2(new_n820), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT100), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n815), .A2(G311), .ZN(new_n843));
  INV_X1    g0643(.A(G294), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n382), .B1(new_n505), .B2(new_n830), .C1(new_n827), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G283), .B2(new_n835), .ZN(new_n846));
  INV_X1    g0646(.A(new_n834), .ZN(new_n847));
  XNOR2_X1  g0647(.A(KEYINPUT33), .B(G317), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G329), .A2(new_n823), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G322), .A2(new_n817), .B1(new_n838), .B2(G326), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n843), .A2(new_n846), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n840), .A2(new_n841), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n842), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n808), .B1(new_n853), .B2(new_n793), .ZN(new_n854));
  INV_X1    g0654(.A(new_n792), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n854), .B1(new_n788), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n789), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G396));
  OAI211_X1 g0658(.A(new_n361), .B(new_n730), .C1(new_n700), .C2(new_n709), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n704), .A2(new_n708), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n720), .B1(new_n778), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n674), .A2(new_n359), .A3(new_n675), .A4(new_n720), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n720), .A2(new_n359), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n361), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n859), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n763), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n807), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n867), .B2(new_n866), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n793), .A2(new_n790), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n807), .B1(G77), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n815), .A2(G116), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n382), .B1(new_n830), .B2(new_n205), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n874), .B(new_n828), .C1(G283), .C2(new_n847), .ZN(new_n875));
  AOI22_X1  g0675(.A1(G311), .A2(new_n823), .B1(new_n835), .B2(G87), .ZN(new_n876));
  AOI22_X1  g0676(.A1(G294), .A2(new_n817), .B1(new_n838), .B2(G303), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n873), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n817), .A2(G143), .B1(G150), .B2(new_n847), .ZN(new_n879));
  INV_X1    g0679(.A(G137), .ZN(new_n880));
  INV_X1    g0680(.A(new_n838), .ZN(new_n881));
  INV_X1    g0681(.A(G159), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n879), .B1(new_n880), .B2(new_n881), .C1(new_n814), .C2(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT34), .Z(new_n884));
  NOR2_X1   g0684(.A1(new_n836), .A2(new_n270), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n280), .B1(new_n830), .B2(new_n227), .ZN(new_n887));
  INV_X1    g0687(.A(new_n827), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(new_n888), .B2(G58), .ZN(new_n889));
  INV_X1    g0689(.A(G132), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n886), .B(new_n889), .C1(new_n890), .C2(new_n822), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n878), .B1(new_n884), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n872), .B1(new_n892), .B2(new_n793), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n791), .B2(new_n865), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n869), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(G384));
  NAND2_X1  g0696(.A1(new_n651), .A2(new_n655), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT35), .ZN(new_n898));
  OAI211_X1 g0698(.A(G116), .B(new_n217), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n898), .B2(new_n897), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT36), .Z(new_n901));
  AOI211_X1 g0701(.A(new_n218), .B(new_n229), .C1(G58), .C2(G68), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n270), .A2(G50), .ZN(new_n903));
  OAI211_X1 g0703(.A(G1), .B(new_n783), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT101), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT102), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n453), .A2(new_n454), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT16), .B1(new_n908), .B2(new_n438), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n445), .B1(new_n467), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n718), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n459), .B2(new_n472), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n457), .A2(new_n422), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n910), .A2(new_n470), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n916), .A3(new_n912), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n468), .A2(new_n470), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n468), .A2(new_n911), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n915), .A2(new_n919), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n914), .A2(new_n923), .A3(KEYINPUT38), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT38), .B1(new_n914), .B2(new_n923), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n907), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n914), .A2(new_n923), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT38), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n914), .A2(new_n923), .A3(KEYINPUT38), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(KEYINPUT102), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n360), .A2(new_n720), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n859), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n279), .A2(new_n720), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n313), .A2(new_n366), .A3(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n279), .B(new_n720), .C1(new_n311), .C2(new_n312), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n932), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n472), .A2(new_n718), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n313), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n730), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n920), .B1(new_n476), .B2(new_n480), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n915), .A2(new_n919), .A3(new_n920), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT37), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n946), .A2(KEYINPUT103), .B1(new_n922), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT103), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n459), .A2(new_n472), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n920), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT38), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT39), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n930), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT104), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n920), .ZN(new_n957));
  OAI211_X1 g0757(.A(KEYINPUT103), .B(new_n957), .C1(new_n459), .C2(new_n472), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n948), .A2(new_n922), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n476), .A2(new_n480), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT103), .B1(new_n961), .B2(new_n957), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n928), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n961), .A2(new_n913), .B1(new_n922), .B2(new_n918), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT39), .B1(new_n964), .B2(KEYINPUT38), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT104), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n954), .B1(new_n929), .B2(new_n930), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n956), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n942), .B1(new_n945), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n766), .A2(new_n780), .A3(new_n685), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n684), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n971), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n757), .A2(new_n762), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n862), .A2(new_n864), .B1(new_n937), .B2(new_n938), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n926), .B2(new_n931), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT40), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n963), .A2(new_n930), .ZN(new_n980));
  NOR4_X1   g0780(.A1(new_n670), .A2(new_n530), .A3(new_n580), .A4(new_n720), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n754), .A2(new_n720), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT31), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n754), .A2(KEYINPUT31), .A3(new_n720), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n976), .B(KEYINPUT40), .C1(new_n981), .C2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n980), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n979), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n482), .B1(new_n762), .B2(new_n757), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n713), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n992), .B2(new_n990), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n974), .A2(new_n994), .B1(new_n255), .B2(new_n784), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n974), .A2(new_n994), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n906), .B1(new_n995), .B2(new_n996), .ZN(G367));
  OAI21_X1  g0797(.A(new_n794), .B1(new_n209), .B2(new_n321), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n242), .B2(new_n797), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n815), .A2(G50), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n280), .B1(new_n830), .B2(new_n373), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n827), .A2(new_n270), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(G159), .C2(new_n847), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G137), .A2(new_n823), .B1(new_n835), .B2(new_n323), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G143), .A2(new_n838), .B1(new_n817), .B2(G150), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1000), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n830), .A2(new_n247), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT46), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n280), .B(new_n1008), .C1(G107), .C2(new_n888), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n835), .A2(G97), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n844), .B2(new_n834), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G317), .B2(new_n823), .ZN(new_n1012));
  INV_X1    g0812(.A(G283), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1009), .B(new_n1012), .C1(new_n1013), .C2(new_n814), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G303), .A2(new_n817), .B1(new_n838), .B2(G311), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT110), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1006), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT47), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n786), .B(new_n999), .C1(new_n1018), .C2(new_n793), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n770), .A2(new_n720), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT105), .Z(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n776), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n703), .B2(new_n1021), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1019), .B1(new_n855), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n785), .A2(G1), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n727), .A2(KEYINPUT109), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n735), .B(new_n737), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n727), .B2(KEYINPUT109), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1026), .B(new_n1028), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n669), .B(new_n663), .C1(new_n668), .C2(new_n730), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n663), .B2(new_n730), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT108), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(new_n739), .A3(KEYINPUT45), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT45), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n1032), .B2(new_n738), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(KEYINPUT44), .B1(new_n1033), .B2(new_n739), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT44), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1032), .A2(new_n1039), .A3(new_n738), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n727), .A2(new_n735), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1037), .A2(new_n736), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1029), .A2(new_n1043), .A3(new_n781), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n781), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n742), .B(KEYINPUT41), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1025), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1023), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT106), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1052), .A2(KEYINPUT43), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n735), .A2(new_n737), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1033), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT42), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT42), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1033), .A2(new_n1059), .A3(new_n1056), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n707), .B1(new_n1033), .B2(new_n733), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1058), .B(new_n1060), .C1(new_n720), .C2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(KEYINPUT107), .B1(new_n736), .B2(new_n1032), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1023), .A2(KEYINPUT43), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT107), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1042), .A2(new_n1065), .A3(new_n1033), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1064), .A2(new_n1062), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1055), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n1054), .A3(new_n1067), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1024), .B1(new_n1048), .B2(new_n1075), .ZN(G387));
  NAND2_X1  g0876(.A1(new_n1029), .A2(new_n1025), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n817), .A2(G317), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n838), .A2(G322), .B1(G311), .B2(new_n847), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n814), .C2(new_n505), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT48), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n830), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n888), .A2(G283), .B1(G294), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT49), .Z(new_n1087));
  AOI21_X1  g0887(.A(new_n280), .B1(new_n823), .B2(G326), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n247), .B2(new_n836), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n814), .A2(new_n270), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n817), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n227), .A2(new_n1092), .B1(new_n881), .B2(new_n882), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n888), .A2(new_n322), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1084), .A2(new_n323), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1094), .A2(new_n1010), .A3(new_n280), .A4(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n448), .A2(new_n834), .B1(new_n370), .B2(new_n822), .ZN(new_n1097));
  NOR4_X1   g0897(.A1(new_n1091), .A2(new_n1093), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n793), .B1(new_n1090), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n735), .A2(new_n792), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n797), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n239), .B2(new_n798), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n744), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n801), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n327), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n227), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT50), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n344), .B1(new_n270), .B2(new_n273), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1107), .A2(new_n1103), .A3(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1104), .A2(new_n1109), .B1(G107), .B2(new_n209), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n786), .B1(new_n1110), .B2(new_n794), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1099), .A2(new_n1100), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1029), .A2(new_n781), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n742), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1029), .A2(new_n781), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1077), .B(new_n1112), .C1(new_n1114), .C2(new_n1115), .ZN(G393));
  NAND3_X1  g0916(.A1(new_n1043), .A2(KEYINPUT111), .A3(new_n1044), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT111), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1041), .A2(new_n1118), .A3(new_n1042), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1117), .A2(new_n1113), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1045), .A2(new_n742), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT114), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1117), .A2(new_n1113), .A3(new_n1119), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT114), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n742), .A4(new_n1045), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1032), .A2(new_n792), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n248), .A2(new_n1101), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n794), .B1(new_n204), .B2(new_n209), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n807), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n834), .A2(new_n227), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n888), .A2(G77), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n382), .B1(new_n1084), .B2(G68), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(new_n536), .C2(new_n836), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1131), .B(new_n1134), .C1(G143), .C2(new_n823), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G150), .A2(new_n838), .B1(new_n817), .B2(G159), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1135), .B(new_n1138), .C1(new_n327), .C2(new_n814), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n823), .A2(G322), .B1(G283), .B2(new_n1084), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT113), .Z(new_n1142));
  NOR2_X1   g0942(.A1(new_n834), .A2(new_n505), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n382), .B1(new_n827), .B2(new_n247), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G107), .C2(new_n835), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1142), .B(new_n1145), .C1(new_n844), .C2(new_n814), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G311), .A2(new_n817), .B1(new_n838), .B2(G317), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT52), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1139), .A2(new_n1140), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1130), .B1(new_n793), .B2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1126), .A2(new_n1025), .B1(new_n1127), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1122), .A2(new_n1125), .A3(new_n1151), .ZN(G390));
  INV_X1    g0952(.A(G330), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n862), .B2(new_n864), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n981), .B2(new_n986), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n939), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n975), .A2(new_n713), .A3(new_n865), .A4(new_n939), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n720), .B1(new_n775), .B2(new_n778), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n933), .B1(new_n1160), .B2(new_n865), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n713), .B(new_n865), .C1(new_n981), .C2(new_n986), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1156), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n975), .A2(new_n939), .A3(new_n1154), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1159), .A2(new_n1161), .B1(new_n1165), .B2(new_n935), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT115), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n991), .B2(G330), .ZN(new_n1168));
  AND4_X1   g0968(.A1(new_n1167), .A2(new_n685), .A3(new_n975), .A4(G330), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n684), .B(new_n972), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n944), .B(new_n980), .C1(new_n1161), .C2(new_n1156), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n945), .B1(new_n935), .B2(new_n939), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1158), .C1(new_n970), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n933), .B1(new_n861), .B2(new_n361), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n944), .B1(new_n1177), .B2(new_n1156), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n963), .A2(new_n965), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n968), .B1(new_n1179), .B2(KEYINPUT104), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1180), .A3(new_n967), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1164), .B1(new_n1181), .B2(new_n1173), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1172), .B1(new_n1176), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1173), .B1(new_n970), .B2(new_n1174), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1164), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(new_n1171), .A3(new_n1175), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1183), .A2(new_n742), .A3(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1176), .A2(new_n1182), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n970), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n790), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n807), .B1(new_n376), .B2(new_n871), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n838), .A2(G283), .B1(G107), .B2(new_n847), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n814), .B2(new_n204), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT118), .Z(new_n1195));
  AOI21_X1  g0995(.A(new_n280), .B1(new_n1084), .B2(G87), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n886), .A2(new_n1132), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G294), .B2(new_n823), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1195), .B(new_n1198), .C1(new_n247), .C2(new_n1092), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(KEYINPUT54), .B(G143), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n815), .A2(new_n1201), .B1(G137), .B2(new_n847), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1202), .A2(KEYINPUT116), .B1(G159), .B2(new_n888), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(KEYINPUT116), .B2(new_n1202), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT117), .Z(new_n1205));
  AOI22_X1  g1005(.A1(G128), .A2(new_n838), .B1(new_n817), .B2(G132), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1084), .A2(G150), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(KEYINPUT53), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n382), .B1(new_n1207), .B2(KEYINPUT53), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G125), .A2(new_n823), .B1(new_n835), .B2(G50), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1206), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1199), .B1(new_n1205), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1192), .B1(new_n1212), .B2(new_n793), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1189), .A2(new_n1025), .B1(new_n1191), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1188), .A2(new_n1214), .ZN(G378));
  INV_X1    g1015(.A(KEYINPUT57), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1166), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1170), .B1(new_n1189), .B2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(G330), .B(new_n989), .C1(new_n978), .C2(KEYINPUT40), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n405), .B(KEYINPUT121), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n911), .A2(new_n378), .ZN(new_n1221));
  XOR2_X1   g1021(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1222));
  XNOR2_X1  g1022(.A(new_n1221), .B(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1220), .B(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1219), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1219), .A2(new_n1224), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1190), .A2(new_n944), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n1225), .A2(new_n1226), .B1(new_n1227), .B2(new_n942), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1224), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n979), .A2(new_n1229), .A3(G330), .A4(new_n989), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1219), .A2(new_n1224), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n971), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1228), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1216), .B1(new_n1218), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1170), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1187), .A2(new_n1235), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1236), .A2(KEYINPUT57), .A3(new_n1232), .A4(new_n1228), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(new_n742), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1228), .A2(new_n1232), .A3(new_n1025), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G97), .A2(new_n847), .B1(new_n835), .B2(G58), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1095), .A2(new_n291), .A3(new_n382), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1240), .B1(new_n1013), .B2(new_n822), .C1(KEYINPUT119), .C2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1002), .B1(new_n1241), .B2(KEYINPUT119), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1243), .B1(new_n1092), .B2(new_n205), .C1(new_n247), .C2(new_n881), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1242), .B(new_n1244), .C1(new_n322), .C2(new_n815), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1245), .A2(KEYINPUT58), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n834), .A2(new_n890), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n827), .A2(new_n370), .B1(new_n830), .B2(new_n1200), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n838), .C2(G125), .ZN(new_n1249));
  INV_X1    g1049(.A(G128), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1092), .C1(new_n880), .C2(new_n814), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1251), .A2(KEYINPUT59), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(KEYINPUT59), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n319), .B(new_n291), .C1(new_n836), .C2(new_n882), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G124), .B2(new_n823), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1245), .A2(KEYINPUT58), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n291), .B1(new_n380), .B2(new_n319), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n227), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1246), .A2(new_n1256), .A3(new_n1257), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n793), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT120), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n786), .B1(new_n227), .B2(new_n870), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(new_n791), .C2(new_n1224), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1239), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1238), .A2(new_n1266), .ZN(G375));
  NAND2_X1  g1067(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1172), .A2(new_n1047), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1156), .A2(new_n790), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(KEYINPUT122), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n888), .A2(new_n322), .B1(G97), .B2(new_n1084), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n1272), .B1(new_n247), .B2(new_n834), .C1(new_n505), .C2(new_n822), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n1013), .A2(new_n1092), .B1(new_n881), .B2(new_n844), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1273), .B(new_n1274), .C1(G107), .C2(new_n815), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n280), .B1(new_n835), .B2(G77), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n1276), .B(KEYINPUT123), .Z(new_n1277));
  NAND2_X1  g1077(.A1(new_n815), .A2(G150), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n890), .A2(new_n881), .B1(new_n1092), .B2(new_n880), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n382), .B1(new_n1084), .B2(G159), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1280), .B1(new_n227), .B2(new_n827), .C1(new_n836), .C2(new_n373), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n1250), .A2(new_n822), .B1(new_n834), .B2(new_n1200), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1279), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n1275), .A2(new_n1277), .B1(new_n1278), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n793), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n807), .B1(G68), .B2(new_n871), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1271), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1217), .B2(new_n1025), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1269), .A2(new_n1288), .ZN(G381));
  AND2_X1   g1089(.A1(new_n1238), .A2(new_n1266), .ZN(new_n1290));
  INV_X1    g1090(.A(G378), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(G390), .A2(G387), .ZN(new_n1292));
  NOR4_X1   g1092(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .A4(new_n1293), .ZN(G407));
  NAND4_X1  g1094(.A1(new_n1290), .A2(G213), .A3(new_n719), .A4(new_n1291), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(G407), .A2(new_n1295), .A3(G213), .ZN(G409));
  NAND2_X1  g1096(.A1(new_n719), .A2(G213), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1165), .A2(new_n935), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1170), .A2(KEYINPUT60), .A3(new_n1298), .A4(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1300), .A2(new_n742), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT60), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1268), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1301), .A2(new_n1302), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1302), .B1(new_n1301), .B2(new_n1304), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1288), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n895), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G384), .B(new_n1288), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1238), .A2(G378), .A3(new_n1266), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1236), .A2(new_n1047), .A3(new_n1232), .A4(new_n1228), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1265), .B1(new_n1312), .B2(KEYINPUT124), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1233), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT124), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1314), .A2(new_n1315), .A3(new_n1047), .A4(new_n1236), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G378), .B1(new_n1313), .B2(new_n1316), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1297), .B(new_n1310), .C1(new_n1311), .C2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(KEYINPUT62), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1297), .B1(new_n1311), .B2(new_n1317), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n719), .A2(G213), .A3(G2897), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1308), .A2(new_n1309), .A3(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1321), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1320), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1312), .A2(KEYINPUT124), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1326), .A2(new_n1316), .A3(new_n1266), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1291), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1238), .A2(G378), .A3(new_n1266), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT62), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1330), .A2(new_n1331), .A3(new_n1297), .A4(new_n1310), .ZN(new_n1332));
  XOR2_X1   g1132(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1333));
  NAND4_X1  g1133(.A1(new_n1319), .A2(new_n1325), .A3(new_n1332), .A4(new_n1333), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(G393), .B(new_n857), .ZN(new_n1335));
  AND2_X1   g1135(.A1(G390), .A2(G387), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1335), .B1(new_n1336), .B2(new_n1292), .ZN(new_n1337));
  OR2_X1    g1137(.A1(G390), .A2(G387), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1335), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(G390), .A2(G387), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1338), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1337), .A2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1334), .A2(new_n1342), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1342), .A2(KEYINPUT61), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT63), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1318), .A2(new_n1345), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1330), .A2(KEYINPUT63), .A3(new_n1297), .A4(new_n1310), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1344), .A2(new_n1346), .A3(new_n1325), .A4(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1343), .A2(new_n1348), .ZN(G405));
  NAND2_X1  g1149(.A1(new_n1329), .A2(KEYINPUT127), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1310), .A2(new_n1291), .A3(G375), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1352), .B1(new_n1290), .B2(G378), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1342), .A2(new_n1351), .A3(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1342), .B1(new_n1351), .B2(new_n1353), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1350), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1353), .A2(new_n1351), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1358), .A2(new_n1337), .A3(new_n1341), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1359), .A2(KEYINPUT127), .A3(new_n1329), .A4(new_n1354), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1357), .A2(new_n1360), .ZN(G402));
endmodule


