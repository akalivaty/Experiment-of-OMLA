

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(G651), .A2(n625), .ZN(n645) );
  NOR2_X1 U553 ( .A1(n673), .A2(G1384), .ZN(n788) );
  INV_X2 U554 ( .A(G2105), .ZN(n519) );
  AND2_X2 U555 ( .A1(n519), .A2(G2104), .ZN(n896) );
  NOR2_X2 U556 ( .A1(G2104), .A2(n519), .ZN(n891) );
  INV_X1 U557 ( .A(n911), .ZN(n976) );
  OR2_X1 U558 ( .A1(n687), .A2(n976), .ZN(n686) );
  XNOR2_X1 U559 ( .A(n680), .B(n679), .ZN(n687) );
  INV_X1 U560 ( .A(KEYINPUT95), .ZN(n679) );
  XNOR2_X1 U561 ( .A(n520), .B(KEYINPUT17), .ZN(n556) );
  INV_X1 U562 ( .A(KEYINPUT92), .ZN(n676) );
  XNOR2_X1 U563 ( .A(n725), .B(n676), .ZN(n691) );
  BUF_X1 U564 ( .A(n691), .Z(n704) );
  INV_X1 U565 ( .A(KEYINPUT30), .ZN(n714) );
  XNOR2_X1 U566 ( .A(n714), .B(KEYINPUT97), .ZN(n715) );
  XNOR2_X1 U567 ( .A(n716), .B(n715), .ZN(n717) );
  INV_X1 U568 ( .A(KEYINPUT29), .ZN(n701) );
  INV_X1 U569 ( .A(KEYINPUT31), .ZN(n721) );
  INV_X1 U570 ( .A(KEYINPUT91), .ZN(n711) );
  XNOR2_X1 U571 ( .A(n712), .B(n711), .ZN(n739) );
  INV_X1 U572 ( .A(KEYINPUT101), .ZN(n747) );
  XNOR2_X1 U573 ( .A(n748), .B(n747), .ZN(n749) );
  INV_X1 U574 ( .A(G2104), .ZN(n518) );
  NAND2_X1 U575 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U576 ( .A(KEYINPUT14), .B(KEYINPUT68), .ZN(n585) );
  XNOR2_X1 U577 ( .A(n586), .B(n585), .ZN(n587) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n642) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n530), .Z(n640) );
  BUF_X1 U580 ( .A(n674), .Z(G160) );
  INV_X1 U581 ( .A(n556), .ZN(n521) );
  INV_X2 U582 ( .A(n521), .ZN(n895) );
  NAND2_X1 U583 ( .A1(n895), .A2(G137), .ZN(n524) );
  NAND2_X1 U584 ( .A1(G101), .A2(n896), .ZN(n522) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n522), .Z(n523) );
  NAND2_X1 U586 ( .A1(n524), .A2(n523), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n891), .A2(G125), .ZN(n527) );
  NAND2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XOR2_X2 U589 ( .A(KEYINPUT64), .B(n525), .Z(n892) );
  NAND2_X1 U590 ( .A1(G113), .A2(n892), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n674) );
  INV_X1 U593 ( .A(G651), .ZN(n537) );
  NOR2_X1 U594 ( .A1(G543), .A2(n537), .ZN(n530) );
  NAND2_X1 U595 ( .A1(G63), .A2(n640), .ZN(n532) );
  XOR2_X1 U596 ( .A(KEYINPUT0), .B(G543), .Z(n625) );
  NAND2_X1 U597 ( .A1(G51), .A2(n645), .ZN(n531) );
  NAND2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n534) );
  XOR2_X1 U599 ( .A(KEYINPUT6), .B(KEYINPUT71), .Z(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n542) );
  NAND2_X1 U601 ( .A1(G89), .A2(n642), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n535), .B(KEYINPUT70), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT4), .ZN(n539) );
  NOR2_X1 U604 ( .A1(n625), .A2(n537), .ZN(n641) );
  NAND2_X1 U605 ( .A1(G76), .A2(n641), .ZN(n538) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U607 ( .A(KEYINPUT5), .B(n540), .Z(n541) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n544) );
  XOR2_X1 U609 ( .A(KEYINPUT7), .B(KEYINPUT72), .Z(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G168) );
  XOR2_X1 U611 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U613 ( .A1(G99), .A2(n896), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n545), .B(KEYINPUT76), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G123), .A2(n891), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n546), .B(KEYINPUT74), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n547), .B(KEYINPUT18), .ZN(n549) );
  NAND2_X1 U618 ( .A1(G135), .A2(n895), .ZN(n548) );
  NAND2_X1 U619 ( .A1(n549), .A2(n548), .ZN(n552) );
  NAND2_X1 U620 ( .A1(G111), .A2(n892), .ZN(n550) );
  XNOR2_X1 U621 ( .A(KEYINPUT75), .B(n550), .ZN(n551) );
  NOR2_X1 U622 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U623 ( .A1(n554), .A2(n553), .ZN(n1005) );
  XNOR2_X1 U624 ( .A(G2096), .B(n1005), .ZN(n555) );
  OR2_X1 U625 ( .A1(G2100), .A2(n555), .ZN(G156) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G132), .ZN(G219) );
  INV_X1 U628 ( .A(G82), .ZN(G220) );
  NAND2_X1 U629 ( .A1(n896), .A2(G102), .ZN(n559) );
  NAND2_X1 U630 ( .A1(n556), .A2(G138), .ZN(n557) );
  XOR2_X1 U631 ( .A(n557), .B(KEYINPUT83), .Z(n558) );
  NAND2_X1 U632 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n891), .A2(G126), .ZN(n561) );
  NAND2_X1 U634 ( .A1(G114), .A2(n892), .ZN(n560) );
  NAND2_X1 U635 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U636 ( .A1(n563), .A2(n562), .ZN(n673) );
  BUF_X1 U637 ( .A(n673), .Z(G164) );
  NAND2_X1 U638 ( .A1(G64), .A2(n640), .ZN(n565) );
  NAND2_X1 U639 ( .A1(G52), .A2(n645), .ZN(n564) );
  NAND2_X1 U640 ( .A1(n565), .A2(n564), .ZN(n571) );
  NAND2_X1 U641 ( .A1(G77), .A2(n641), .ZN(n567) );
  NAND2_X1 U642 ( .A1(G90), .A2(n642), .ZN(n566) );
  NAND2_X1 U643 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U644 ( .A(KEYINPUT66), .B(n568), .Z(n569) );
  XNOR2_X1 U645 ( .A(KEYINPUT9), .B(n569), .ZN(n570) );
  NOR2_X1 U646 ( .A1(n571), .A2(n570), .ZN(G171) );
  NAND2_X1 U647 ( .A1(G62), .A2(n640), .ZN(n573) );
  NAND2_X1 U648 ( .A1(G50), .A2(n645), .ZN(n572) );
  NAND2_X1 U649 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U650 ( .A(KEYINPUT81), .B(n574), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n641), .A2(G75), .ZN(n576) );
  NAND2_X1 U652 ( .A1(G88), .A2(n642), .ZN(n575) );
  AND2_X1 U653 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(G303) );
  NAND2_X1 U655 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U656 ( .A(n579), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U657 ( .A(G223), .ZN(n828) );
  NAND2_X1 U658 ( .A1(n828), .A2(G567), .ZN(n580) );
  XOR2_X1 U659 ( .A(KEYINPUT11), .B(n580), .Z(G234) );
  NAND2_X1 U660 ( .A1(n642), .A2(G81), .ZN(n581) );
  XNOR2_X1 U661 ( .A(n581), .B(KEYINPUT12), .ZN(n583) );
  NAND2_X1 U662 ( .A1(G68), .A2(n641), .ZN(n582) );
  NAND2_X1 U663 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U664 ( .A(n584), .B(KEYINPUT13), .ZN(n588) );
  NAND2_X1 U665 ( .A1(G56), .A2(n640), .ZN(n586) );
  NAND2_X1 U666 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U667 ( .A(n589), .B(KEYINPUT69), .ZN(n591) );
  NAND2_X1 U668 ( .A1(G43), .A2(n645), .ZN(n590) );
  NAND2_X1 U669 ( .A1(n591), .A2(n590), .ZN(n991) );
  INV_X1 U670 ( .A(G860), .ZN(n610) );
  OR2_X1 U671 ( .A1(n991), .A2(n610), .ZN(G153) );
  INV_X1 U672 ( .A(G171), .ZN(G301) );
  NAND2_X1 U673 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U674 ( .A1(G79), .A2(n641), .ZN(n593) );
  NAND2_X1 U675 ( .A1(G92), .A2(n642), .ZN(n592) );
  NAND2_X1 U676 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U677 ( .A1(G66), .A2(n640), .ZN(n595) );
  NAND2_X1 U678 ( .A1(G54), .A2(n645), .ZN(n594) );
  NAND2_X1 U679 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U680 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U681 ( .A(KEYINPUT15), .B(n598), .Z(n911) );
  INV_X1 U682 ( .A(G868), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n976), .A2(n613), .ZN(n599) );
  NAND2_X1 U684 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U685 ( .A1(G78), .A2(n641), .ZN(n602) );
  NAND2_X1 U686 ( .A1(G91), .A2(n642), .ZN(n601) );
  NAND2_X1 U687 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U688 ( .A1(G65), .A2(n640), .ZN(n603) );
  XNOR2_X1 U689 ( .A(KEYINPUT67), .B(n603), .ZN(n604) );
  NOR2_X1 U690 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U691 ( .A1(n645), .A2(G53), .ZN(n606) );
  NAND2_X1 U692 ( .A1(n607), .A2(n606), .ZN(G299) );
  NAND2_X1 U693 ( .A1(G868), .A2(G286), .ZN(n609) );
  NAND2_X1 U694 ( .A1(G299), .A2(n613), .ZN(n608) );
  NAND2_X1 U695 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U696 ( .A1(n610), .A2(G559), .ZN(n611) );
  NAND2_X1 U697 ( .A1(n611), .A2(n911), .ZN(n612) );
  XNOR2_X1 U698 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U699 ( .A1(n976), .A2(n613), .ZN(n614) );
  XNOR2_X1 U700 ( .A(n614), .B(KEYINPUT73), .ZN(n615) );
  NOR2_X1 U701 ( .A1(G559), .A2(n615), .ZN(n617) );
  NOR2_X1 U702 ( .A1(G868), .A2(n991), .ZN(n616) );
  NOR2_X1 U703 ( .A1(n617), .A2(n616), .ZN(G282) );
  INV_X1 U704 ( .A(G303), .ZN(G166) );
  NAND2_X1 U705 ( .A1(G86), .A2(n642), .ZN(n619) );
  NAND2_X1 U706 ( .A1(G61), .A2(n640), .ZN(n618) );
  NAND2_X1 U707 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U708 ( .A1(n641), .A2(G73), .ZN(n620) );
  XOR2_X1 U709 ( .A(KEYINPUT2), .B(n620), .Z(n621) );
  NOR2_X1 U710 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U711 ( .A1(n645), .A2(G48), .ZN(n623) );
  NAND2_X1 U712 ( .A1(n624), .A2(n623), .ZN(G305) );
  NAND2_X1 U713 ( .A1(G87), .A2(n625), .ZN(n626) );
  XNOR2_X1 U714 ( .A(n626), .B(KEYINPUT80), .ZN(n631) );
  NAND2_X1 U715 ( .A1(G49), .A2(n645), .ZN(n628) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U717 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U718 ( .A1(n640), .A2(n629), .ZN(n630) );
  NAND2_X1 U719 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U720 ( .A1(G60), .A2(n640), .ZN(n633) );
  NAND2_X1 U721 ( .A1(G47), .A2(n645), .ZN(n632) );
  NAND2_X1 U722 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U723 ( .A1(G72), .A2(n641), .ZN(n634) );
  XNOR2_X1 U724 ( .A(KEYINPUT65), .B(n634), .ZN(n635) );
  NOR2_X1 U725 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U726 ( .A1(n642), .A2(G85), .ZN(n637) );
  NAND2_X1 U727 ( .A1(n638), .A2(n637), .ZN(G290) );
  NAND2_X1 U728 ( .A1(G559), .A2(n911), .ZN(n639) );
  XNOR2_X1 U729 ( .A(n639), .B(n991), .ZN(n836) );
  NAND2_X1 U730 ( .A1(G67), .A2(n640), .ZN(n650) );
  NAND2_X1 U731 ( .A1(G80), .A2(n641), .ZN(n644) );
  NAND2_X1 U732 ( .A1(G93), .A2(n642), .ZN(n643) );
  NAND2_X1 U733 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U734 ( .A1(n645), .A2(G55), .ZN(n646) );
  XOR2_X1 U735 ( .A(KEYINPUT78), .B(n646), .Z(n647) );
  NOR2_X1 U736 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U737 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U738 ( .A(n651), .B(KEYINPUT79), .ZN(n839) );
  XNOR2_X1 U739 ( .A(G166), .B(n839), .ZN(n657) );
  XNOR2_X1 U740 ( .A(KEYINPUT82), .B(G305), .ZN(n652) );
  XNOR2_X1 U741 ( .A(n652), .B(G288), .ZN(n653) );
  XNOR2_X1 U742 ( .A(KEYINPUT19), .B(n653), .ZN(n655) );
  INV_X1 U743 ( .A(G299), .ZN(n979) );
  XNOR2_X1 U744 ( .A(G290), .B(n979), .ZN(n654) );
  XNOR2_X1 U745 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U746 ( .A(n657), .B(n656), .ZN(n914) );
  XNOR2_X1 U747 ( .A(n836), .B(n914), .ZN(n658) );
  NAND2_X1 U748 ( .A1(n658), .A2(G868), .ZN(n660) );
  OR2_X1 U749 ( .A1(G868), .A2(n839), .ZN(n659) );
  NAND2_X1 U750 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2078), .A2(G2084), .ZN(n661) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U755 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n665) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n665), .Z(n666) );
  NOR2_X1 U759 ( .A1(G218), .A2(n666), .ZN(n667) );
  NAND2_X1 U760 ( .A1(G96), .A2(n667), .ZN(n834) );
  NAND2_X1 U761 ( .A1(n834), .A2(G2106), .ZN(n671) );
  NAND2_X1 U762 ( .A1(G120), .A2(G69), .ZN(n668) );
  NOR2_X1 U763 ( .A1(G237), .A2(n668), .ZN(n669) );
  NAND2_X1 U764 ( .A1(G108), .A2(n669), .ZN(n835) );
  NAND2_X1 U765 ( .A1(n835), .A2(G567), .ZN(n670) );
  NAND2_X1 U766 ( .A1(n671), .A2(n670), .ZN(n924) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U768 ( .A1(n924), .A2(n672), .ZN(n833) );
  NAND2_X1 U769 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U770 ( .A1(n674), .A2(G40), .ZN(n787) );
  INV_X1 U771 ( .A(n787), .ZN(n675) );
  NAND2_X2 U772 ( .A1(n788), .A2(n675), .ZN(n725) );
  NAND2_X1 U773 ( .A1(G8), .A2(n725), .ZN(n817) );
  NAND2_X1 U774 ( .A1(n691), .A2(G2067), .ZN(n678) );
  NAND2_X1 U775 ( .A1(G1348), .A2(n725), .ZN(n677) );
  NAND2_X1 U776 ( .A1(n678), .A2(n677), .ZN(n680) );
  INV_X1 U777 ( .A(n725), .ZN(n703) );
  NAND2_X1 U778 ( .A1(G1996), .A2(n703), .ZN(n681) );
  XOR2_X1 U779 ( .A(KEYINPUT26), .B(n681), .Z(n682) );
  NOR2_X1 U780 ( .A1(n991), .A2(n682), .ZN(n684) );
  NAND2_X1 U781 ( .A1(G1341), .A2(n725), .ZN(n683) );
  NAND2_X1 U782 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U783 ( .A1(n686), .A2(n685), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n976), .A2(n687), .ZN(n688) );
  NAND2_X1 U785 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U786 ( .A(n690), .B(KEYINPUT96), .ZN(n696) );
  NAND2_X1 U787 ( .A1(G2072), .A2(n704), .ZN(n692) );
  XNOR2_X1 U788 ( .A(n692), .B(KEYINPUT27), .ZN(n694) );
  XOR2_X1 U789 ( .A(G1956), .B(KEYINPUT94), .Z(n930) );
  NOR2_X1 U790 ( .A1(n704), .A2(n930), .ZN(n693) );
  NOR2_X1 U791 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U792 ( .A1(n697), .A2(n979), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n696), .A2(n695), .ZN(n700) );
  NOR2_X1 U794 ( .A1(n697), .A2(n979), .ZN(n698) );
  XOR2_X1 U795 ( .A(n698), .B(KEYINPUT28), .Z(n699) );
  NAND2_X1 U796 ( .A1(n700), .A2(n699), .ZN(n702) );
  XNOR2_X1 U797 ( .A(n702), .B(n701), .ZN(n710) );
  NOR2_X1 U798 ( .A1(n703), .A2(G1961), .ZN(n707) );
  XOR2_X1 U799 ( .A(G2078), .B(KEYINPUT25), .Z(n959) );
  INV_X1 U800 ( .A(n704), .ZN(n705) );
  NOR2_X1 U801 ( .A1(n959), .A2(n705), .ZN(n706) );
  NOR2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U803 ( .A(n708), .B(KEYINPUT93), .ZN(n718) );
  NAND2_X1 U804 ( .A1(n718), .A2(G171), .ZN(n709) );
  NAND2_X1 U805 ( .A1(n710), .A2(n709), .ZN(n724) );
  NOR2_X1 U806 ( .A1(G1966), .A2(n817), .ZN(n712) );
  NOR2_X1 U807 ( .A1(G2084), .A2(n725), .ZN(n735) );
  NOR2_X1 U808 ( .A1(n739), .A2(n735), .ZN(n713) );
  NAND2_X1 U809 ( .A1(G8), .A2(n713), .ZN(n716) );
  NOR2_X1 U810 ( .A1(n717), .A2(G168), .ZN(n720) );
  NOR2_X1 U811 ( .A1(G171), .A2(n718), .ZN(n719) );
  NOR2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n722) );
  XNOR2_X1 U813 ( .A(n722), .B(n721), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n737) );
  NAND2_X1 U815 ( .A1(n737), .A2(G286), .ZN(n730) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n817), .ZN(n727) );
  NOR2_X1 U817 ( .A1(G2090), .A2(n725), .ZN(n726) );
  NOR2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U819 ( .A1(n728), .A2(G303), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U821 ( .A(n731), .B(KEYINPUT98), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n732), .A2(G8), .ZN(n734) );
  XOR2_X1 U823 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n733) );
  XNOR2_X1 U824 ( .A(n734), .B(n733), .ZN(n743) );
  NAND2_X1 U825 ( .A1(G8), .A2(n735), .ZN(n736) );
  XNOR2_X1 U826 ( .A(KEYINPUT90), .B(n736), .ZN(n741) );
  INV_X1 U827 ( .A(n737), .ZN(n738) );
  NOR2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n811) );
  NOR2_X1 U831 ( .A1(G1971), .A2(G303), .ZN(n744) );
  XNOR2_X1 U832 ( .A(n744), .B(KEYINPUT100), .ZN(n745) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n983) );
  NOR2_X1 U834 ( .A1(n745), .A2(n983), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n811), .A2(n746), .ZN(n748) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n980) );
  NAND2_X1 U837 ( .A1(n749), .A2(n980), .ZN(n750) );
  XNOR2_X1 U838 ( .A(n750), .B(KEYINPUT102), .ZN(n751) );
  NOR2_X1 U839 ( .A1(n817), .A2(n751), .ZN(n752) );
  NOR2_X1 U840 ( .A1(KEYINPUT33), .A2(n752), .ZN(n753) );
  XNOR2_X1 U841 ( .A(n753), .B(KEYINPUT103), .ZN(n810) );
  NAND2_X1 U842 ( .A1(n983), .A2(KEYINPUT33), .ZN(n754) );
  NOR2_X1 U843 ( .A1(n754), .A2(n817), .ZN(n755) );
  XOR2_X1 U844 ( .A(n755), .B(KEYINPUT104), .Z(n756) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n973) );
  AND2_X1 U846 ( .A1(n756), .A2(n973), .ZN(n808) );
  NAND2_X1 U847 ( .A1(n895), .A2(G140), .ZN(n757) );
  XOR2_X1 U848 ( .A(KEYINPUT85), .B(n757), .Z(n759) );
  NAND2_X1 U849 ( .A1(n896), .A2(G104), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U851 ( .A(KEYINPUT34), .B(n760), .ZN(n766) );
  NAND2_X1 U852 ( .A1(G116), .A2(n892), .ZN(n761) );
  XNOR2_X1 U853 ( .A(n761), .B(KEYINPUT86), .ZN(n763) );
  NAND2_X1 U854 ( .A1(G128), .A2(n891), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U856 ( .A(KEYINPUT35), .B(n764), .Z(n765) );
  NOR2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U858 ( .A(n767), .B(KEYINPUT36), .ZN(n768) );
  XOR2_X1 U859 ( .A(n768), .B(KEYINPUT87), .Z(n907) );
  XNOR2_X1 U860 ( .A(G2067), .B(KEYINPUT37), .ZN(n796) );
  AND2_X1 U861 ( .A1(n907), .A2(n796), .ZN(n769) );
  XNOR2_X1 U862 ( .A(KEYINPUT107), .B(n769), .ZN(n1012) );
  NAND2_X1 U863 ( .A1(G141), .A2(n895), .ZN(n771) );
  NAND2_X1 U864 ( .A1(G129), .A2(n891), .ZN(n770) );
  NAND2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n896), .A2(G105), .ZN(n772) );
  XOR2_X1 U867 ( .A(KEYINPUT38), .B(n772), .Z(n773) );
  NOR2_X1 U868 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U869 ( .A1(G117), .A2(n892), .ZN(n775) );
  NAND2_X1 U870 ( .A1(n776), .A2(n775), .ZN(n877) );
  NOR2_X1 U871 ( .A1(G1996), .A2(n877), .ZN(n999) );
  NAND2_X1 U872 ( .A1(G131), .A2(n895), .ZN(n778) );
  NAND2_X1 U873 ( .A1(G95), .A2(n896), .ZN(n777) );
  NAND2_X1 U874 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U875 ( .A(KEYINPUT88), .B(n779), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n891), .A2(G119), .ZN(n781) );
  NAND2_X1 U877 ( .A1(G107), .A2(n892), .ZN(n780) );
  NAND2_X1 U878 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U880 ( .A(KEYINPUT89), .B(n784), .ZN(n906) );
  AND2_X1 U881 ( .A1(n906), .A2(G1991), .ZN(n786) );
  AND2_X1 U882 ( .A1(n877), .A2(G1996), .ZN(n785) );
  NOR2_X1 U883 ( .A1(n786), .A2(n785), .ZN(n1002) );
  NOR2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n801) );
  INV_X1 U885 ( .A(n801), .ZN(n789) );
  NOR2_X1 U886 ( .A1(n1002), .A2(n789), .ZN(n802) );
  NOR2_X1 U887 ( .A1(G1986), .A2(G290), .ZN(n790) );
  NOR2_X1 U888 ( .A1(G1991), .A2(n906), .ZN(n1004) );
  NOR2_X1 U889 ( .A1(n790), .A2(n1004), .ZN(n791) );
  NOR2_X1 U890 ( .A1(n802), .A2(n791), .ZN(n792) );
  XOR2_X1 U891 ( .A(KEYINPUT105), .B(n792), .Z(n793) );
  NOR2_X1 U892 ( .A1(n999), .A2(n793), .ZN(n794) );
  XNOR2_X1 U893 ( .A(KEYINPUT39), .B(n794), .ZN(n795) );
  XNOR2_X1 U894 ( .A(n795), .B(KEYINPUT106), .ZN(n797) );
  NOR2_X1 U895 ( .A1(n907), .A2(n796), .ZN(n1007) );
  NAND2_X1 U896 ( .A1(n801), .A2(n1007), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n797), .A2(n804), .ZN(n798) );
  NAND2_X1 U898 ( .A1(n1012), .A2(n798), .ZN(n799) );
  NAND2_X1 U899 ( .A1(n799), .A2(n801), .ZN(n820) );
  XNOR2_X1 U900 ( .A(G1986), .B(KEYINPUT84), .ZN(n800) );
  XNOR2_X1 U901 ( .A(n800), .B(G290), .ZN(n987) );
  AND2_X1 U902 ( .A1(n987), .A2(n801), .ZN(n806) );
  INV_X1 U903 ( .A(n802), .ZN(n803) );
  NAND2_X1 U904 ( .A1(n804), .A2(n803), .ZN(n805) );
  OR2_X1 U905 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U906 ( .A1(n820), .A2(n807), .ZN(n824) );
  AND2_X1 U907 ( .A1(n808), .A2(n824), .ZN(n809) );
  NAND2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n826) );
  NOR2_X1 U909 ( .A1(G2090), .A2(G303), .ZN(n812) );
  NAND2_X1 U910 ( .A1(G8), .A2(n812), .ZN(n813) );
  NAND2_X1 U911 ( .A1(n811), .A2(n813), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n814), .A2(n817), .ZN(n819) );
  NOR2_X1 U913 ( .A1(G1981), .A2(G305), .ZN(n815) );
  XOR2_X1 U914 ( .A(n815), .B(KEYINPUT24), .Z(n816) );
  OR2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n822) );
  INV_X1 U917 ( .A(n820), .ZN(n821) );
  OR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U921 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n828), .ZN(G217) );
  INV_X1 U923 ( .A(G661), .ZN(n830) );
  NAND2_X1 U924 ( .A1(G2), .A2(G15), .ZN(n829) );
  NOR2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  XOR2_X1 U926 ( .A(KEYINPUT112), .B(n831), .Z(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U929 ( .A(G69), .B(KEYINPUT113), .ZN(G235) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  NOR2_X1 U935 ( .A1(G860), .A2(n836), .ZN(n837) );
  XOR2_X1 U936 ( .A(KEYINPUT77), .B(n837), .Z(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(G145) );
  XNOR2_X1 U938 ( .A(G1348), .B(G1341), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n840), .B(G2427), .ZN(n850) );
  XOR2_X1 U940 ( .A(G2446), .B(KEYINPUT109), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2430), .B(G2451), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U943 ( .A(KEYINPUT110), .B(G2438), .Z(n844) );
  XNOR2_X1 U944 ( .A(G2435), .B(G2454), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U946 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U947 ( .A(KEYINPUT108), .B(G2443), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  NAND2_X1 U950 ( .A1(n851), .A2(G14), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n852), .B(KEYINPUT111), .ZN(G401) );
  XOR2_X1 U952 ( .A(G2100), .B(G2096), .Z(n854) );
  XNOR2_X1 U953 ( .A(KEYINPUT42), .B(G2678), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U955 ( .A(KEYINPUT43), .B(G2090), .Z(n856) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U958 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U959 ( .A(G2078), .B(G2084), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U961 ( .A(G1976), .B(G1981), .Z(n862) );
  XNOR2_X1 U962 ( .A(G1961), .B(G1956), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(n863), .B(KEYINPUT41), .Z(n865) );
  XNOR2_X1 U965 ( .A(G1986), .B(G1971), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U967 ( .A(G2474), .B(G1966), .Z(n867) );
  XNOR2_X1 U968 ( .A(G1996), .B(G1991), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(G229) );
  NAND2_X1 U971 ( .A1(G124), .A2(n891), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n870), .B(KEYINPUT44), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n896), .A2(G100), .ZN(n871) );
  NAND2_X1 U974 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G136), .A2(n895), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G112), .A2(n892), .ZN(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U978 ( .A1(n876), .A2(n875), .ZN(G162) );
  XOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n879) );
  XOR2_X1 U980 ( .A(n877), .B(KEYINPUT114), .Z(n878) );
  XNOR2_X1 U981 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n1005), .B(n880), .ZN(n890) );
  NAND2_X1 U983 ( .A1(G139), .A2(n895), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G103), .A2(n896), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n888) );
  NAND2_X1 U986 ( .A1(n891), .A2(G127), .ZN(n884) );
  NAND2_X1 U987 ( .A1(G115), .A2(n892), .ZN(n883) );
  NAND2_X1 U988 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U989 ( .A(KEYINPUT47), .B(n885), .ZN(n886) );
  XNOR2_X1 U990 ( .A(KEYINPUT115), .B(n886), .ZN(n887) );
  NOR2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n1014) );
  XNOR2_X1 U992 ( .A(G164), .B(n1014), .ZN(n889) );
  XNOR2_X1 U993 ( .A(n890), .B(n889), .ZN(n905) );
  XNOR2_X1 U994 ( .A(G160), .B(G162), .ZN(n903) );
  NAND2_X1 U995 ( .A1(n891), .A2(G130), .ZN(n894) );
  NAND2_X1 U996 ( .A1(G118), .A2(n892), .ZN(n893) );
  NAND2_X1 U997 ( .A1(n894), .A2(n893), .ZN(n901) );
  NAND2_X1 U998 ( .A1(G142), .A2(n895), .ZN(n898) );
  NAND2_X1 U999 ( .A1(G106), .A2(n896), .ZN(n897) );
  NAND2_X1 U1000 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U1001 ( .A(KEYINPUT45), .B(n899), .Z(n900) );
  NOR2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(n905), .B(n904), .Z(n909) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1008 ( .A(G286), .B(KEYINPUT116), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(G171), .B(n911), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n916) );
  XOR2_X1 U1011 ( .A(n991), .B(n914), .Z(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n917), .ZN(G397) );
  OR2_X1 U1014 ( .A1(n924), .A2(G401), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n918) );
  XOR2_X1 U1016 ( .A(KEYINPUT117), .B(n918), .Z(n919) );
  XNOR2_X1 U1017 ( .A(n919), .B(KEYINPUT49), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(n924), .ZN(G319) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1024 ( .A(G1976), .B(G23), .Z(n926) );
  XOR2_X1 U1025 ( .A(G1971), .B(G22), .Z(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(G24), .B(G1986), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1029 ( .A(KEYINPUT58), .B(n929), .Z(n946) );
  XOR2_X1 U1030 ( .A(G1961), .B(G5), .Z(n941) );
  XOR2_X1 U1031 ( .A(G1981), .B(G6), .Z(n932) );
  XNOR2_X1 U1032 ( .A(n930), .B(G20), .ZN(n931) );
  NAND2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n938) );
  XOR2_X1 U1034 ( .A(G1341), .B(G19), .Z(n936) );
  XOR2_X1 U1035 ( .A(G1348), .B(G4), .Z(n933) );
  XNOR2_X1 U1036 ( .A(KEYINPUT125), .B(n933), .ZN(n934) );
  XNOR2_X1 U1037 ( .A(n934), .B(KEYINPUT59), .ZN(n935) );
  NAND2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1040 ( .A(KEYINPUT60), .B(n939), .ZN(n940) );
  NAND2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(G21), .B(G1966), .ZN(n942) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1044 ( .A(KEYINPUT126), .B(n944), .Z(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1046 ( .A(KEYINPUT61), .B(n947), .Z(n948) );
  NOR2_X1 U1047 ( .A1(G16), .A2(n948), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(KEYINPUT127), .B(n949), .ZN(n1029) );
  XNOR2_X1 U1049 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n1021) );
  XNOR2_X1 U1050 ( .A(n1021), .B(KEYINPUT123), .ZN(n970) );
  XNOR2_X1 U1051 ( .A(G2090), .B(G35), .ZN(n964) );
  XNOR2_X1 U1052 ( .A(KEYINPUT121), .B(G2067), .ZN(n950) );
  XNOR2_X1 U1053 ( .A(n950), .B(G26), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G1996), .B(G32), .ZN(n952) );
  XNOR2_X1 U1055 ( .A(G33), .B(G2072), .ZN(n951) );
  NOR2_X1 U1056 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1057 ( .A1(G28), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1058 ( .A(G25), .B(G1991), .ZN(n954) );
  XNOR2_X1 U1059 ( .A(KEYINPUT120), .B(n954), .ZN(n955) );
  NOR2_X1 U1060 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1061 ( .A1(n958), .A2(n957), .ZN(n961) );
  XNOR2_X1 U1062 ( .A(G27), .B(n959), .ZN(n960) );
  NOR2_X1 U1063 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1064 ( .A(KEYINPUT53), .B(n962), .ZN(n963) );
  NOR2_X1 U1065 ( .A1(n964), .A2(n963), .ZN(n968) );
  XOR2_X1 U1066 ( .A(KEYINPUT122), .B(G34), .Z(n966) );
  XNOR2_X1 U1067 ( .A(G2084), .B(KEYINPUT54), .ZN(n965) );
  XNOR2_X1 U1068 ( .A(n966), .B(n965), .ZN(n967) );
  NAND2_X1 U1069 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1070 ( .A(n970), .B(n969), .ZN(n971) );
  OR2_X1 U1071 ( .A1(G29), .A2(n971), .ZN(n972) );
  NAND2_X1 U1072 ( .A1(G11), .A2(n972), .ZN(n1027) );
  XNOR2_X1 U1073 ( .A(KEYINPUT56), .B(G16), .ZN(n997) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G168), .ZN(n974) );
  NAND2_X1 U1075 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1076 ( .A(KEYINPUT57), .B(n975), .ZN(n995) );
  XNOR2_X1 U1077 ( .A(G301), .B(G1961), .ZN(n978) );
  XNOR2_X1 U1078 ( .A(n976), .B(G1348), .ZN(n977) );
  NOR2_X1 U1079 ( .A1(n978), .A2(n977), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(G166), .B(G1971), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(n979), .B(G1956), .ZN(n981) );
  NAND2_X1 U1082 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1083 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1084 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1085 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1086 ( .A(n988), .B(KEYINPUT124), .ZN(n989) );
  NAND2_X1 U1087 ( .A1(n990), .A2(n989), .ZN(n993) );
  XNOR2_X1 U1088 ( .A(G1341), .B(n991), .ZN(n992) );
  NOR2_X1 U1089 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1090 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n1025) );
  XOR2_X1 U1092 ( .A(G2090), .B(G162), .Z(n998) );
  NOR2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1094 ( .A(KEYINPUT51), .B(n1000), .Z(n1001) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1011) );
  XOR2_X1 U1096 ( .A(G160), .B(G2084), .Z(n1003) );
  NOR2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1100 ( .A(KEYINPUT118), .B(n1009), .Z(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1019) );
  XOR2_X1 U1103 ( .A(G2072), .B(n1014), .Z(n1016) );
  XOR2_X1 U1104 ( .A(G164), .B(G2078), .Z(n1015) );
  NOR2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1106 ( .A(KEYINPUT50), .B(n1017), .Z(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(G29), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

