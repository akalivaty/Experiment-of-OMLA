//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n527, new_n528,
    new_n529, new_n530, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT68), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n460), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n464), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT69), .Z(new_n480));
  AND2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  AOI211_X1 g059(.A(new_n477), .B(new_n480), .C1(G136), .C2(new_n484), .ZN(G162));
  AND2_X1   g060(.A1(KEYINPUT70), .A2(G138), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n464), .B(new_n486), .C1(new_n481), .C2(new_n482), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n463), .A2(KEYINPUT4), .A3(new_n464), .A4(new_n486), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n463), .A2(G126), .A3(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n464), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT71), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(G543), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n500), .A2(new_n503), .B1(KEYINPUT5), .B2(new_n499), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n504), .A2(G62), .ZN(new_n505));
  AND2_X1   g080(.A1(G75), .A2(G543), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n498), .B(G651), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n509), .A2(G88), .B1(G50), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n506), .B1(new_n504), .B2(G62), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT72), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n507), .A2(new_n512), .A3(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND2_X1  g092(.A1(new_n511), .A2(G51), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n504), .A2(G89), .A3(new_n508), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  AOI22_X1  g101(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(new_n514), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT73), .B(G52), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n509), .A2(G90), .B1(new_n511), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(G301));
  INV_X1    g106(.A(G301), .ZN(G171));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n504), .A2(G56), .ZN(new_n534));
  AND2_X1   g109(.A1(G68), .A2(G543), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n533), .B(G651), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n509), .A2(G81), .B1(G43), .B2(new_n511), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n535), .B1(new_n504), .B2(G56), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT74), .B1(new_n538), .B2(new_n514), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT75), .ZN(G188));
  NAND2_X1  g122(.A1(new_n509), .A2(G91), .ZN(new_n548));
  INV_X1    g123(.A(G53), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT9), .B1(new_n510), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT9), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n508), .A2(new_n551), .A3(G53), .A4(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n548), .B(new_n553), .C1(new_n514), .C2(new_n554), .ZN(G299));
  NAND2_X1  g130(.A1(new_n509), .A2(G87), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n511), .A2(G49), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(G288));
  AOI22_X1  g134(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n514), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n504), .A2(new_n508), .ZN(new_n562));
  INV_X1    g137(.A(G86), .ZN(new_n563));
  INV_X1    g138(.A(G48), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n562), .A2(new_n563), .B1(new_n564), .B2(new_n510), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G305));
  AOI22_X1  g142(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n514), .ZN(new_n569));
  INV_X1    g144(.A(G85), .ZN(new_n570));
  INV_X1    g145(.A(G47), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n562), .A2(new_n570), .B1(new_n571), .B2(new_n510), .ZN(new_n572));
  OR3_X1    g147(.A1(new_n569), .A2(new_n572), .A3(KEYINPUT76), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT76), .B1(new_n569), .B2(new_n572), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G290));
  INV_X1    g150(.A(G868), .ZN(new_n576));
  NOR2_X1   g151(.A1(G301), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n504), .A2(G92), .A3(new_n508), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g154(.A1(G79), .A2(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n500), .A2(new_n503), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n511), .A2(G54), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n578), .B(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n585), .A2(G651), .B1(G54), .B2(new_n511), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT77), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n577), .B1(new_n597), .B2(new_n576), .ZN(G284));
  AOI21_X1  g173(.A(new_n577), .B1(new_n597), .B2(new_n576), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(G299), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  XOR2_X1   g177(.A(G280), .B(KEYINPUT78), .Z(G297));
  XNOR2_X1  g178(.A(KEYINPUT79), .B(G559), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(G860), .B2(new_n605), .ZN(G148));
  NAND3_X1  g181(.A1(new_n591), .A2(new_n596), .A3(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n463), .A2(new_n461), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(KEYINPUT12), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT12), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n463), .A2(new_n613), .A3(new_n461), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(G2100), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n475), .A2(G123), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n464), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(G135), .ZN(new_n623));
  OAI221_X1 g198(.A(new_n620), .B1(new_n621), .B2(new_n622), .C1(new_n623), .C2(new_n465), .ZN(new_n624));
  INV_X1    g199(.A(G2096), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n618), .A2(new_n619), .A3(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2430), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2435), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT15), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT15), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G2435), .ZN(new_n635));
  INV_X1    g210(.A(G2438), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT80), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT80), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G2438), .ZN(new_n639));
  AND4_X1   g214(.A1(new_n633), .A2(new_n635), .A3(new_n637), .A4(new_n639), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n633), .A2(new_n635), .B1(new_n637), .B2(new_n639), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n631), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n633), .A2(new_n635), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(new_n639), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g220(.A1(new_n633), .A2(new_n635), .A3(new_n637), .A4(new_n639), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(new_n630), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT81), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n645), .A2(new_n646), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n650), .B1(new_n651), .B2(new_n631), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT81), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(new_n647), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n649), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n656), .B1(new_n649), .B2(new_n654), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n629), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n656), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n653), .B1(new_n652), .B2(new_n647), .ZN(new_n663));
  AND4_X1   g238(.A1(new_n653), .A2(new_n642), .A3(KEYINPUT14), .A4(new_n647), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n649), .A2(new_n654), .A3(new_n656), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n628), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n659), .A2(new_n661), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT82), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n670));
  NAND4_X1  g245(.A1(new_n659), .A2(new_n670), .A3(new_n667), .A4(new_n661), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G14), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n659), .A2(new_n667), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT83), .B1(new_n674), .B2(new_n660), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n676));
  AOI211_X1 g251(.A(new_n676), .B(new_n661), .C1(new_n659), .C2(new_n667), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n673), .A2(new_n678), .ZN(G401));
  INV_X1    g254(.A(KEYINPUT18), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(KEYINPUT17), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(new_n617), .ZN(new_n687));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n683), .B2(KEYINPUT18), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(new_n625), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G1971), .ZN(new_n699));
  INV_X1    g274(.A(G1976), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(G1971), .A2(G1976), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n701), .A2(KEYINPUT19), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT19), .ZN(new_n704));
  INV_X1    g279(.A(new_n702), .ZN(new_n705));
  NOR2_X1   g280(.A1(G1971), .A2(G1976), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1956), .B(G2474), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1961), .B(G1966), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n698), .A2(new_n703), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(new_n703), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n712), .A2(new_n708), .A3(new_n709), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n708), .A2(new_n709), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(KEYINPUT20), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n712), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n721));
  AND3_X1   g296(.A1(new_n714), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n714), .B2(new_n720), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n695), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n714), .A2(new_n720), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(KEYINPUT84), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n714), .A2(new_n720), .A3(new_n721), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n726), .A2(new_n727), .A3(new_n694), .ZN(new_n728));
  XOR2_X1   g303(.A(G1991), .B(G1996), .Z(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n724), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n724), .B2(new_n728), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n693), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n722), .A2(new_n723), .A3(new_n695), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n694), .B1(new_n726), .B2(new_n727), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n729), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n724), .A2(new_n728), .A3(new_n730), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n736), .A2(new_n737), .A3(new_n692), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n733), .A2(new_n738), .ZN(G229));
  INV_X1    g314(.A(G16), .ZN(new_n740));
  NOR2_X1   g315(.A1(G171), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G5), .B2(new_n740), .ZN(new_n742));
  INV_X1    g317(.A(G1961), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n740), .A2(G21), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G168), .B2(new_n740), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n742), .A2(new_n743), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT85), .B(G29), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(G27), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G164), .B2(new_n751), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT96), .B(G2078), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n744), .A2(new_n748), .A3(new_n749), .A4(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G32), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT26), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n475), .A2(G129), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n461), .A2(G105), .ZN(new_n763));
  INV_X1    g338(.A(G141), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n465), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n758), .B1(new_n766), .B2(new_n757), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT27), .B(G1996), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT94), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n767), .B(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT31), .B(G11), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n624), .A2(new_n750), .ZN(new_n773));
  INV_X1    g348(.A(G28), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT30), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(KEYINPUT30), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n772), .B(new_n773), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G2084), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(G34), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(G34), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n750), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT93), .Z(new_n783));
  NAND2_X1  g358(.A1(G160), .A2(G29), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n770), .B(new_n777), .C1(new_n778), .C2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G127), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n483), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(G115), .A2(G2104), .ZN(new_n789));
  OAI21_X1  g364(.A(G2105), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n484), .A2(G139), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT25), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n790), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(new_n757), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n757), .B2(G33), .ZN(new_n798));
  INV_X1    g373(.A(G2072), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n798), .A2(new_n799), .B1(new_n785), .B2(new_n778), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n799), .B2(new_n798), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n756), .A2(new_n786), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT97), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n740), .A2(G4), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n597), .B2(new_n740), .ZN(new_n805));
  INV_X1    g380(.A(G1348), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n751), .A2(G35), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G162), .B2(new_n751), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT29), .B(G2090), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT98), .B(KEYINPUT23), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n740), .A2(G20), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n601), .B2(new_n740), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1956), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n750), .A2(G26), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT28), .ZN(new_n818));
  OAI211_X1 g393(.A(G140), .B(new_n464), .C1(new_n481), .C2(new_n482), .ZN(new_n819));
  OAI211_X1 g394(.A(G128), .B(G2105), .C1(new_n481), .C2(new_n482), .ZN(new_n820));
  OR2_X1    g395(.A1(G104), .A2(G2105), .ZN(new_n821));
  INV_X1    g396(.A(G116), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G2105), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n821), .A2(new_n823), .A3(G2104), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n819), .A2(new_n820), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n818), .B1(new_n757), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT91), .ZN(new_n827));
  INV_X1    g402(.A(G2067), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n811), .A2(new_n816), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(G16), .A2(G19), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n541), .B2(G16), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(G1341), .Z(new_n833));
  NAND3_X1  g408(.A1(new_n807), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n803), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n740), .A2(G22), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G166), .B2(new_n740), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT89), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(new_n699), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n699), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n740), .A2(G23), .ZN(new_n841));
  INV_X1    g416(.A(G288), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n740), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT33), .B(G1976), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(G6), .A2(G16), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n566), .B2(G16), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT32), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G1981), .ZN(new_n852));
  INV_X1    g427(.A(G1981), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n849), .A2(new_n853), .A3(new_n850), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n845), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n839), .A2(new_n840), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(G16), .A2(G24), .ZN(new_n860));
  INV_X1    g435(.A(G290), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(G16), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G1986), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n751), .A2(G25), .ZN(new_n864));
  NOR2_X1   g439(.A1(G95), .A2(G2105), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n460), .B1(new_n865), .B2(KEYINPUT86), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT86), .ZN(new_n867));
  INV_X1    g442(.A(G107), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(G2105), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n866), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n463), .A2(G131), .A3(new_n464), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n463), .A2(G119), .A3(G2105), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT87), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n864), .B1(new_n875), .B2(new_n751), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT88), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G1991), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n863), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n839), .A2(new_n840), .A3(new_n855), .A4(new_n857), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n859), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT36), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT36), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n859), .A2(new_n884), .A3(new_n881), .A4(new_n880), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n835), .A2(new_n886), .ZN(G150));
  INV_X1    g462(.A(G150), .ZN(G311));
  AOI22_X1  g463(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(new_n514), .ZN(new_n890));
  INV_X1    g465(.A(G93), .ZN(new_n891));
  XOR2_X1   g466(.A(KEYINPUT99), .B(G55), .Z(new_n892));
  OAI22_X1  g467(.A1(new_n562), .A2(new_n891), .B1(new_n510), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G860), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT37), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n597), .A2(G559), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(KEYINPUT100), .Z(new_n899));
  INV_X1    g474(.A(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n898), .B(KEYINPUT100), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n890), .A2(new_n893), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n540), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n894), .A2(new_n536), .A3(new_n539), .A4(new_n537), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT39), .ZN(new_n910));
  INV_X1    g485(.A(new_n908), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n901), .A2(new_n911), .A3(new_n903), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n895), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n910), .B1(new_n909), .B2(new_n912), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n897), .B1(new_n914), .B2(new_n915), .ZN(G145));
  OR2_X1    g491(.A1(G106), .A2(G2105), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n917), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n918));
  OAI211_X1 g493(.A(G142), .B(new_n464), .C1(new_n481), .C2(new_n482), .ZN(new_n919));
  OAI211_X1 g494(.A(G130), .B(G2105), .C1(new_n481), .C2(new_n482), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT101), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n918), .A2(new_n919), .A3(new_n920), .A4(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n615), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n615), .A3(new_n924), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n875), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n873), .B(KEYINPUT87), .ZN(new_n929));
  INV_X1    g504(.A(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n929), .B1(new_n930), .B2(new_n925), .ZN(new_n931));
  INV_X1    g506(.A(new_n766), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n819), .A2(new_n820), .A3(new_n824), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n496), .A2(new_n933), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n475), .A2(G126), .B1(new_n492), .B2(new_n494), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n825), .A2(new_n490), .A3(new_n489), .A4(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n934), .A2(new_n936), .A3(new_n795), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n795), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n796), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n934), .A2(new_n936), .A3(new_n795), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n766), .A3(new_n942), .ZN(new_n943));
  AOI221_X4 g518(.A(KEYINPUT102), .B1(new_n928), .B2(new_n931), .C1(new_n939), .C2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n943), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n928), .A2(new_n931), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT103), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n937), .A2(new_n938), .A3(new_n932), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n766), .B1(new_n941), .B2(new_n942), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT102), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n946), .A2(new_n945), .A3(new_n947), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n946), .ZN(new_n957));
  INV_X1    g532(.A(new_n947), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n949), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(G160), .B(new_n624), .ZN(new_n961));
  XNOR2_X1  g536(.A(G162), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT104), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n960), .A2(new_n965), .A3(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n953), .A2(new_n955), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n962), .B1(new_n958), .B2(new_n957), .ZN(new_n968));
  AOI21_X1  g543(.A(G37), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g546(.A1(new_n597), .A2(new_n605), .A3(new_n908), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n607), .A2(new_n911), .ZN(new_n974));
  OAI21_X1  g549(.A(G299), .B1(new_n579), .B2(new_n588), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n554), .A2(new_n514), .ZN(new_n976));
  AOI22_X1  g551(.A1(G91), .A2(new_n509), .B1(new_n550), .B2(new_n552), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n593), .A2(new_n594), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n972), .A2(new_n973), .A3(new_n974), .A4(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n972), .A2(new_n974), .A3(new_n980), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT105), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT41), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n975), .A2(KEYINPUT41), .A3(new_n978), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n972), .B2(new_n974), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n981), .B1(new_n983), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT107), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n991), .B(new_n981), .C1(new_n983), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g567(.A1(G305), .A2(G303), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n566), .A2(new_n507), .A3(new_n515), .A4(new_n512), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n994), .A3(G288), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G288), .B1(new_n993), .B2(new_n994), .ZN(new_n997));
  OAI21_X1  g572(.A(G290), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(new_n994), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n842), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(new_n861), .A3(new_n995), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n1003));
  XNOR2_X1  g578(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n990), .A2(new_n992), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1004), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(new_n989), .A3(KEYINPUT107), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1007), .A3(G868), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n905), .A2(new_n576), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1005), .A2(new_n1007), .A3(KEYINPUT108), .A4(G868), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(G295));
  NAND3_X1  g588(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(G331));
  INV_X1    g589(.A(new_n1002), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n511), .A2(new_n529), .ZN(new_n1016));
  INV_X1    g591(.A(G90), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(new_n562), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n527), .A2(new_n514), .ZN(new_n1019));
  OAI21_X1  g594(.A(G286), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n518), .A2(new_n520), .A3(new_n524), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1021), .A2(new_n528), .A3(new_n519), .A4(new_n530), .ZN(new_n1022));
  AND4_X1   g597(.A1(new_n906), .A2(new_n907), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n906), .A2(new_n907), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n979), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1020), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT109), .B1(new_n908), .B2(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1022), .A2(new_n1020), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n906), .A4(new_n907), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n908), .A2(new_n1026), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n987), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1025), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1033), .A3(KEYINPUT110), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1015), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G37), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n979), .B1(new_n908), .B2(new_n1026), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n985), .B(new_n986), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1039), .B1(new_n1043), .B2(new_n1002), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT43), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1041), .A2(new_n1042), .B1(new_n998), .B2(new_n1001), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1047), .B(new_n1039), .C1(new_n1043), .C2(new_n1002), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1045), .B(KEYINPUT44), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT43), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n1038), .B2(new_n1048), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1049), .B1(new_n1054), .B2(new_n1055), .ZN(G397));
  INV_X1    g631(.A(G1384), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT45), .B1(new_n496), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G125), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n483), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n469), .ZN(new_n1062));
  OAI21_X1  g637(.A(G2105), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n484), .A2(G137), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(G40), .A3(new_n462), .A4(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1059), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  OR3_X1    g642(.A1(new_n1067), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT46), .B1(new_n1067), .B2(G1996), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n933), .B(new_n828), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n766), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1068), .A2(new_n1069), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1072), .B(KEYINPUT47), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1067), .A2(G290), .A3(G1986), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1074), .A2(KEYINPUT48), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n875), .A2(new_n878), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n766), .B(G1996), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n875), .A2(new_n878), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1070), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1066), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(KEYINPUT48), .B2(new_n1074), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1077), .A2(new_n1070), .ZN(new_n1083));
  OAI22_X1  g658(.A1(new_n1083), .A2(new_n1078), .B1(G2067), .B2(new_n933), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1073), .B(new_n1082), .C1(new_n1066), .C2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1057), .A2(KEYINPUT45), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1065), .B1(new_n496), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1059), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n747), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n496), .A2(new_n1057), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1065), .B1(KEYINPUT50), .B2(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1091), .A2(KEYINPUT50), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n778), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G40), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n467), .A2(new_n470), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n496), .A2(new_n1086), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(new_n1058), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT118), .B1(new_n1100), .B2(G1966), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(G8), .B(G168), .C1(new_n1095), .C2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT49), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n566), .A2(new_n853), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT115), .B(G1981), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n561), .A2(new_n565), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1105), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1107), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n566), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1111), .B(KEYINPUT49), .C1(new_n853), .C2(new_n566), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1097), .A2(new_n1057), .A3(new_n496), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G8), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1109), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n556), .A2(G1976), .A3(new_n557), .A4(new_n558), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(G8), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT52), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT52), .B1(G288), .B2(new_n700), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(G8), .A3(new_n1113), .A4(new_n1117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1104), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1109), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1124), .A2(KEYINPUT116), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1103), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT55), .ZN(new_n1127));
  INV_X1    g702(.A(G8), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(G166), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT113), .B(G1971), .Z(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1099), .B2(new_n1058), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT114), .ZN(new_n1135));
  INV_X1    g710(.A(G2090), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1092), .A2(new_n1093), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT114), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1139), .B(new_n1133), .C1(new_n1099), .C2(new_n1058), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  OAI211_X1 g716(.A(G8), .B(new_n1131), .C1(new_n1138), .C2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(G8), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1126), .A2(KEYINPUT63), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1111), .B1(new_n853), .B2(new_n566), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1114), .B1(new_n1147), .B2(new_n1105), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1122), .B1(new_n1112), .B2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1137), .A2(new_n1134), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1129), .B(new_n1130), .C1(new_n1150), .C2(new_n1128), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1142), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1146), .B1(new_n1152), .B2(new_n1103), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1145), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1090), .A2(new_n1101), .A3(G168), .A4(new_n1094), .ZN(new_n1155));
  OAI21_X1  g730(.A(G8), .B1(KEYINPUT122), .B2(KEYINPUT51), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(G8), .B(G286), .C1(new_n1095), .C2(new_n1102), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1158), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT62), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1162), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1164), .A2(new_n1165), .A3(new_n1160), .A4(new_n1159), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT53), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n1088), .B2(G2078), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n743), .ZN(new_n1170));
  INV_X1    g745(.A(G2078), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1100), .A2(KEYINPUT53), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1168), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(G171), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1152), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1163), .A2(new_n1166), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1142), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1124), .A2(new_n700), .A3(new_n842), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1108), .B(KEYINPUT117), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1114), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1154), .A2(new_n1176), .A3(new_n1181), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1168), .A2(new_n1170), .A3(new_n1172), .A4(G301), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1174), .A2(KEYINPUT54), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(KEYINPUT124), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1174), .A2(new_n1186), .A3(KEYINPUT54), .A4(new_n1183), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT123), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1174), .A2(new_n1189), .A3(new_n1183), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1183), .ZN(new_n1191));
  AOI21_X1  g766(.A(KEYINPUT54), .B1(new_n1191), .B2(KEYINPUT123), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1152), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1164), .A2(new_n1160), .A3(new_n1159), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1188), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT57), .ZN(new_n1197));
  XNOR2_X1  g772(.A(G299), .B(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(G1956), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1169), .A2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(KEYINPUT56), .B(G2072), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1100), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1198), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  OR2_X1    g778(.A1(new_n1203), .A2(KEYINPUT119), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1203), .A2(KEYINPUT119), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1113), .A2(G2067), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1206), .B1(new_n1169), .B2(new_n806), .ZN(new_n1207));
  OAI211_X1 g782(.A(new_n1204), .B(new_n1205), .C1(new_n595), .C2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1200), .A2(new_n1198), .A3(new_n1202), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  XOR2_X1   g785(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1211));
  INV_X1    g786(.A(G1996), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1087), .A2(new_n1212), .A3(new_n1059), .ZN(new_n1213));
  XOR2_X1   g788(.A(KEYINPUT58), .B(G1341), .Z(new_n1214));
  NAND2_X1  g789(.A1(new_n1113), .A2(new_n1214), .ZN(new_n1215));
  AOI211_X1 g790(.A(new_n540), .B(new_n1211), .C1(new_n1213), .C2(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT120), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1219), .A2(new_n541), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1216), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1209), .B1(new_n1203), .B2(KEYINPUT61), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n1223));
  NAND4_X1  g798(.A1(new_n1200), .A2(new_n1198), .A3(new_n1223), .A4(new_n1202), .ZN(new_n1224));
  AND3_X1   g799(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n589), .B1(new_n1207), .B2(KEYINPUT60), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1226), .A2(KEYINPUT121), .ZN(new_n1227));
  AND2_X1   g802(.A1(new_n1207), .A2(KEYINPUT60), .ZN(new_n1228));
  INV_X1    g803(.A(KEYINPUT121), .ZN(new_n1229));
  OAI211_X1 g804(.A(new_n1229), .B(new_n589), .C1(new_n1207), .C2(KEYINPUT60), .ZN(new_n1230));
  AND3_X1   g805(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g806(.A(new_n1228), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1225), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  AOI22_X1  g808(.A1(new_n1195), .A2(new_n1196), .B1(new_n1210), .B2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g809(.A1(new_n1188), .A2(new_n1193), .A3(KEYINPUT125), .A4(new_n1194), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1182), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  AND3_X1   g811(.A1(G290), .A2(G1986), .A3(new_n1066), .ZN(new_n1237));
  NOR2_X1   g812(.A1(new_n1074), .A2(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g813(.A(new_n1238), .B(KEYINPUT112), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1239), .A2(new_n1080), .ZN(new_n1240));
  OAI21_X1  g815(.A(new_n1085), .B1(new_n1236), .B2(new_n1240), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g816(.A(new_n969), .ZN(new_n1243));
  AOI21_X1  g817(.A(new_n1243), .B1(new_n963), .B2(KEYINPUT104), .ZN(new_n1244));
  OR2_X1    g818(.A1(G227), .A2(new_n458), .ZN(new_n1245));
  AOI21_X1  g819(.A(new_n1245), .B1(new_n733), .B2(new_n738), .ZN(new_n1246));
  OAI21_X1  g820(.A(new_n1246), .B1(new_n673), .B2(new_n678), .ZN(new_n1247));
  NAND2_X1  g821(.A1(new_n1247), .A2(KEYINPUT126), .ZN(new_n1248));
  INV_X1    g822(.A(KEYINPUT126), .ZN(new_n1249));
  OAI211_X1 g823(.A(new_n1246), .B(new_n1249), .C1(new_n673), .C2(new_n678), .ZN(new_n1250));
  AOI22_X1  g824(.A1(new_n1244), .A2(new_n966), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g825(.A(KEYINPUT127), .B1(new_n1251), .B2(new_n1051), .ZN(new_n1252));
  NAND2_X1  g826(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1253));
  AND4_X1   g827(.A1(KEYINPUT127), .A2(new_n970), .A3(new_n1253), .A4(new_n1051), .ZN(new_n1254));
  NOR2_X1   g828(.A1(new_n1252), .A2(new_n1254), .ZN(G308));
  NAND2_X1  g829(.A1(new_n1251), .A2(new_n1051), .ZN(G225));
endmodule


