//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n206), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT65), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(new_n203), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT66), .Z(new_n229));
  AOI211_X1 g0029(.A(new_n214), .B(new_n229), .C1(KEYINPUT1), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G20), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G50), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT69), .ZN(new_n250));
  INV_X1    g0050(.A(G13), .ZN(new_n251));
  NOR3_X1   g0051(.A1(new_n251), .A2(new_n208), .A3(G1), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n207), .B1(new_n203), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G50), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n250), .A2(new_n255), .B1(new_n256), .B2(new_n252), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n253), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n258), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G50), .A2(G58), .ZN(new_n265));
  INV_X1    g0065(.A(G68), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n208), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n254), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n257), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g0069(.A(new_n269), .B(KEYINPUT9), .Z(new_n270));
  AND2_X1   g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  OAI21_X1  g0071(.A(G274), .B1(new_n271), .B2(new_n207), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT67), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  AND2_X1   g0075(.A1(G1), .A2(G13), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n278), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n271), .A2(new_n207), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n285), .B1(G226), .B2(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n288), .A2(KEYINPUT68), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G222), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G77), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(G1698), .ZN(new_n294));
  INV_X1    g0094(.A(G223), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n292), .B1(new_n293), .B2(new_n290), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n286), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(new_n288), .B2(KEYINPUT68), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n270), .B1(new_n299), .B2(G190), .ZN(new_n300));
  OAI21_X1  g0100(.A(G200), .B1(new_n289), .B2(new_n298), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n300), .A2(new_n304), .A3(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n299), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(new_n269), .C1(G169), .C2(new_n299), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n252), .A2(new_n266), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT12), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n259), .A2(G77), .B1(G20), .B2(new_n266), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n256), .B2(new_n263), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n255), .A2(G68), .A3(new_n248), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT11), .B1(new_n313), .B2(new_n254), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G97), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n232), .A2(G1698), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(G226), .B2(G1698), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n320), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(new_n286), .B1(new_n287), .B2(G238), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n284), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT13), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(new_n331), .A3(new_n284), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(G179), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n332), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n331), .B1(new_n328), .B2(new_n284), .ZN(new_n335));
  OAI21_X1  g0135(.A(G169), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n333), .B1(new_n336), .B2(KEYINPUT14), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT14), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n330), .A2(new_n332), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(G169), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n319), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(G200), .ZN(new_n342));
  INV_X1    g0142(.A(G190), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n342), .B(new_n318), .C1(new_n343), .C2(new_n339), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n285), .B1(G244), .B2(new_n287), .ZN(new_n346));
  INV_X1    g0146(.A(G238), .ZN(new_n347));
  INV_X1    g0147(.A(G107), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n294), .A2(new_n347), .B1(new_n348), .B2(new_n290), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n326), .A2(new_n232), .A3(G1698), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n286), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G200), .ZN(new_n353));
  INV_X1    g0153(.A(new_n254), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n357));
  INV_X1    g0157(.A(new_n258), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n262), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n354), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n255), .A2(G77), .A3(new_n248), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT70), .B1(new_n252), .B2(new_n293), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n252), .A2(KEYINPUT70), .A3(new_n293), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n353), .B(new_n365), .C1(new_n343), .C2(new_n352), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n352), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n346), .A2(new_n307), .A3(new_n351), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n306), .A2(new_n309), .A3(new_n345), .A4(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT7), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(G20), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT71), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n253), .ZN(new_n377));
  NAND2_X1  g0177(.A1(KEYINPUT71), .A2(G33), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT3), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n325), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n375), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n374), .B1(new_n290), .B2(G20), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n266), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G58), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n266), .ZN(new_n385));
  NOR2_X1   g0185(.A1(G58), .A2(G68), .ZN(new_n386));
  OAI21_X1  g0186(.A(G20), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n262), .A2(G159), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n373), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n373), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n377), .A2(KEYINPUT3), .A3(new_n378), .ZN(new_n392));
  AOI21_X1  g0192(.A(G20), .B1(new_n392), .B2(new_n324), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n393), .B2(new_n374), .ZN(new_n394));
  AOI211_X1 g0194(.A(KEYINPUT7), .B(G20), .C1(new_n392), .C2(new_n324), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n391), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(new_n396), .A3(new_n254), .ZN(new_n397));
  INV_X1    g0197(.A(G200), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n287), .A2(G232), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n272), .A2(KEYINPUT67), .A3(new_n273), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n279), .B1(new_n278), .B2(new_n282), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n403));
  MUX2_X1   g0203(.A(G223), .B(G226), .S(G1698), .Z(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(new_n392), .A3(new_n324), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n398), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n274), .A2(new_n283), .B1(new_n287), .B2(G232), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n405), .A2(new_n406), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n409), .B(new_n343), .C1(new_n410), .C2(new_n403), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n358), .A2(new_n248), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n255), .B1(new_n252), .B2(new_n258), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n397), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT17), .ZN(new_n417));
  INV_X1    g0217(.A(new_n415), .ZN(new_n418));
  INV_X1    g0218(.A(new_n324), .ZN(new_n419));
  AND2_X1   g0219(.A1(KEYINPUT71), .A2(G33), .ZN(new_n420));
  NOR2_X1   g0220(.A1(KEYINPUT71), .A2(G33), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n419), .B1(new_n422), .B2(KEYINPUT3), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT7), .B1(new_n423), .B2(G20), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n393), .A2(new_n374), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(G68), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n354), .B1(new_n426), .B2(new_n391), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n418), .B1(new_n427), .B2(new_n390), .ZN(new_n428));
  OAI21_X1  g0228(.A(G169), .B1(new_n402), .B2(new_n407), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n409), .B(G179), .C1(new_n410), .C2(new_n403), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT18), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT72), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n397), .A2(new_n415), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n429), .A2(new_n430), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n433), .B1(new_n432), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n417), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n372), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G283), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n442), .B(new_n208), .C1(G33), .C2(new_n218), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT20), .ZN(new_n444));
  INV_X1    g0244(.A(G116), .ZN(new_n445));
  AOI22_X1  g0245(.A1(KEYINPUT80), .A2(new_n444), .B1(new_n445), .B2(G20), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n446), .A3(new_n254), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n444), .A2(KEYINPUT80), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n448), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n443), .A2(new_n446), .A3(new_n450), .A4(new_n254), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n252), .A2(new_n445), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT73), .B1(new_n253), .B2(G1), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT73), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(new_n247), .A3(G33), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n255), .A2(new_n454), .A3(G116), .A4(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n255), .A2(G116), .A3(new_n458), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT79), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n453), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(G257), .A2(G1698), .ZN(new_n463));
  INV_X1    g0263(.A(G264), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n464), .B2(G1698), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(new_n392), .A3(new_n324), .ZN(new_n466));
  XOR2_X1   g0266(.A(KEYINPUT78), .B(G303), .Z(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n326), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n286), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n247), .B(G45), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G270), .A3(new_n403), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n247), .A2(G45), .ZN(new_n475));
  INV_X1    g0275(.A(new_n472), .ZN(new_n476));
  NAND2_X1  g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n278), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n470), .A2(G179), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT81), .B1(new_n462), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n461), .A2(new_n459), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT81), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n403), .B1(new_n466), .B2(new_n468), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n474), .A2(new_n479), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n487), .A2(new_n488), .A3(new_n307), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n470), .A2(new_n480), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G169), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n494), .B2(new_n462), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n485), .A2(new_n493), .A3(KEYINPUT21), .A4(G169), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(G200), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(new_n462), .C1(new_n343), .C2(new_n493), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n491), .A2(new_n495), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n478), .A2(new_n464), .A3(new_n286), .ZN(new_n500));
  NOR2_X1   g0300(.A1(G250), .A2(G1698), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n219), .B2(G1698), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(new_n392), .A3(new_n324), .ZN(new_n503));
  XNOR2_X1  g0303(.A(KEYINPUT71), .B(G33), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G294), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n500), .B1(new_n506), .B2(new_n286), .ZN(new_n507));
  AOI21_X1  g0307(.A(G169), .B1(new_n507), .B2(new_n479), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n403), .B1(new_n503), .B2(new_n505), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n473), .A2(new_n272), .ZN(new_n510));
  NOR4_X1   g0310(.A1(new_n509), .A2(new_n500), .A3(G179), .A4(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n392), .A2(new_n208), .A3(G87), .A4(new_n324), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT22), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(new_n208), .A3(G87), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT82), .B1(new_n326), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT82), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n216), .A2(KEYINPUT22), .A3(G20), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n290), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n513), .A2(KEYINPUT22), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n504), .A2(new_n208), .A3(G116), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT23), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n208), .B2(G107), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n348), .A2(KEYINPUT23), .A3(G20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT24), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n513), .A2(KEYINPUT22), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n516), .A2(new_n519), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  INV_X1    g0331(.A(new_n526), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n354), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n255), .A2(new_n458), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G107), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n252), .A2(new_n348), .ZN(new_n538));
  XNOR2_X1  g0338(.A(KEYINPUT83), .B(KEYINPUT25), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n512), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n531), .B1(new_n530), .B2(new_n532), .ZN(new_n543));
  AOI211_X1 g0343(.A(KEYINPUT24), .B(new_n526), .C1(new_n528), .C2(new_n529), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n254), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n541), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n506), .A2(new_n286), .ZN(new_n547));
  INV_X1    g0347(.A(new_n500), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n547), .A2(new_n343), .A3(new_n548), .A4(new_n479), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n509), .A2(new_n500), .A3(new_n510), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(G200), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n545), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n542), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n499), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n348), .B1(new_n381), .B2(new_n382), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT6), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n556), .A2(new_n218), .A3(G107), .ZN(new_n557));
  XNOR2_X1  g0357(.A(G97), .B(G107), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n557), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n559), .A2(new_n208), .B1(new_n293), .B2(new_n263), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n254), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n252), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(G97), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n536), .B2(G97), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g0365(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n392), .A2(new_n324), .ZN(new_n567));
  INV_X1    g0367(.A(G244), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(G1698), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n566), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n569), .A2(new_n324), .A3(new_n325), .A4(KEYINPUT4), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n324), .A2(new_n325), .A3(G250), .A4(G1698), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n572), .A2(new_n573), .A3(new_n442), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n403), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n473), .A2(new_n403), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n479), .B1(new_n576), .B2(new_n219), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n398), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n575), .A2(G190), .A3(new_n577), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n565), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n561), .A2(new_n564), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n367), .B1(new_n575), .B2(new_n577), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n571), .A2(new_n574), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n577), .B1(new_n584), .B2(new_n286), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n582), .B(new_n583), .C1(new_n586), .C2(G179), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n535), .A2(new_n216), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n259), .A2(new_n590), .A3(G97), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G97), .A2(G107), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n216), .B1(new_n320), .B2(new_n208), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n591), .B1(new_n593), .B2(new_n590), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n392), .A2(new_n208), .A3(G68), .A4(new_n324), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n354), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n356), .A2(new_n562), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n589), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT75), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n281), .B2(G1), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n247), .A2(KEYINPUT75), .A3(G45), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n217), .B1(new_n276), .B2(new_n277), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT76), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT76), .B1(new_n602), .B2(new_n603), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n604), .A2(new_n605), .B1(new_n272), .B2(new_n475), .ZN(new_n606));
  NOR2_X1   g0406(.A1(G238), .A2(G1698), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n568), .B2(G1698), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n392), .A3(new_n324), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n504), .A2(G116), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n403), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(G200), .B1(new_n606), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n611), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n272), .A2(new_n475), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n602), .A2(new_n603), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT76), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT76), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n598), .B(new_n612), .C1(new_n343), .C2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n597), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n594), .A2(new_n595), .ZN(new_n623));
  OAI221_X1 g0423(.A(new_n622), .B1(new_n355), .B2(new_n535), .C1(new_n623), .C2(new_n354), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n613), .A2(new_n619), .A3(new_n307), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n367), .B1(new_n606), .B2(new_n611), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT77), .B1(new_n588), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n585), .A2(new_n343), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n578), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n307), .A2(new_n585), .B1(new_n561), .B2(new_n564), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n565), .A2(new_n631), .B1(new_n632), .B2(new_n583), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT77), .ZN(new_n634));
  INV_X1    g0434(.A(new_n628), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n441), .A2(new_n554), .A3(new_n629), .A4(new_n636), .ZN(G372));
  INV_X1    g0437(.A(KEYINPUT84), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n628), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n621), .A2(new_n627), .A3(KEYINPUT84), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n639), .A2(new_n633), .A3(new_n552), .A4(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n491), .A2(new_n495), .A3(new_n496), .ZN(new_n642));
  INV_X1    g0442(.A(new_n542), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(new_n587), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n639), .A2(new_n646), .A3(new_n647), .A4(new_n640), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT26), .B1(new_n628), .B2(new_n587), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n627), .A3(new_n649), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n441), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n428), .A2(KEYINPUT85), .A3(new_n431), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT85), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n434), .B2(new_n436), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n435), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT85), .B1(new_n428), .B2(new_n431), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n434), .A2(new_n654), .A3(new_n436), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(KEYINPUT18), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT17), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n416), .B(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n370), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n344), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n664), .B2(new_n341), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n306), .B1(new_n660), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(new_n309), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n652), .A2(new_n667), .ZN(G369));
  INV_X1    g0468(.A(G330), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n247), .A2(new_n208), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n485), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT86), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n499), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n642), .A2(new_n677), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n669), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n643), .A2(new_n675), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n675), .B1(new_n534), .B2(new_n541), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n542), .A2(new_n682), .A3(new_n552), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n675), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n642), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(new_n553), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n643), .A2(new_n686), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(KEYINPUT87), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT87), .B1(new_n688), .B2(new_n689), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n685), .B1(new_n691), .B2(new_n692), .ZN(G399));
  NAND3_X1  g0493(.A1(new_n592), .A2(new_n216), .A3(new_n445), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n204), .A2(new_n280), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(new_n696), .A3(G1), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n213), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n554), .A2(new_n629), .A3(new_n636), .A4(new_n686), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n606), .A2(new_n611), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n585), .A2(new_n701), .A3(new_n489), .A4(new_n507), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n507), .A2(new_n619), .A3(new_n613), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(KEYINPUT30), .A3(new_n489), .A4(new_n585), .ZN(new_n706));
  INV_X1    g0506(.A(new_n550), .ZN(new_n707));
  AOI21_X1  g0507(.A(G179), .B1(new_n470), .B2(new_n480), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n586), .A2(new_n707), .A3(new_n620), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n704), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT31), .B1(new_n710), .B2(new_n675), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n700), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT88), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT88), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n717), .A3(G330), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n627), .A2(KEYINPUT89), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT89), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n624), .A2(new_n626), .A3(new_n721), .A4(new_n625), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n628), .A2(new_n587), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n646), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n621), .A2(new_n627), .A3(KEYINPUT84), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT84), .B1(new_n621), .B2(new_n627), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n726), .A2(new_n727), .A3(new_n587), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n725), .B1(new_n728), .B2(new_n646), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n686), .B1(new_n729), .B2(new_n645), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n645), .A2(new_n650), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n732), .A2(KEYINPUT29), .A3(new_n675), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n719), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n699), .B1(new_n734), .B2(G1), .ZN(G364));
  NOR2_X1   g0535(.A1(new_n251), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n247), .B1(new_n736), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n696), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n290), .A2(new_n204), .ZN(new_n741));
  INV_X1    g0541(.A(G355), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n741), .A2(new_n742), .B1(G116), .B2(new_n204), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n242), .A2(G45), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n567), .A2(new_n204), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n281), .B2(new_n212), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n743), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n207), .B1(G20), .B2(new_n367), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n740), .B1(new_n747), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n208), .A2(new_n307), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G190), .A3(new_n398), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n290), .B1(new_n756), .B2(new_n384), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G190), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n757), .B1(G77), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n755), .A2(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n343), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(G190), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G50), .A2(new_n763), .B1(new_n764), .B2(G68), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n208), .A2(G179), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n758), .ZN(new_n767));
  INV_X1    g0567(.A(G159), .ZN(new_n768));
  OR3_X1    g0568(.A1(new_n767), .A2(KEYINPUT32), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(KEYINPUT32), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n761), .A2(new_n765), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n766), .A2(G190), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n216), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n343), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n208), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n218), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n766), .A2(new_n343), .A3(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n348), .ZN(new_n778));
  NOR4_X1   g0578(.A1(new_n771), .A2(new_n773), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT90), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT90), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  INV_X1    g0582(.A(G329), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n777), .A2(new_n782), .B1(new_n767), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT91), .ZN(new_n785));
  INV_X1    g0585(.A(new_n764), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT33), .B(G317), .Z(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n775), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n763), .A2(G326), .ZN(new_n790));
  INV_X1    g0590(.A(G303), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n791), .B2(new_n772), .ZN(new_n792));
  INV_X1    g0592(.A(G311), .ZN(new_n793));
  INV_X1    g0593(.A(G322), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n326), .B1(new_n759), .B2(new_n793), .C1(new_n794), .C2(new_n756), .ZN(new_n795));
  OR4_X1    g0595(.A1(new_n785), .A2(new_n789), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n780), .A2(new_n781), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n754), .B1(new_n797), .B2(new_n751), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n678), .A2(new_n679), .ZN(new_n799));
  INV_X1    g0599(.A(new_n750), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n680), .A2(new_n740), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n799), .A2(G330), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT92), .Z(G396));
  INV_X1    g0605(.A(KEYINPUT96), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n370), .A2(new_n675), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n366), .B1(new_n365), .B2(new_n686), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n370), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n732), .B2(new_n675), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n686), .B(new_n809), .C1(new_n645), .C2(new_n650), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n719), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n806), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n740), .B(new_n816), .C1(new_n719), .C2(new_n813), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n814), .A2(new_n815), .A3(new_n806), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n751), .ZN(new_n820));
  INV_X1    g0620(.A(new_n756), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n776), .B1(G294), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT93), .Z(new_n823));
  OAI21_X1  g0623(.A(new_n326), .B1(new_n767), .B2(new_n793), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G116), .B2(new_n760), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n777), .A2(new_n216), .ZN(new_n826));
  INV_X1    g0626(.A(new_n772), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(G107), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G283), .A2(new_n764), .B1(new_n763), .B2(G303), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n823), .A2(new_n825), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n821), .A2(G143), .B1(new_n760), .B2(G159), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  INV_X1    g0632(.A(new_n763), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n831), .B1(new_n786), .B2(new_n261), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT94), .Z(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n836));
  INV_X1    g0636(.A(new_n777), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(G68), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(new_n256), .B2(new_n772), .C1(new_n384), .C2(new_n775), .ZN(new_n839));
  INV_X1    g0639(.A(new_n767), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n567), .B(new_n839), .C1(G132), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n830), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT95), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n820), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n845), .B2(new_n844), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n751), .A2(new_n748), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n739), .B(new_n738), .C1(new_n293), .C2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(new_n749), .C2(new_n809), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n819), .A2(new_n850), .ZN(G384));
  INV_X1    g0651(.A(new_n559), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n445), .B(new_n210), .C1(new_n852), .C2(KEYINPUT35), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(KEYINPUT35), .B2(new_n852), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT36), .Z(new_n855));
  OAI211_X1 g0655(.A(new_n212), .B(G77), .C1(new_n384), .C2(new_n266), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n256), .A2(G68), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n247), .B(G13), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n807), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n812), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n318), .A2(new_n686), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n341), .A2(new_n344), .A3(new_n864), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n337), .A2(new_n340), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n865), .A2(KEYINPUT97), .B1(new_n866), .B2(new_n863), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT97), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n341), .A2(new_n344), .A3(new_n868), .A4(new_n864), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n862), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n397), .A2(new_n412), .A3(new_n415), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n673), .B1(new_n397), .B2(new_n415), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT98), .B1(new_n428), .B2(new_n431), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT98), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n434), .A2(new_n878), .A3(new_n436), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n394), .A2(new_n395), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n373), .B1(new_n881), .B2(new_n389), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n418), .B1(new_n882), .B2(new_n427), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n416), .B1(new_n883), .B2(new_n673), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n431), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n880), .A2(KEYINPUT99), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT99), .B1(new_n880), .B2(new_n886), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n432), .A2(new_n437), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT72), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n662), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n883), .A2(new_n673), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n887), .A2(new_n888), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n440), .A2(new_n893), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n898), .B(KEYINPUT38), .C1(new_n888), .C2(new_n887), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n872), .A2(new_n900), .B1(new_n660), .B2(new_n673), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n416), .B1(new_n428), .B2(new_n673), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n657), .B2(new_n658), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n880), .B1(new_n903), .B2(new_n876), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n662), .B1(new_n656), .B2(new_n659), .ZN(new_n905));
  INV_X1    g0705(.A(new_n874), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n896), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n897), .A2(KEYINPUT39), .A3(new_n899), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n866), .A2(new_n319), .A3(new_n686), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n901), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n441), .B1(new_n731), .B2(new_n733), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n667), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n916), .B(new_n918), .Z(new_n919));
  AOI21_X1  g0719(.A(new_n810), .B1(new_n867), .B2(new_n869), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n710), .A2(new_n675), .ZN(new_n921));
  NOR2_X1   g0721(.A1(KEYINPUT100), .A2(KEYINPUT31), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n700), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT101), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT40), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n920), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n899), .B2(new_n897), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n920), .A2(new_n925), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n909), .B(new_n928), .C1(new_n930), .C2(KEYINPUT101), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n931), .B2(KEYINPUT40), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n441), .A2(new_n925), .ZN(new_n933));
  OAI21_X1  g0733(.A(G330), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n933), .B2(new_n932), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n919), .A2(new_n935), .B1(new_n247), .B2(new_n736), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n919), .A2(new_n935), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n859), .B1(new_n936), .B2(new_n937), .ZN(G367));
  INV_X1    g0738(.A(KEYINPUT109), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n688), .B(KEYINPUT107), .Z(new_n940));
  OR2_X1    g0740(.A1(new_n680), .A2(KEYINPUT108), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n687), .A2(new_n681), .A3(new_n683), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n680), .A2(KEYINPUT108), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n734), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n685), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n688), .A2(new_n689), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT87), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n633), .B1(new_n565), .B2(new_n686), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n647), .A2(new_n675), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n951), .A2(new_n690), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT105), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT44), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n951), .A2(new_n690), .A3(new_n955), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n957), .A2(new_n958), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n954), .B1(new_n691), .B2(new_n692), .ZN(new_n964));
  XNOR2_X1  g0764(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n954), .B(new_n965), .C1(new_n691), .C2(new_n692), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(KEYINPUT106), .B(new_n948), .C1(new_n963), .C2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n969), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n685), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n947), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n972), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT106), .B1(new_n975), .B2(new_n948), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n734), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n696), .B(KEYINPUT41), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n738), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n955), .A2(new_n688), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT42), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n587), .B1(new_n952), .B2(new_n542), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n686), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n598), .A2(new_n686), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n639), .A2(new_n640), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n627), .B2(new_n986), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n988), .A2(KEYINPUT102), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(KEYINPUT102), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT43), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n985), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT103), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n948), .A2(new_n954), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n991), .B1(new_n985), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n994), .A2(new_n993), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n939), .B1(new_n980), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n948), .B1(new_n963), .B2(new_n969), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT106), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1005), .A2(new_n970), .A3(new_n947), .A4(new_n973), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n978), .B1(new_n1006), .B2(new_n734), .ZN(new_n1007));
  OAI211_X1 g0807(.A(KEYINPUT109), .B(new_n1000), .C1(new_n1007), .C2(new_n738), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n752), .B1(new_n204), .B2(new_n355), .C1(new_n238), .C2(new_n745), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n290), .B1(new_n767), .B2(new_n832), .C1(new_n256), .C2(new_n759), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n837), .A2(G77), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n786), .B2(new_n768), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(G58), .C2(new_n827), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT111), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n763), .A2(G143), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n266), .B2(new_n775), .C1(new_n261), .C2(new_n756), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1014), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT112), .Z(new_n1020));
  NAND3_X1  g0820(.A1(new_n827), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT110), .Z(new_n1022));
  INV_X1    g0822(.A(new_n775), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1023), .A2(G107), .B1(new_n837), .B2(G97), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n788), .B2(new_n786), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n821), .A2(new_n467), .B1(new_n840), .B2(G317), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n782), .B2(new_n759), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT46), .B1(new_n827), .B2(G116), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n567), .B1(new_n833), .B2(new_n793), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1020), .B1(new_n1022), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT47), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n740), .B(new_n1010), .C1(new_n1032), .C2(new_n820), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n988), .A2(new_n800), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1009), .A2(new_n1036), .ZN(G387));
  NOR2_X1   g0837(.A1(new_n947), .A2(new_n696), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n944), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n943), .B(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1038), .B1(new_n734), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n681), .A2(new_n683), .A3(new_n750), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n741), .A2(new_n695), .B1(G107), .B2(new_n204), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n235), .A2(new_n281), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n258), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI211_X1 g0846(.A(G45), .B(new_n694), .C1(G68), .C2(G77), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n745), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1043), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n740), .B1(new_n1049), .B2(new_n753), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n772), .A2(new_n293), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G97), .B2(new_n837), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(KEYINPUT113), .B(G150), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1052), .B(new_n423), .C1(new_n767), .C2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT114), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n756), .A2(new_n256), .B1(new_n759), .B2(new_n266), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G159), .B2(new_n763), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n356), .A2(new_n1023), .B1(new_n764), .B2(new_n358), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n423), .B1(G326), .B2(new_n840), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n775), .A2(new_n782), .B1(new_n772), .B2(new_n788), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n821), .A2(G317), .B1(new_n760), .B2(new_n467), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n786), .B2(new_n793), .C1(new_n794), .C2(new_n833), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT49), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1060), .B1(new_n445), .B2(new_n777), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1059), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT115), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n820), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1050), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1040), .A2(new_n738), .B1(new_n1042), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1041), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT116), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1041), .A2(KEYINPUT116), .A3(new_n1075), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(G393));
  OAI221_X1 g0880(.A(new_n752), .B1(new_n218), .B2(new_n204), .C1(new_n245), .C2(new_n745), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n740), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n833), .A2(new_n261), .B1(new_n768), .B2(new_n756), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT51), .Z(new_n1084));
  OAI22_X1  g0884(.A1(new_n786), .A2(new_n256), .B1(new_n772), .B2(new_n266), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n775), .A2(new_n293), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1085), .A2(new_n826), .A3(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n358), .A2(new_n760), .B1(new_n840), .B2(G143), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n423), .A3(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G317), .A2(new_n763), .B1(new_n821), .B2(G311), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n326), .B1(new_n759), .B2(new_n788), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G322), .B2(new_n840), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n778), .B1(G116), .B2(new_n1023), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n764), .A2(new_n467), .B1(new_n827), .B2(G283), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1084), .A2(new_n1089), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1082), .B1(new_n1097), .B2(new_n751), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n954), .B2(new_n800), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1003), .A2(new_n973), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n737), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1040), .A2(new_n734), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n696), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1101), .B1(new_n1006), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(G390));
  AOI21_X1  g0905(.A(new_n669), .B1(new_n924), .B2(new_n700), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n920), .A2(new_n1106), .A3(KEYINPUT117), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT117), .B1(new_n920), .B2(new_n1106), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n914), .B1(new_n861), .B2(new_n870), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n897), .A2(KEYINPUT39), .A3(new_n899), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT39), .B1(new_n899), .B2(new_n908), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n808), .A2(new_n370), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n686), .B(new_n1115), .C1(new_n729), .C2(new_n645), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n860), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n870), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n913), .A3(new_n909), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1109), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1110), .B1(new_n911), .B2(new_n912), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1118), .A2(new_n909), .A3(new_n913), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n717), .B1(new_n714), .B2(G330), .ZN(new_n1123));
  AOI211_X1 g0923(.A(KEYINPUT88), .B(new_n669), .C1(new_n700), .C2(new_n713), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n809), .B(new_n870), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1121), .A2(new_n1122), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1120), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n748), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n848), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n740), .B1(new_n358), .B2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT119), .Z(new_n1132));
  NOR2_X1   g0932(.A1(new_n786), .A2(new_n348), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1086), .B(new_n1133), .C1(G283), .C2(new_n763), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n773), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n756), .A2(new_n445), .B1(new_n767), .B2(new_n788), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n290), .B(new_n1136), .C1(G97), .C2(new_n760), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n838), .A4(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n772), .A2(new_n1053), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT53), .ZN(new_n1140));
  INV_X1    g0940(.A(G132), .ZN(new_n1141));
  INV_X1    g0941(.A(G125), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n756), .A2(new_n1141), .B1(new_n767), .B2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT54), .B(G143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n290), .B1(new_n759), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n763), .A2(G128), .B1(new_n837), .B2(G50), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G159), .A2(new_n1023), .B1(new_n764), .B2(G137), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1140), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT120), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1150), .A2(new_n820), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1138), .A2(KEYINPUT120), .A3(new_n1149), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1132), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1128), .A2(new_n738), .B1(new_n1129), .B2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT121), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1114), .A2(new_n1119), .A3(new_n1125), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n920), .A2(new_n1106), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT117), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n920), .A2(new_n1106), .A3(KEYINPUT117), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1156), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n441), .A2(new_n1106), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n917), .A2(new_n667), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n809), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n871), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n862), .B1(new_n1168), .B2(new_n1109), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1106), .A2(new_n809), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1117), .B1(new_n871), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1125), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1166), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(KEYINPUT118), .B1(new_n1163), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n870), .B1(new_n719), .B2(new_n809), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n861), .B1(new_n1176), .B2(new_n1161), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1165), .B1(new_n1177), .B2(new_n1172), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT118), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1178), .A2(new_n1179), .A3(new_n1156), .A4(new_n1162), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n739), .C1(new_n1128), .C2(new_n1178), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1155), .A2(new_n1182), .ZN(G378));
  NAND2_X1  g0983(.A1(new_n306), .A2(new_n309), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n673), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n269), .A2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1184), .B(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1187), .B(new_n1188), .Z(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n932), .A2(new_n669), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1189), .B1(new_n932), .B2(new_n669), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n916), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n915), .A3(new_n901), .A4(new_n1193), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n738), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n740), .B1(G50), .B2(new_n1130), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n356), .A2(new_n760), .B1(new_n840), .B2(G283), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n348), .B2(new_n756), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1051), .B(new_n1201), .C1(G68), .C2(new_n1023), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n833), .A2(new_n445), .B1(new_n777), .B2(new_n384), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G97), .B2(new_n764), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1202), .A2(new_n280), .A3(new_n567), .A4(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT58), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n567), .A2(new_n280), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G50), .B1(new_n253), .B2(new_n280), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1205), .A2(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n1142), .A2(new_n833), .B1(new_n786), .B2(new_n1141), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n821), .A2(G128), .B1(new_n760), .B2(G137), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n772), .B2(new_n1144), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(G150), .C2(new_n1023), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT122), .B(G124), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n840), .C2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT59), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1217), .B1(new_n768), .B2(new_n777), .C1(new_n1213), .C2(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1209), .B1(new_n1206), .B2(new_n1205), .C1(new_n1215), .C2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1199), .B1(new_n1220), .B2(new_n751), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1190), .B2(new_n749), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1198), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1179), .B1(new_n1128), .B2(new_n1178), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1163), .A2(new_n1174), .A3(KEYINPUT118), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1166), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT123), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1181), .A2(KEYINPUT123), .A3(new_n1166), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1197), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT123), .B1(new_n1181), .B2(new_n1166), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1228), .B(new_n1165), .C1(new_n1175), .C2(new_n1180), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1234), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n739), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1224), .B1(new_n1232), .B2(new_n1238), .ZN(G375));
  NOR2_X1   g1039(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n871), .A2(new_n748), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n740), .B1(G68), .B2(new_n1130), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n423), .B1(new_n384), .B2(new_n777), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT125), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1023), .A2(G50), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n827), .A2(G159), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G150), .A2(new_n760), .B1(new_n840), .B2(G128), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT126), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n763), .A2(G132), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1251), .B1(new_n832), .B2(new_n756), .C1(new_n786), .C2(new_n1144), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n764), .A2(G116), .B1(new_n760), .B2(G107), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n788), .B2(new_n833), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT124), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1012), .B1(new_n218), .B2(new_n772), .C1(new_n355), .C2(new_n775), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n326), .B1(new_n767), .B2(new_n791), .C1(new_n756), .C2(new_n782), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n1250), .A2(new_n1252), .B1(new_n1255), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1243), .B1(new_n1259), .B2(new_n751), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1241), .A2(new_n738), .B1(new_n1242), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1240), .A2(new_n1165), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n979), .A3(new_n1174), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(G381));
  NOR2_X1   g1064(.A1(G393), .A2(G396), .ZN(new_n1265));
  INV_X1    g1065(.A(G384), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1267), .A2(G378), .A3(G381), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n696), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1197), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1233), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1223), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1035), .B(G390), .C1(new_n1002), .C2(new_n1008), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1268), .A2(new_n1272), .A3(new_n1273), .ZN(G407));
  INV_X1    g1074(.A(G378), .ZN(new_n1275));
  INV_X1    g1075(.A(G213), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(G343), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1272), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(G407), .A2(new_n1278), .A3(G213), .ZN(G409));
  OAI211_X1 g1079(.A(G378), .B(new_n1224), .C1(new_n1232), .C2(new_n1238), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1197), .B(new_n979), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1275), .B1(new_n1282), .B2(new_n1223), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1277), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1262), .B(KEYINPUT60), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(new_n739), .A3(new_n1174), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1261), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1266), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(G384), .A3(new_n1261), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1284), .A2(new_n1285), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1277), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(new_n1297), .A3(new_n1292), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1277), .A2(G2897), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1289), .A2(new_n1290), .A3(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1299), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(G378), .B1(new_n1224), .B2(new_n1281), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1272), .B2(G378), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1305), .B2(new_n1277), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1294), .A2(new_n1295), .A3(new_n1298), .A4(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G387), .A2(G390), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1009), .A2(new_n1036), .A3(new_n1104), .ZN(new_n1309));
  INV_X1    g1109(.A(G396), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1310), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1265), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1308), .A2(new_n1309), .A3(new_n1312), .ZN(new_n1313));
  OR2_X1    g1113(.A1(new_n1265), .A2(new_n1311), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1104), .B1(new_n1009), .B2(new_n1036), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1314), .B1(new_n1315), .B2(new_n1273), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1307), .A2(new_n1318), .ZN(new_n1319));
  OR2_X1    g1119(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1317), .B(new_n1295), .C1(new_n1296), .C2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT63), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1293), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT127), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1325), .B1(new_n1293), .B2(new_n1323), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1296), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1292), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1322), .A2(new_n1324), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1319), .A2(new_n1328), .ZN(G405));
  NAND2_X1  g1129(.A1(G375), .A2(new_n1275), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1280), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1292), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1330), .A2(new_n1280), .A3(new_n1291), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1334), .B(new_n1318), .ZN(G402));
endmodule


