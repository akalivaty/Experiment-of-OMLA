

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U548 ( .A1(n516), .A2(G2105), .ZN(n613) );
  NOR2_X1 U549 ( .A1(G2104), .A2(G2105), .ZN(n554) );
  NOR2_X2 U550 ( .A1(G1966), .A2(n733), .ZN(n743) );
  XOR2_X1 U551 ( .A(KEYINPUT105), .B(n830), .Z(n831) );
  BUF_X1 U552 ( .A(n609), .Z(n610) );
  XNOR2_X1 U553 ( .A(G2104), .B(KEYINPUT65), .ZN(n516) );
  OR2_X1 U554 ( .A1(n766), .A2(n754), .ZN(n761) );
  NOR2_X2 U555 ( .A1(n727), .A2(n726), .ZN(n729) );
  XNOR2_X1 U556 ( .A(KEYINPUT28), .B(KEYINPUT95), .ZN(n691) );
  NAND2_X1 U557 ( .A1(G171), .A2(n721), .ZN(n719) );
  XNOR2_X1 U558 ( .A(n742), .B(n741), .ZN(n766) );
  NAND2_X1 U559 ( .A1(n740), .A2(G8), .ZN(n742) );
  INV_X1 U560 ( .A(G299), .ZN(n932) );
  AND2_X1 U561 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U562 ( .A1(G543), .A2(G651), .ZN(n639) );
  XOR2_X1 U563 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U564 ( .A1(n693), .A2(n932), .ZN(n692) );
  NOR2_X1 U565 ( .A1(n690), .A2(n689), .ZN(n693) );
  AND2_X1 U566 ( .A1(n571), .A2(n570), .ZN(n517) );
  INV_X1 U567 ( .A(n931), .ZN(n702) );
  NAND2_X1 U568 ( .A1(n703), .A2(n702), .ZN(n704) );
  INV_X1 U569 ( .A(KEYINPUT29), .ZN(n713) );
  INV_X1 U570 ( .A(KEYINPUT31), .ZN(n728) );
  INV_X1 U571 ( .A(KEYINPUT32), .ZN(n741) );
  XOR2_X1 U572 ( .A(G543), .B(KEYINPUT0), .Z(n653) );
  NOR2_X2 U573 ( .A1(G651), .A2(n653), .ZN(n648) );
  NAND2_X1 U574 ( .A1(G52), .A2(n648), .ZN(n520) );
  INV_X1 U575 ( .A(G651), .ZN(n521) );
  NOR2_X1 U576 ( .A1(G543), .A2(n521), .ZN(n518) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n518), .Z(n652) );
  NAND2_X1 U578 ( .A1(G64), .A2(n652), .ZN(n519) );
  NAND2_X1 U579 ( .A1(n520), .A2(n519), .ZN(n527) );
  NOR2_X1 U580 ( .A1(n653), .A2(n521), .ZN(n640) );
  NAND2_X1 U581 ( .A1(G77), .A2(n640), .ZN(n523) );
  NAND2_X1 U582 ( .A1(G90), .A2(n639), .ZN(n522) );
  NAND2_X1 U583 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U584 ( .A(KEYINPUT69), .B(n524), .ZN(n525) );
  XNOR2_X1 U585 ( .A(KEYINPUT9), .B(n525), .ZN(n526) );
  NOR2_X1 U586 ( .A1(n527), .A2(n526), .ZN(G171) );
  NAND2_X1 U587 ( .A1(G78), .A2(n640), .ZN(n529) );
  NAND2_X1 U588 ( .A1(G91), .A2(n639), .ZN(n528) );
  NAND2_X1 U589 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U590 ( .A(KEYINPUT70), .B(n530), .Z(n534) );
  NAND2_X1 U591 ( .A1(G53), .A2(n648), .ZN(n532) );
  NAND2_X1 U592 ( .A1(G65), .A2(n652), .ZN(n531) );
  AND2_X1 U593 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U594 ( .A1(n534), .A2(n533), .ZN(G299) );
  NAND2_X1 U595 ( .A1(n639), .A2(G89), .ZN(n535) );
  XNOR2_X1 U596 ( .A(n535), .B(KEYINPUT4), .ZN(n537) );
  NAND2_X1 U597 ( .A1(G76), .A2(n640), .ZN(n536) );
  NAND2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U599 ( .A(n538), .B(KEYINPUT5), .ZN(n544) );
  XNOR2_X1 U600 ( .A(KEYINPUT75), .B(KEYINPUT6), .ZN(n542) );
  NAND2_X1 U601 ( .A1(G51), .A2(n648), .ZN(n540) );
  NAND2_X1 U602 ( .A1(G63), .A2(n652), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U604 ( .A(n542), .B(n541), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U606 ( .A(KEYINPUT7), .B(n545), .ZN(G168) );
  XNOR2_X2 U607 ( .A(G2104), .B(KEYINPUT65), .ZN(n549) );
  NOR2_X2 U608 ( .A1(n549), .A2(G2105), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n546), .B(KEYINPUT66), .ZN(n567) );
  NAND2_X1 U610 ( .A1(n567), .A2(G101), .ZN(n548) );
  INV_X1 U611 ( .A(KEYINPUT23), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n613), .A2(G125), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n553) );
  INV_X1 U615 ( .A(KEYINPUT67), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n553), .B(n552), .ZN(n559) );
  AND2_X1 U617 ( .A1(G2104), .A2(G2105), .ZN(n892) );
  NAND2_X1 U618 ( .A1(G113), .A2(n892), .ZN(n557) );
  XOR2_X1 U619 ( .A(KEYINPUT17), .B(n554), .Z(n555) );
  XNOR2_X2 U620 ( .A(KEYINPUT68), .B(n555), .ZN(n895) );
  NAND2_X1 U621 ( .A1(G137), .A2(n895), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X2 U623 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(KEYINPUT64), .ZN(n684) );
  BUF_X1 U625 ( .A(n684), .Z(G160) );
  NAND2_X1 U626 ( .A1(G72), .A2(n640), .ZN(n562) );
  NAND2_X1 U627 ( .A1(G85), .A2(n639), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G47), .A2(n648), .ZN(n564) );
  NAND2_X1 U630 ( .A1(G60), .A2(n652), .ZN(n563) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  OR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(G290) );
  AND2_X1 U633 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U634 ( .A(G132), .ZN(G219) );
  INV_X1 U635 ( .A(G82), .ZN(G220) );
  INV_X1 U636 ( .A(G57), .ZN(G237) );
  BUF_X1 U637 ( .A(n567), .Z(n609) );
  NAND2_X1 U638 ( .A1(G102), .A2(n609), .ZN(n568) );
  XNOR2_X1 U639 ( .A(KEYINPUT85), .B(n568), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G138), .A2(n895), .ZN(n572) );
  NAND2_X1 U641 ( .A1(G126), .A2(n613), .ZN(n569) );
  XNOR2_X1 U642 ( .A(n569), .B(KEYINPUT84), .ZN(n571) );
  NAND2_X1 U643 ( .A1(n892), .A2(G114), .ZN(n570) );
  NAND2_X1 U644 ( .A1(n572), .A2(n517), .ZN(n573) );
  NOR2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U646 ( .A(KEYINPUT86), .B(n575), .ZN(G164) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U648 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U649 ( .A(G223), .ZN(n834) );
  NAND2_X1 U650 ( .A1(n834), .A2(G567), .ZN(n577) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  NAND2_X1 U652 ( .A1(n639), .A2(G81), .ZN(n578) );
  XNOR2_X1 U653 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U654 ( .A1(G68), .A2(n640), .ZN(n579) );
  NAND2_X1 U655 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U656 ( .A(n581), .B(KEYINPUT13), .ZN(n583) );
  NAND2_X1 U657 ( .A1(G43), .A2(n648), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n652), .A2(G56), .ZN(n584) );
  XOR2_X1 U660 ( .A(KEYINPUT14), .B(n584), .Z(n585) );
  NOR2_X1 U661 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U662 ( .A(KEYINPUT71), .B(n587), .ZN(n935) );
  INV_X1 U663 ( .A(G860), .ZN(n623) );
  NOR2_X1 U664 ( .A1(n935), .A2(n623), .ZN(n588) );
  XOR2_X1 U665 ( .A(KEYINPUT72), .B(n588), .Z(G153) );
  INV_X1 U666 ( .A(G171), .ZN(G301) );
  NAND2_X1 U667 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G92), .A2(n639), .ZN(n590) );
  NAND2_X1 U669 ( .A1(G66), .A2(n652), .ZN(n589) );
  NAND2_X1 U670 ( .A1(n590), .A2(n589), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n648), .A2(G54), .ZN(n591) );
  XOR2_X1 U672 ( .A(KEYINPUT73), .B(n591), .Z(n593) );
  NAND2_X1 U673 ( .A1(n640), .A2(G79), .ZN(n592) );
  NAND2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U675 ( .A(KEYINPUT74), .B(n594), .ZN(n595) );
  NOR2_X1 U676 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U677 ( .A(n597), .B(KEYINPUT15), .ZN(n931) );
  INV_X1 U678 ( .A(G868), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n931), .A2(n606), .ZN(n598) );
  NAND2_X1 U680 ( .A1(n599), .A2(n598), .ZN(G284) );
  NOR2_X1 U681 ( .A1(G286), .A2(n606), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n600), .B(KEYINPUT76), .ZN(n602) );
  NOR2_X1 U683 ( .A1(G299), .A2(G868), .ZN(n601) );
  NOR2_X1 U684 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U685 ( .A1(n623), .A2(G559), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n603), .A2(n702), .ZN(n604) );
  XNOR2_X1 U687 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  OR2_X1 U688 ( .A1(G559), .A2(n931), .ZN(n605) );
  NAND2_X1 U689 ( .A1(n605), .A2(G868), .ZN(n608) );
  NAND2_X1 U690 ( .A1(n935), .A2(n606), .ZN(n607) );
  NAND2_X1 U691 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U692 ( .A1(G111), .A2(n892), .ZN(n612) );
  NAND2_X1 U693 ( .A1(G99), .A2(n610), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n613), .A2(G123), .ZN(n614) );
  XNOR2_X1 U696 ( .A(n614), .B(KEYINPUT18), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G135), .A2(n895), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U699 ( .A(KEYINPUT77), .B(n617), .Z(n618) );
  NOR2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n1000) );
  XNOR2_X1 U701 ( .A(n1000), .B(G2096), .ZN(n621) );
  INV_X1 U702 ( .A(G2100), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n621), .A2(n620), .ZN(G156) );
  NAND2_X1 U704 ( .A1(G559), .A2(n702), .ZN(n622) );
  XOR2_X1 U705 ( .A(n935), .B(n622), .Z(n662) );
  NAND2_X1 U706 ( .A1(n623), .A2(n662), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G55), .A2(n648), .ZN(n625) );
  NAND2_X1 U708 ( .A1(G67), .A2(n652), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G80), .A2(n640), .ZN(n627) );
  NAND2_X1 U711 ( .A1(G93), .A2(n639), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n664) );
  XOR2_X1 U714 ( .A(n630), .B(n664), .Z(G145) );
  NAND2_X1 U715 ( .A1(n639), .A2(G86), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G48), .A2(n648), .ZN(n632) );
  NAND2_X1 U717 ( .A1(G61), .A2(n652), .ZN(n631) );
  NAND2_X1 U718 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U719 ( .A1(G73), .A2(n640), .ZN(n633) );
  XOR2_X1 U720 ( .A(KEYINPUT2), .B(n633), .Z(n634) );
  NOR2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U723 ( .A(n638), .B(KEYINPUT78), .ZN(G305) );
  NAND2_X1 U724 ( .A1(n639), .A2(G88), .ZN(n643) );
  NAND2_X1 U725 ( .A1(G75), .A2(n640), .ZN(n641) );
  XOR2_X1 U726 ( .A(KEYINPUT79), .B(n641), .Z(n642) );
  NAND2_X1 U727 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U728 ( .A1(G50), .A2(n648), .ZN(n645) );
  NAND2_X1 U729 ( .A1(G62), .A2(n652), .ZN(n644) );
  NAND2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U731 ( .A1(n647), .A2(n646), .ZN(G166) );
  NAND2_X1 U732 ( .A1(G49), .A2(n648), .ZN(n650) );
  NAND2_X1 U733 ( .A1(G74), .A2(G651), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U735 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U736 ( .A1(n653), .A2(G87), .ZN(n654) );
  NAND2_X1 U737 ( .A1(n655), .A2(n654), .ZN(G288) );
  XNOR2_X1 U738 ( .A(n932), .B(G166), .ZN(n658) );
  XOR2_X1 U739 ( .A(KEYINPUT19), .B(KEYINPUT80), .Z(n656) );
  XNOR2_X1 U740 ( .A(G290), .B(n656), .ZN(n657) );
  XNOR2_X1 U741 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U742 ( .A(n664), .B(n659), .ZN(n660) );
  XNOR2_X1 U743 ( .A(n660), .B(G288), .ZN(n661) );
  XNOR2_X1 U744 ( .A(G305), .B(n661), .ZN(n912) );
  XNOR2_X1 U745 ( .A(n662), .B(n912), .ZN(n663) );
  NAND2_X1 U746 ( .A1(n663), .A2(G868), .ZN(n666) );
  OR2_X1 U747 ( .A1(G868), .A2(n664), .ZN(n665) );
  NAND2_X1 U748 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U753 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XOR2_X1 U754 ( .A(KEYINPUT81), .B(G44), .Z(n671) );
  XNOR2_X1 U755 ( .A(KEYINPUT3), .B(n671), .ZN(G218) );
  NAND2_X1 U756 ( .A1(G120), .A2(G69), .ZN(n672) );
  NOR2_X1 U757 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U758 ( .A1(G108), .A2(n673), .ZN(n839) );
  NAND2_X1 U759 ( .A1(G567), .A2(n839), .ZN(n674) );
  XNOR2_X1 U760 ( .A(KEYINPUT83), .B(n674), .ZN(n680) );
  NOR2_X1 U761 ( .A1(G220), .A2(G219), .ZN(n675) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(n675), .Z(n676) );
  NOR2_X1 U763 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U764 ( .A1(G96), .A2(n677), .ZN(n838) );
  NAND2_X1 U765 ( .A1(G2106), .A2(n838), .ZN(n678) );
  XOR2_X1 U766 ( .A(KEYINPUT82), .B(n678), .Z(n679) );
  NOR2_X1 U767 ( .A1(n680), .A2(n679), .ZN(G319) );
  INV_X1 U768 ( .A(G319), .ZN(n682) );
  NAND2_X1 U769 ( .A1(G661), .A2(G483), .ZN(n681) );
  NOR2_X1 U770 ( .A1(n682), .A2(n681), .ZN(n837) );
  NAND2_X1 U771 ( .A1(n837), .A2(G36), .ZN(G176) );
  XNOR2_X1 U772 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  XNOR2_X1 U773 ( .A(G1981), .B(G305), .ZN(n683) );
  XNOR2_X1 U774 ( .A(n683), .B(KEYINPUT98), .ZN(n943) );
  NAND2_X1 U775 ( .A1(n684), .A2(G40), .ZN(n781) );
  INV_X1 U776 ( .A(KEYINPUT92), .ZN(n685) );
  XNOR2_X1 U777 ( .A(n781), .B(n685), .ZN(n686) );
  NOR2_X1 U778 ( .A1(G1384), .A2(G164), .ZN(n783) );
  NAND2_X2 U779 ( .A1(n686), .A2(n783), .ZN(n722) );
  INV_X1 U780 ( .A(n722), .ZN(n687) );
  NAND2_X1 U781 ( .A1(n687), .A2(G2072), .ZN(n688) );
  XNOR2_X1 U782 ( .A(n688), .B(KEYINPUT27), .ZN(n690) );
  BUF_X2 U783 ( .A(n722), .Z(n734) );
  AND2_X2 U784 ( .A1(G1956), .A2(n734), .ZN(n689) );
  XNOR2_X1 U785 ( .A(n692), .B(n691), .ZN(n712) );
  BUF_X1 U786 ( .A(n693), .Z(n694) );
  NAND2_X1 U787 ( .A1(n694), .A2(n932), .ZN(n710) );
  INV_X1 U788 ( .A(G1996), .ZN(n695) );
  NOR2_X1 U789 ( .A1(n722), .A2(n695), .ZN(n696) );
  XOR2_X1 U790 ( .A(n696), .B(KEYINPUT26), .Z(n699) );
  AND2_X1 U791 ( .A1(n734), .A2(G1341), .ZN(n697) );
  NOR2_X1 U792 ( .A1(n697), .A2(n935), .ZN(n698) );
  NAND2_X1 U793 ( .A1(n699), .A2(n698), .ZN(n705) );
  NAND2_X1 U794 ( .A1(G1348), .A2(n734), .ZN(n701) );
  INV_X1 U795 ( .A(n722), .ZN(n716) );
  NAND2_X1 U796 ( .A1(G2067), .A2(n716), .ZN(n700) );
  NAND2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n706) );
  INV_X1 U798 ( .A(n706), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n705), .A2(n704), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n931), .A2(n706), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U803 ( .A1(n712), .A2(n711), .ZN(n714) );
  XNOR2_X1 U804 ( .A(n714), .B(n713), .ZN(n720) );
  XNOR2_X1 U805 ( .A(G1961), .B(KEYINPUT93), .ZN(n961) );
  NAND2_X1 U806 ( .A1(n734), .A2(n961), .ZN(n715) );
  XNOR2_X1 U807 ( .A(n715), .B(KEYINPUT94), .ZN(n718) );
  XNOR2_X1 U808 ( .A(KEYINPUT25), .B(G2078), .ZN(n985) );
  NAND2_X1 U809 ( .A1(n716), .A2(n985), .ZN(n717) );
  NAND2_X1 U810 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U811 ( .A1(n720), .A2(n719), .ZN(n731) );
  NOR2_X1 U812 ( .A1(G171), .A2(n721), .ZN(n727) );
  NAND2_X1 U813 ( .A1(G8), .A2(n722), .ZN(n733) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n722), .ZN(n745) );
  NOR2_X1 U815 ( .A1(n743), .A2(n745), .ZN(n723) );
  NAND2_X1 U816 ( .A1(n723), .A2(G8), .ZN(n724) );
  XNOR2_X1 U817 ( .A(n724), .B(KEYINPUT30), .ZN(n725) );
  NOR2_X1 U818 ( .A1(G168), .A2(n725), .ZN(n726) );
  XNOR2_X1 U819 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n744) );
  NAND2_X1 U821 ( .A1(n744), .A2(G286), .ZN(n732) );
  XNOR2_X1 U822 ( .A(n732), .B(KEYINPUT96), .ZN(n739) );
  BUF_X1 U823 ( .A(n733), .Z(n750) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n750), .ZN(n736) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n734), .ZN(n735) );
  NOR2_X1 U826 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U827 ( .A1(n737), .A2(G303), .ZN(n738) );
  NAND2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n740) );
  BUF_X1 U829 ( .A(n744), .Z(n747) );
  NAND2_X1 U830 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U831 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U832 ( .A1(n743), .A2(n748), .ZN(n765) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n756) );
  INV_X1 U834 ( .A(n750), .ZN(n775) );
  NAND2_X1 U835 ( .A1(n756), .A2(n775), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n749), .A2(KEYINPUT33), .ZN(n757) );
  INV_X1 U837 ( .A(n757), .ZN(n753) );
  NOR2_X1 U838 ( .A1(n750), .A2(KEYINPUT33), .ZN(n751) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n928) );
  AND2_X1 U840 ( .A1(n751), .A2(n928), .ZN(n752) );
  NOR2_X1 U841 ( .A1(n753), .A2(n752), .ZN(n759) );
  OR2_X1 U842 ( .A1(n765), .A2(n759), .ZN(n754) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n924) );
  AND2_X1 U845 ( .A1(n924), .A2(n757), .ZN(n758) );
  OR2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U848 ( .A(n762), .B(KEYINPUT97), .ZN(n763) );
  NOR2_X1 U849 ( .A1(n943), .A2(n763), .ZN(n764) );
  XNOR2_X1 U850 ( .A(n764), .B(KEYINPUT99), .ZN(n779) );
  NOR2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n770) );
  NOR2_X1 U852 ( .A1(G2090), .A2(G303), .ZN(n767) );
  NAND2_X1 U853 ( .A1(G8), .A2(n767), .ZN(n768) );
  XOR2_X1 U854 ( .A(KEYINPUT100), .B(n768), .Z(n769) );
  NOR2_X1 U855 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U856 ( .A1(n775), .A2(n771), .ZN(n772) );
  XNOR2_X1 U857 ( .A(n772), .B(KEYINPUT101), .ZN(n777) );
  NOR2_X1 U858 ( .A1(G1981), .A2(G305), .ZN(n773) );
  XNOR2_X1 U859 ( .A(n773), .B(KEYINPUT24), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U863 ( .A(n780), .B(KEYINPUT102), .ZN(n816) );
  BUF_X1 U864 ( .A(n781), .Z(n782) );
  NOR2_X1 U865 ( .A1(n783), .A2(n782), .ZN(n829) );
  NAND2_X1 U866 ( .A1(G104), .A2(n610), .ZN(n785) );
  NAND2_X1 U867 ( .A1(G140), .A2(n895), .ZN(n784) );
  NAND2_X1 U868 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U869 ( .A(KEYINPUT34), .B(n786), .ZN(n791) );
  NAND2_X1 U870 ( .A1(G116), .A2(n892), .ZN(n788) );
  NAND2_X1 U871 ( .A1(G128), .A2(n613), .ZN(n787) );
  NAND2_X1 U872 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U873 ( .A(KEYINPUT35), .B(n789), .Z(n790) );
  NOR2_X1 U874 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U875 ( .A(KEYINPUT36), .B(n792), .ZN(n904) );
  XNOR2_X1 U876 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NOR2_X1 U877 ( .A1(n904), .A2(n826), .ZN(n1003) );
  NAND2_X1 U878 ( .A1(n829), .A2(n1003), .ZN(n824) );
  NAND2_X1 U879 ( .A1(G117), .A2(n892), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G129), .A2(n613), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U882 ( .A(n795), .B(KEYINPUT89), .ZN(n797) );
  NAND2_X1 U883 ( .A1(G141), .A2(n895), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n610), .A2(G105), .ZN(n798) );
  XOR2_X1 U886 ( .A(KEYINPUT38), .B(n798), .Z(n799) );
  NOR2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U888 ( .A(KEYINPUT90), .B(n801), .Z(n908) );
  NAND2_X1 U889 ( .A1(G1996), .A2(n908), .ZN(n810) );
  NAND2_X1 U890 ( .A1(n610), .A2(G95), .ZN(n806) );
  NAND2_X1 U891 ( .A1(G107), .A2(n892), .ZN(n803) );
  NAND2_X1 U892 ( .A1(G119), .A2(n613), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U894 ( .A(KEYINPUT88), .B(n804), .Z(n805) );
  AND2_X1 U895 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U896 ( .A1(G131), .A2(n895), .ZN(n807) );
  NAND2_X1 U897 ( .A1(n808), .A2(n807), .ZN(n889) );
  NAND2_X1 U898 ( .A1(G1991), .A2(n889), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n1007) );
  NAND2_X1 U900 ( .A1(n829), .A2(n1007), .ZN(n811) );
  XNOR2_X1 U901 ( .A(KEYINPUT91), .B(n811), .ZN(n821) );
  INV_X1 U902 ( .A(n821), .ZN(n812) );
  AND2_X1 U903 ( .A1(n824), .A2(n812), .ZN(n814) );
  XNOR2_X1 U904 ( .A(G1986), .B(G290), .ZN(n927) );
  NAND2_X1 U905 ( .A1(n927), .A2(n829), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n832) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n908), .ZN(n817) );
  XOR2_X1 U908 ( .A(KEYINPUT103), .B(n817), .Z(n998) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n889), .ZN(n1001) );
  NOR2_X1 U911 ( .A1(n818), .A2(n1001), .ZN(n819) );
  XNOR2_X1 U912 ( .A(n819), .B(KEYINPUT104), .ZN(n820) );
  NOR2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U914 ( .A1(n998), .A2(n822), .ZN(n823) );
  XNOR2_X1 U915 ( .A(KEYINPUT39), .B(n823), .ZN(n825) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n904), .A2(n826), .ZN(n1012) );
  NAND2_X1 U918 ( .A1(n827), .A2(n1012), .ZN(n828) );
  NAND2_X1 U919 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U920 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U921 ( .A(KEYINPUT40), .B(n833), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U924 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U926 ( .A1(n837), .A2(n836), .ZN(G188) );
  XOR2_X1 U927 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  NOR2_X1 U931 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U933 ( .A(KEYINPUT106), .B(G2446), .ZN(n849) );
  XOR2_X1 U934 ( .A(G2430), .B(G2427), .Z(n841) );
  XNOR2_X1 U935 ( .A(G2435), .B(G2438), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U937 ( .A(G2454), .B(KEYINPUT107), .Z(n843) );
  XNOR2_X1 U938 ( .A(G1341), .B(G1348), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U940 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U941 ( .A(G2451), .B(G2443), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U943 ( .A(n849), .B(n848), .ZN(n850) );
  NAND2_X1 U944 ( .A1(n850), .A2(G14), .ZN(n851) );
  XNOR2_X1 U945 ( .A(KEYINPUT108), .B(n851), .ZN(n918) );
  XNOR2_X1 U946 ( .A(n918), .B(KEYINPUT109), .ZN(G401) );
  XOR2_X1 U947 ( .A(G2100), .B(G2096), .Z(n853) );
  XNOR2_X1 U948 ( .A(KEYINPUT42), .B(G2678), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U950 ( .A(KEYINPUT43), .B(G2090), .Z(n855) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U953 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U954 ( .A(G2078), .B(G2084), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n859), .B(n858), .ZN(G227) );
  XOR2_X1 U956 ( .A(G1986), .B(G1971), .Z(n861) );
  XNOR2_X1 U957 ( .A(G1981), .B(G1966), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(n871) );
  XOR2_X1 U959 ( .A(KEYINPUT112), .B(G2474), .Z(n863) );
  XNOR2_X1 U960 ( .A(G1996), .B(KEYINPUT111), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U962 ( .A(G1976), .B(G1956), .Z(n865) );
  XNOR2_X1 U963 ( .A(G1991), .B(G1961), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U965 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U966 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U968 ( .A(n871), .B(n870), .Z(G229) );
  NAND2_X1 U969 ( .A1(G136), .A2(n895), .ZN(n872) );
  XNOR2_X1 U970 ( .A(KEYINPUT114), .B(n872), .ZN(n875) );
  NAND2_X1 U971 ( .A1(n613), .A2(G124), .ZN(n873) );
  XNOR2_X1 U972 ( .A(KEYINPUT44), .B(n873), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n876), .B(KEYINPUT115), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G100), .A2(n610), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n892), .A2(G112), .ZN(n879) );
  XOR2_X1 U978 ( .A(KEYINPUT116), .B(n879), .Z(n880) );
  NOR2_X1 U979 ( .A1(n881), .A2(n880), .ZN(G162) );
  XNOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n891) );
  NAND2_X1 U981 ( .A1(G103), .A2(n610), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G139), .A2(n895), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G115), .A2(n892), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G127), .A2(n613), .ZN(n884) );
  NAND2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U987 ( .A(KEYINPUT47), .B(n886), .Z(n887) );
  NOR2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n1015) );
  XNOR2_X1 U989 ( .A(n889), .B(n1015), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n902) );
  NAND2_X1 U991 ( .A1(G118), .A2(n892), .ZN(n894) );
  NAND2_X1 U992 ( .A1(G130), .A2(n613), .ZN(n893) );
  NAND2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n900) );
  NAND2_X1 U994 ( .A1(G106), .A2(n610), .ZN(n897) );
  NAND2_X1 U995 ( .A1(G142), .A2(n895), .ZN(n896) );
  NAND2_X1 U996 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(n898), .B(KEYINPUT45), .Z(n899) );
  NOR2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U999 ( .A(n902), .B(n901), .Z(n903) );
  XNOR2_X1 U1000 ( .A(G162), .B(n903), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n904), .B(n1000), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1003 ( .A(n908), .B(n907), .Z(n909) );
  XNOR2_X1 U1004 ( .A(G164), .B(n909), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n910), .B(G160), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n911), .ZN(G395) );
  XNOR2_X1 U1007 ( .A(G286), .B(n912), .ZN(n915) );
  XNOR2_X1 U1008 ( .A(KEYINPUT117), .B(G301), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(n913), .B(n935), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1011 ( .A(n916), .B(n931), .Z(n917) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n917), .ZN(G397) );
  NAND2_X1 U1013 ( .A1(n918), .A2(G319), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n919), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1021 ( .A(KEYINPUT56), .B(G16), .ZN(n948) );
  XNOR2_X1 U1022 ( .A(G171), .B(G1961), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n929) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n941) );
  XOR2_X1 U1026 ( .A(G1348), .B(KEYINPUT122), .Z(n930) );
  XNOR2_X1 U1027 ( .A(n931), .B(n930), .ZN(n939) );
  XNOR2_X1 U1028 ( .A(n932), .B(G1956), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(G1971), .A2(G303), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(G1341), .B(n935), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n946) );
  XOR2_X1 U1035 ( .A(G168), .B(G1966), .Z(n942) );
  NOR2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1037 ( .A(KEYINPUT57), .B(n944), .Z(n945) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1039 ( .A1(n948), .A2(n947), .ZN(n1030) );
  XOR2_X1 U1040 ( .A(G1341), .B(G19), .Z(n951) );
  XNOR2_X1 U1041 ( .A(G20), .B(KEYINPUT123), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(n949), .B(G1956), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(G6), .B(G1981), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1046 ( .A(KEYINPUT124), .B(n954), .Z(n958) );
  XNOR2_X1 U1047 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(n955), .B(G4), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G1348), .B(n956), .ZN(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(KEYINPUT60), .B(n959), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(n960), .B(KEYINPUT126), .ZN(n972) );
  XOR2_X1 U1053 ( .A(G1966), .B(G21), .Z(n963) );
  XNOR2_X1 U1054 ( .A(n961), .B(G5), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n970) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G22), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(G23), .B(G1976), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n967) );
  XOR2_X1 U1059 ( .A(G1986), .B(G24), .Z(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT58), .B(n968), .ZN(n969) );
  NOR2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n974), .B(n973), .ZN(n976) );
  INV_X1 U1066 ( .A(G16), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n977), .A2(G11), .ZN(n1028) );
  XNOR2_X1 U1069 ( .A(G2090), .B(G35), .ZN(n990) );
  XNOR2_X1 U1070 ( .A(G1996), .B(G32), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(G33), .B(G2072), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n984) );
  XOR2_X1 U1073 ( .A(G1991), .B(G25), .Z(n980) );
  NAND2_X1 U1074 ( .A1(n980), .A2(G28), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(G26), .B(G2067), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1078 ( .A(G27), .B(n985), .Z(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT53), .B(n988), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1082 ( .A(G2084), .B(KEYINPUT54), .Z(n991) );
  XNOR2_X1 U1083 ( .A(G34), .B(n991), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(KEYINPUT55), .B(n994), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(G29), .A2(n995), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n996), .B(KEYINPUT121), .ZN(n1026) );
  XOR2_X1 U1088 ( .A(G2090), .B(G162), .Z(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1090 ( .A(KEYINPUT51), .B(n999), .Z(n1010) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1005) );
  XOR2_X1 U1092 ( .A(G2084), .B(G160), .Z(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(KEYINPUT118), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(n1011), .B(KEYINPUT119), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(KEYINPUT120), .B(n1014), .ZN(n1020) );
  XOR2_X1 U1101 ( .A(G2072), .B(n1015), .Z(n1017) );
  XOR2_X1 U1102 ( .A(G164), .B(G2078), .Z(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(KEYINPUT50), .B(n1018), .Z(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1021), .B(KEYINPUT52), .ZN(n1023) );
  INV_X1 U1107 ( .A(KEYINPUT55), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(G29), .A2(n1024), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1112 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

