//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  AOI22_X1  g003(.A1(new_n203), .A2(new_n204), .B1(G211gat), .B2(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n203), .B2(new_n204), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G226gat), .A2(G233gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT64), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n214), .B1(G169gat), .B2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT26), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n216), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT65), .B1(new_n225), .B2(new_n212), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n217), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT27), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT27), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G183gat), .ZN(new_n231));
  INV_X1    g030(.A(G190gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT28), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT27), .B(G183gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT28), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n236), .A3(new_n232), .ZN(new_n237));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n234), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n240), .A2(new_n241), .B1(G169gat), .B2(G176gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n228), .A2(new_n232), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(KEYINPUT24), .A3(new_n238), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n223), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n242), .A2(new_n244), .A3(new_n245), .A4(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n218), .B1(new_n238), .B2(KEYINPUT24), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT23), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n244), .A4(new_n254), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n227), .A2(new_n239), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n211), .B1(new_n256), .B2(KEYINPUT29), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n250), .A2(new_n255), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n240), .B1(new_n233), .B2(KEYINPUT28), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n227), .A2(new_n259), .A3(new_n237), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n211), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT74), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT74), .ZN(new_n264));
  AOI211_X1 g063(.A(new_n264), .B(new_n211), .C1(new_n258), .C2(new_n260), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n210), .B(new_n257), .C1(new_n263), .C2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n210), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT29), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n262), .B1(new_n261), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n256), .A2(new_n211), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G8gat), .B(G36gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(G64gat), .B(G92gat), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  AND3_X1   g073(.A1(new_n266), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n274), .B1(new_n266), .B2(new_n271), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AND4_X1   g077(.A1(new_n277), .A2(new_n266), .A3(new_n271), .A4(new_n274), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n202), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n276), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n271), .A3(new_n274), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(KEYINPUT30), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n279), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT83), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G228gat), .A2(G233gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n288));
  INV_X1    g087(.A(G148gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(G141gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(G141gat), .ZN(new_n291));
  INV_X1    g090(.A(G141gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n292), .A2(KEYINPUT75), .A3(G148gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n297));
  INV_X1    g096(.A(G162gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT2), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(G155gat), .ZN(new_n300));
  INV_X1    g099(.A(G155gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G162gat), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n290), .A2(new_n293), .A3(KEYINPUT76), .A4(new_n291), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n296), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307));
  INV_X1    g106(.A(new_n291), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n289), .A2(G141gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n300), .A2(new_n302), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n305), .A2(new_n306), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n210), .B1(new_n268), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n287), .B1(new_n314), .B2(KEYINPUT80), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G22gat), .ZN(new_n316));
  INV_X1    g115(.A(G22gat), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n317), .B(new_n287), .C1(new_n314), .C2(KEYINPUT80), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n306), .B1(new_n267), .B2(KEYINPUT29), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n312), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n314), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G78gat), .B(G106gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(G50gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(KEYINPUT81), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n320), .A2(new_n321), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n268), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n267), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n332), .A3(new_n318), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n323), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n327), .B(KEYINPUT81), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n323), .B2(new_n333), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G120gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G113gat), .ZN(new_n339));
  INV_X1    g138(.A(G113gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G120gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G127gat), .B(G134gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT68), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT1), .B1(new_n339), .B2(new_n341), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT68), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n343), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G134gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G127gat), .ZN(new_n352));
  INV_X1    g151(.A(G127gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G134gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT66), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n358), .A2(KEYINPUT67), .A3(new_n347), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT67), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n353), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n343), .B2(new_n355), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n344), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n350), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(new_n258), .A3(new_n260), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT67), .B1(new_n358), .B2(new_n347), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n363), .A2(new_n360), .A3(new_n356), .A4(new_n357), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n367), .A2(new_n368), .B1(new_n346), .B2(new_n349), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n254), .A2(KEYINPUT25), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n242), .A2(new_n244), .A3(new_n247), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n370), .A2(new_n371), .B1(new_n248), .B2(new_n249), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n227), .A2(new_n259), .A3(new_n237), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n366), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT32), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT33), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT69), .ZN(new_n382));
  INV_X1    g181(.A(G15gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G43gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n378), .A2(new_n380), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n384), .B(G43gat), .ZN(new_n388));
  OAI211_X1 g187(.A(KEYINPUT32), .B(new_n377), .C1(new_n388), .C2(new_n379), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT72), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT71), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n256), .A2(new_n365), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n369), .A2(new_n372), .A3(new_n373), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n375), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT70), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n376), .B1(new_n366), .B2(new_n374), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n398), .A2(KEYINPUT70), .A3(KEYINPUT71), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT34), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n395), .A2(new_n396), .A3(new_n392), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT71), .B1(new_n398), .B2(KEYINPUT70), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT34), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n390), .A2(new_n391), .A3(new_n400), .A4(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n391), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n403), .B1(new_n401), .B2(new_n402), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n391), .B1(new_n387), .B2(new_n389), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n286), .A2(new_n337), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n294), .B2(new_n295), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n419), .A2(new_n304), .B1(new_n310), .B2(new_n311), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n369), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(new_n365), .A3(new_n313), .ZN(new_n425));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n369), .A2(new_n420), .A3(KEYINPUT4), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n423), .A2(new_n425), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n365), .A2(new_n321), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n421), .ZN(new_n430));
  INV_X1    g229(.A(new_n426), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(KEYINPUT5), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n427), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT4), .B1(new_n369), .B2(new_n420), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT5), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n426), .A4(new_n425), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(new_n438), .A3(KEYINPUT84), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT84), .B1(new_n433), .B2(new_n438), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n417), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n433), .A2(new_n438), .A3(new_n416), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n416), .B1(new_n433), .B2(new_n438), .ZN(new_n448));
  INV_X1    g247(.A(new_n444), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT35), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n412), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n445), .B2(new_n448), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n283), .A2(new_n284), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n411), .A2(new_n337), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT82), .B1(new_n334), .B2(new_n336), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n454), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n323), .A2(new_n333), .ZN(new_n460));
  INV_X1    g259(.A(new_n335), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n323), .A2(new_n328), .A3(new_n333), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n458), .A2(new_n459), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n411), .A2(KEYINPUT36), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n400), .A2(new_n404), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n387), .A2(new_n389), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT72), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n406), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT36), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n405), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n423), .A2(new_n425), .A3(new_n427), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT39), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n431), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n479), .A2(new_n416), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n426), .B1(new_n436), .B2(new_n425), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT39), .B1(new_n430), .B2(new_n431), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n480), .B(KEYINPUT40), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT40), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n481), .A2(new_n482), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n479), .A2(new_n416), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n442), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n337), .B1(new_n286), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n266), .A2(new_n271), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT37), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n274), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n261), .A2(new_n262), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n257), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(new_n494), .B2(new_n210), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n267), .B(new_n257), .C1(new_n263), .C2(new_n265), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT38), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n275), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n433), .A2(new_n438), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n416), .B1(new_n501), .B2(new_n439), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n498), .B(new_n450), .C1(new_n502), .C2(new_n445), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n492), .B1(new_n491), .B2(new_n490), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n503), .A2(KEYINPUT85), .B1(KEYINPUT38), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT85), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n447), .A2(new_n506), .A3(new_n450), .A4(new_n498), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n489), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n457), .B1(new_n476), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(G197gat), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT11), .B(G169gat), .Z(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT12), .Z(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n317), .A2(G15gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n383), .A2(G22gat), .ZN(new_n517));
  INV_X1    g316(.A(G1gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT16), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT87), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n516), .A2(new_n517), .ZN(new_n524));
  AOI21_X1  g323(.A(G8gat), .B1(new_n524), .B2(new_n518), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n526), .A2(KEYINPUT88), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(KEYINPUT88), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n524), .A2(new_n518), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(new_n520), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G43gat), .B(G50gat), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n537));
  NOR2_X1   g336(.A1(G29gat), .A2(G36gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT14), .ZN(new_n539));
  INV_X1    g338(.A(G29gat), .ZN(new_n540));
  INV_X1    g339(.A(G36gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OR4_X1    g341(.A1(new_n536), .A2(new_n537), .A3(new_n539), .A4(new_n542), .ZN(new_n543));
  OAI22_X1  g342(.A1(new_n539), .A2(KEYINPUT86), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n539), .A2(KEYINPUT86), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n536), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n534), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n532), .B1(new_n527), .B2(new_n528), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n543), .A2(new_n546), .A3(KEYINPUT17), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n548), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT18), .B1(new_n555), .B2(KEYINPUT89), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT89), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n548), .A2(new_n553), .A3(new_n557), .A4(new_n554), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n549), .B1(new_n546), .B2(new_n543), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n534), .A2(new_n547), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n554), .B(KEYINPUT13), .Z(new_n562));
  AOI22_X1  g361(.A1(new_n556), .A2(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n548), .A2(new_n553), .A3(KEYINPUT18), .A4(new_n554), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT90), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n515), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n515), .A3(new_n566), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n509), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G64gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(G57gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT91), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(G57gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  OR2_X1    g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n575), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT9), .B1(new_n584), .B2(new_n573), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(new_n579), .A3(new_n580), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G127gat), .B(G155gat), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT20), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n591), .B(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G183gat), .B(G211gat), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n594), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n587), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n534), .B1(KEYINPUT21), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n594), .A2(new_n596), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n594), .A2(new_n596), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G99gat), .B(G106gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(KEYINPUT8), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT94), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT7), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n608), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(new_n608), .A3(new_n616), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(KEYINPUT95), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(KEYINPUT95), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n617), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n547), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n551), .A2(new_n552), .A3(new_n622), .A4(new_n620), .ZN(new_n625));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT96), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n624), .A2(new_n625), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT97), .ZN(new_n631));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n627), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n630), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n607), .A2(KEYINPUT98), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT98), .B1(new_n607), .B2(new_n642), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n620), .A2(new_n622), .A3(new_n587), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n598), .A2(new_n618), .A3(new_n619), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT99), .B(KEYINPUT10), .Z(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n598), .A2(KEYINPUT10), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n623), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n645), .A2(new_n646), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n653), .B1(new_n654), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n655), .A2(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n643), .A2(new_n644), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n571), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n453), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(new_n518), .ZN(G1324gat));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  INV_X1    g469(.A(new_n286), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n571), .A2(new_n671), .A3(new_n666), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT16), .B(G8gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT100), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n670), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n675), .A2(KEYINPUT101), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(KEYINPUT101), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n672), .A2(G8gat), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n672), .A2(new_n670), .A3(new_n673), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT102), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT103), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n678), .A2(new_n684), .A3(new_n679), .A4(new_n681), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(G1325gat));
  INV_X1    g485(.A(new_n411), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n383), .B1(new_n667), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT104), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n472), .A2(new_n473), .A3(new_n405), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n473), .B1(new_n472), .B2(new_n405), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n468), .A2(KEYINPUT105), .A3(new_n474), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n667), .A2(new_n383), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n689), .A2(new_n696), .ZN(G1326gat));
  AND2_X1   g496(.A1(new_n458), .A2(new_n465), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n571), .A2(new_n698), .A3(new_n666), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(new_n607), .ZN(new_n702));
  INV_X1    g501(.A(new_n642), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n702), .A2(new_n703), .A3(new_n663), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n571), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(G29gat), .A3(new_n453), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT45), .Z(new_n707));
  AOI22_X1  g506(.A1(new_n412), .A2(new_n451), .B1(new_n455), .B2(KEYINPUT35), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n466), .B1(new_n693), .B2(new_n694), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n503), .A2(KEYINPUT85), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n504), .A2(KEYINPUT38), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n507), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n489), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n708), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n642), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n640), .A2(KEYINPUT108), .A3(new_n641), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n715), .A2(new_n716), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n509), .B2(new_n642), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n663), .B(KEYINPUT106), .Z(new_n727));
  INV_X1    g526(.A(new_n569), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n567), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n727), .A2(new_n729), .A3(new_n702), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G29gat), .B1(new_n731), .B2(new_n453), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n707), .A2(new_n732), .ZN(G1328gat));
  NOR3_X1   g532(.A1(new_n705), .A2(G36gat), .A3(new_n286), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT46), .ZN(new_n735));
  INV_X1    g534(.A(new_n731), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n671), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n738), .B2(new_n541), .ZN(G1329gat));
  NAND2_X1  g538(.A1(new_n411), .A2(new_n385), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n705), .A2(new_n740), .B1(new_n741), .B2(KEYINPUT47), .ZN(new_n742));
  INV_X1    g541(.A(new_n695), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n742), .B1(new_n744), .B2(G43gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(KEYINPUT47), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n745), .B(new_n746), .Z(G1330gat));
  OAI21_X1  g546(.A(G50gat), .B1(new_n731), .B2(new_n337), .ZN(new_n748));
  INV_X1    g547(.A(new_n698), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n705), .A2(G50gat), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n748), .A2(KEYINPUT48), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n698), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n750), .B1(new_n753), .B2(G50gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n754), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g554(.A1(new_n727), .A2(new_n643), .A3(new_n729), .A4(new_n644), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n715), .ZN(new_n757));
  INV_X1    g556(.A(new_n453), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g559(.A(new_n286), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT110), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n763), .B(new_n764), .Z(G1333gat));
  NAND2_X1  g564(.A1(new_n757), .A2(new_n743), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n687), .A2(G71gat), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n766), .A2(G71gat), .B1(new_n757), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n757), .A2(new_n698), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n702), .A2(new_n570), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n664), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n726), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G85gat), .B1(new_n775), .B2(new_n453), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n772), .A2(new_n642), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n709), .A2(new_n714), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n457), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(KEYINPUT51), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT111), .B1(new_n779), .B2(KEYINPUT51), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n715), .A2(new_n782), .A3(new_n783), .A4(new_n777), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT112), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n691), .A2(new_n692), .A3(new_n690), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT105), .B1(new_n468), .B2(new_n474), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n467), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n457), .B1(new_n788), .B2(new_n508), .ZN(new_n789));
  INV_X1    g588(.A(new_n777), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n782), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n779), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n780), .B1(new_n785), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n663), .A2(new_n758), .A3(new_n610), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n776), .B1(new_n796), .B2(new_n797), .ZN(G1336gat));
  INV_X1    g597(.A(new_n780), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n781), .A2(new_n784), .A3(KEYINPUT112), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n793), .B1(new_n792), .B2(new_n794), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  INV_X1    g602(.A(new_n727), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n804), .A2(G92gat), .A3(new_n286), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n805), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT113), .B1(new_n796), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n726), .A2(new_n809), .A3(new_n671), .A4(new_n774), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n671), .B(new_n774), .C1(new_n722), .C2(new_n724), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n611), .B1(new_n811), .B2(KEYINPUT114), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n806), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n780), .B1(new_n792), .B2(new_n794), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n807), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n811), .A2(G92gat), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT52), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n814), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(G1337gat));
  OAI21_X1  g622(.A(G99gat), .B1(new_n775), .B2(new_n695), .ZN(new_n824));
  OR3_X1    g623(.A1(new_n664), .A2(G99gat), .A3(new_n687), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n796), .B2(new_n825), .ZN(G1338gat));
  INV_X1    g625(.A(G106gat), .ZN(new_n827));
  INV_X1    g626(.A(new_n775), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n698), .ZN(new_n829));
  INV_X1    g628(.A(new_n337), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n727), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT53), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n827), .B1(new_n828), .B2(new_n830), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n796), .A2(new_n831), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(G1339gat));
  NOR3_X1   g636(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n554), .B1(new_n548), .B2(new_n553), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n513), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT117), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n663), .A2(new_n569), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n652), .B1(new_n623), .B2(new_n649), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n648), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n653), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n653), .A2(KEYINPUT116), .A3(new_n845), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n659), .B1(new_n653), .B2(KEYINPUT54), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n851), .B1(new_n848), .B2(new_n849), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n854), .B(new_n661), .C1(KEYINPUT55), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n842), .B1(new_n856), .B2(new_n729), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n721), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n854), .A2(new_n661), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n855), .A2(KEYINPUT55), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n841), .A2(new_n569), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n720), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n702), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n643), .A2(new_n729), .A3(new_n644), .A4(new_n664), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT118), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n861), .A2(new_n720), .A3(new_n862), .ZN(new_n868));
  INV_X1    g667(.A(new_n851), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n850), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n852), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n660), .B1(new_n850), .B2(new_n853), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n570), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n720), .B1(new_n873), .B2(new_n842), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n607), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n865), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n867), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n698), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n671), .A2(new_n453), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n411), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G113gat), .B1(new_n881), .B2(new_n729), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n877), .A3(new_n758), .A4(new_n412), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT119), .Z(new_n884));
  NAND2_X1  g683(.A1(new_n570), .A2(new_n340), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G1340gat));
  OAI21_X1  g685(.A(G120gat), .B1(new_n881), .B2(new_n804), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n663), .A2(new_n338), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n884), .B2(new_n888), .ZN(G1341gat));
  OAI21_X1  g688(.A(G127gat), .B1(new_n881), .B2(new_n607), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n702), .A2(new_n353), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n883), .B2(new_n891), .ZN(G1342gat));
  OAI21_X1  g691(.A(G134gat), .B1(new_n881), .B2(new_n703), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n642), .A2(new_n351), .ZN(new_n894));
  OR3_X1    g693(.A1(new_n883), .A2(KEYINPUT56), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT56), .B1(new_n883), .B2(new_n894), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(G1343gat));
  NAND2_X1  g696(.A1(new_n695), .A2(new_n880), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n867), .A2(new_n830), .A3(new_n877), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT120), .B1(new_n859), .B2(new_n860), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n871), .A2(new_n903), .A3(new_n872), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n570), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n642), .B1(new_n905), .B2(new_n842), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n607), .B1(new_n906), .B2(new_n868), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n865), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(KEYINPUT57), .A3(new_n698), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n898), .B1(new_n901), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n570), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G141gat), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n743), .A2(new_n337), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n867), .A2(new_n877), .A3(new_n758), .A4(new_n913), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT121), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n671), .B1(new_n914), .B2(KEYINPUT121), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n915), .A2(new_n916), .A3(new_n292), .A4(new_n570), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n912), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NOR4_X1   g718(.A1(new_n914), .A2(G141gat), .A3(new_n729), .A4(new_n671), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n911), .B2(G141gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n919), .B1(new_n921), .B2(new_n918), .ZN(G1344gat));
  NAND4_X1  g721(.A1(new_n915), .A2(new_n916), .A3(new_n289), .A4(new_n663), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n289), .A2(KEYINPUT59), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AOI211_X1 g724(.A(KEYINPUT122), .B(new_n925), .C1(new_n910), .C2(new_n663), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n901), .A2(new_n909), .ZN(new_n928));
  INV_X1    g727(.A(new_n898), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n663), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n927), .B1(new_n930), .B2(new_n924), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT59), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n861), .A2(new_n642), .A3(new_n862), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n934), .B1(new_n906), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n729), .B1(new_n856), .B2(KEYINPUT120), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n938), .A2(new_n904), .B1(new_n663), .B2(new_n862), .ZN(new_n939));
  OAI211_X1 g738(.A(KEYINPUT123), .B(new_n935), .C1(new_n939), .C2(new_n642), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n940), .A3(new_n607), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n865), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT124), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n941), .A2(new_n944), .A3(new_n865), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n749), .A2(KEYINPUT57), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n899), .A2(KEYINPUT57), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n947), .A2(new_n663), .A3(new_n929), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n933), .B1(new_n949), .B2(G148gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n923), .B1(new_n932), .B2(new_n950), .ZN(G1345gat));
  NAND3_X1  g750(.A1(new_n915), .A2(new_n702), .A3(new_n916), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n607), .A2(new_n301), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT125), .ZN(new_n954));
  AOI22_X1  g753(.A1(new_n952), .A2(new_n301), .B1(new_n910), .B2(new_n954), .ZN(G1346gat));
  XNOR2_X1  g754(.A(KEYINPUT77), .B(G162gat), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n703), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n915), .A2(new_n916), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n910), .A2(KEYINPUT126), .A3(new_n720), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(new_n956), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT126), .B1(new_n910), .B2(new_n720), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G1347gat));
  NAND2_X1  g761(.A1(new_n671), .A2(new_n453), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(new_n687), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n879), .A2(new_n964), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n965), .A2(new_n221), .A3(new_n729), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n878), .A2(new_n758), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n687), .A2(new_n830), .A3(new_n286), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n570), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n966), .B1(new_n221), .B2(new_n969), .ZN(G1348gat));
  OAI21_X1  g769(.A(G176gat), .B1(new_n965), .B2(new_n804), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n967), .A2(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n663), .A2(new_n222), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT127), .ZN(G1349gat));
  OAI21_X1  g774(.A(G183gat), .B1(new_n965), .B2(new_n607), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n702), .A2(new_n235), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g778(.A1(new_n879), .A2(new_n642), .A3(new_n964), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n980), .A2(new_n981), .A3(G190gat), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n981), .B1(new_n980), .B2(G190gat), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n720), .A2(new_n232), .ZN(new_n985));
  OAI22_X1  g784(.A1(new_n983), .A2(new_n984), .B1(new_n972), .B2(new_n985), .ZN(G1351gat));
  AND2_X1   g785(.A1(new_n947), .A2(new_n948), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n743), .A2(new_n963), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(G197gat), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n729), .A2(new_n990), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n743), .A2(new_n337), .A3(new_n286), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n967), .A2(new_n570), .A3(new_n992), .ZN(new_n993));
  AOI22_X1  g792(.A1(new_n989), .A2(new_n991), .B1(new_n990), .B2(new_n993), .ZN(G1352gat));
  NAND3_X1  g793(.A1(new_n987), .A2(new_n727), .A3(new_n988), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(G204gat), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n967), .A2(new_n992), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n997), .A2(G204gat), .A3(new_n664), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n998), .B(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n996), .A2(new_n999), .ZN(G1353gat));
  OR3_X1    g799(.A1(new_n997), .A2(G211gat), .A3(new_n607), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n947), .A2(new_n702), .A3(new_n948), .A4(new_n988), .ZN(new_n1002));
  AND3_X1   g801(.A1(new_n1002), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1003));
  AOI21_X1  g802(.A(KEYINPUT63), .B1(new_n1002), .B2(G211gat), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(G1354gat));
  NAND3_X1  g804(.A1(new_n987), .A2(new_n642), .A3(new_n988), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(G218gat), .ZN(new_n1007));
  OR3_X1    g806(.A1(new_n997), .A2(G218gat), .A3(new_n721), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n1008), .ZN(G1355gat));
endmodule


