

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581;

  XOR2_X1 U325 ( .A(n330), .B(n416), .Z(n293) );
  XOR2_X1 U326 ( .A(KEYINPUT71), .B(G78GAT), .Z(n294) );
  XOR2_X1 U327 ( .A(G99GAT), .B(G71GAT), .Z(n295) );
  XOR2_X1 U328 ( .A(n368), .B(n367), .Z(n296) );
  NOR2_X1 U329 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U330 ( .A(n320), .B(n295), .ZN(n306) );
  XNOR2_X1 U331 ( .A(n458), .B(KEYINPUT26), .ZN(n567) );
  XOR2_X1 U332 ( .A(n571), .B(KEYINPUT41), .Z(n546) );
  XNOR2_X1 U333 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U334 ( .A(n309), .B(n308), .Z(n525) );
  XNOR2_X1 U335 ( .A(n470), .B(KEYINPUT38), .ZN(n494) );
  XNOR2_X1 U336 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U337 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n471) );
  XNOR2_X1 U338 ( .A(n451), .B(n450), .ZN(G1349GAT) );
  XNOR2_X1 U339 ( .A(n472), .B(n471), .ZN(G1328GAT) );
  XNOR2_X1 U340 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n297), .B(KEYINPUT17), .ZN(n298) );
  XOR2_X1 U342 ( .A(n298), .B(KEYINPUT19), .Z(n300) );
  XNOR2_X1 U343 ( .A(G190GAT), .B(G183GAT), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n400) );
  XOR2_X1 U345 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n302) );
  XNOR2_X1 U346 ( .A(G176GAT), .B(KEYINPUT82), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n400), .B(n303), .ZN(n309) );
  XOR2_X1 U349 ( .A(G134GAT), .B(G43GAT), .Z(n330) );
  XNOR2_X1 U350 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n304), .B(G120GAT), .ZN(n416) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n293), .B(n305), .ZN(n307) );
  XOR2_X1 U354 ( .A(G127GAT), .B(G15GAT), .Z(n320) );
  XOR2_X1 U355 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n311) );
  XNOR2_X1 U356 ( .A(G1GAT), .B(G64GAT), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U358 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n313) );
  XNOR2_X1 U359 ( .A(KEYINPUT79), .B(KEYINPUT12), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n326) );
  XNOR2_X1 U362 ( .A(G57GAT), .B(G71GAT), .ZN(n316) );
  XNOR2_X1 U363 ( .A(n316), .B(KEYINPUT13), .ZN(n365) );
  XOR2_X1 U364 ( .A(n365), .B(KEYINPUT15), .Z(n318) );
  NAND2_X1 U365 ( .A1(G231GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U367 ( .A(G155GAT), .B(G22GAT), .Z(n435) );
  XNOR2_X1 U368 ( .A(n319), .B(n435), .ZN(n324) );
  XOR2_X1 U369 ( .A(G183GAT), .B(G78GAT), .Z(n322) );
  XOR2_X1 U370 ( .A(G211GAT), .B(G8GAT), .Z(n396) );
  XNOR2_X1 U371 ( .A(n320), .B(n396), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n574) );
  XOR2_X1 U375 ( .A(n574), .B(KEYINPUT114), .Z(n558) );
  XOR2_X1 U376 ( .A(G92GAT), .B(G99GAT), .Z(n328) );
  XNOR2_X1 U377 ( .A(G85GAT), .B(KEYINPUT72), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n372) );
  XOR2_X1 U379 ( .A(G29GAT), .B(KEYINPUT8), .Z(n329) );
  XOR2_X1 U380 ( .A(KEYINPUT7), .B(n329), .Z(n344) );
  XOR2_X1 U381 ( .A(n372), .B(n344), .Z(n343) );
  XOR2_X1 U382 ( .A(G218GAT), .B(G36GAT), .Z(n388) );
  XOR2_X1 U383 ( .A(n330), .B(n388), .Z(n332) );
  NAND2_X1 U384 ( .A1(G232GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U386 ( .A(G162GAT), .B(G50GAT), .Z(n443) );
  XOR2_X1 U387 ( .A(n333), .B(n443), .Z(n341) );
  XOR2_X1 U388 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n335) );
  XNOR2_X1 U389 ( .A(KEYINPUT65), .B(KEYINPUT76), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U391 ( .A(G106GAT), .B(G190GAT), .Z(n337) );
  XNOR2_X1 U392 ( .A(KEYINPUT9), .B(KEYINPUT64), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U396 ( .A(n343), .B(n342), .Z(n473) );
  INV_X1 U397 ( .A(n473), .ZN(n561) );
  XOR2_X1 U398 ( .A(G36GAT), .B(G43GAT), .Z(n346) );
  XNOR2_X1 U399 ( .A(n344), .B(G50GAT), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U401 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n348) );
  NAND2_X1 U402 ( .A1(G229GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U404 ( .A(n350), .B(n349), .Z(n352) );
  XNOR2_X1 U405 ( .A(G141GAT), .B(KEYINPUT29), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n360) );
  XOR2_X1 U407 ( .A(G197GAT), .B(G169GAT), .Z(n354) );
  XNOR2_X1 U408 ( .A(G22GAT), .B(G15GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U410 ( .A(KEYINPUT66), .B(G8GAT), .Z(n356) );
  XNOR2_X1 U411 ( .A(G113GAT), .B(G1GAT), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U413 ( .A(n358), .B(n357), .Z(n359) );
  XOR2_X1 U414 ( .A(n360), .B(n359), .Z(n543) );
  INV_X1 U415 ( .A(n543), .ZN(n568) );
  XOR2_X1 U416 ( .A(KEYINPUT70), .B(KEYINPUT74), .Z(n362) );
  XNOR2_X1 U417 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n376) );
  XOR2_X1 U419 ( .A(KEYINPUT73), .B(G176GAT), .Z(n364) );
  XNOR2_X1 U420 ( .A(G64GAT), .B(G204GAT), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n389) );
  XNOR2_X1 U422 ( .A(n365), .B(n389), .ZN(n370) );
  XNOR2_X1 U423 ( .A(G148GAT), .B(G106GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n294), .B(n366), .ZN(n430) );
  XOR2_X1 U425 ( .A(KEYINPUT68), .B(G120GAT), .Z(n368) );
  NAND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n430), .B(n296), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U429 ( .A(n371), .B(KEYINPUT31), .Z(n374) );
  XNOR2_X1 U430 ( .A(n372), .B(KEYINPUT69), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n571) );
  NAND2_X1 U433 ( .A1(n568), .A2(n546), .ZN(n377) );
  XOR2_X1 U434 ( .A(KEYINPUT46), .B(n377), .Z(n378) );
  NOR2_X1 U435 ( .A1(n561), .A2(n378), .ZN(n379) );
  NAND2_X1 U436 ( .A1(n558), .A2(n379), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n380), .B(KEYINPUT47), .ZN(n386) );
  XOR2_X1 U438 ( .A(KEYINPUT36), .B(n473), .Z(n577) );
  NAND2_X1 U439 ( .A1(n574), .A2(n577), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n381), .B(KEYINPUT115), .ZN(n382) );
  XNOR2_X1 U441 ( .A(KEYINPUT45), .B(n382), .ZN(n383) );
  INV_X1 U442 ( .A(n571), .ZN(n452) );
  NAND2_X1 U443 ( .A1(n383), .A2(n452), .ZN(n384) );
  NOR2_X1 U444 ( .A1(n568), .A2(n384), .ZN(n385) );
  NOR2_X1 U445 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U446 ( .A(KEYINPUT48), .B(n387), .ZN(n540) );
  XOR2_X1 U447 ( .A(n389), .B(n388), .Z(n391) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U450 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n393) );
  XNOR2_X1 U451 ( .A(G92GAT), .B(KEYINPUT93), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U453 ( .A(n395), .B(n394), .Z(n398) );
  XOR2_X1 U454 ( .A(KEYINPUT21), .B(G197GAT), .Z(n434) );
  XNOR2_X1 U455 ( .A(n396), .B(n434), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n516) );
  NOR2_X1 U458 ( .A1(n540), .A2(n516), .ZN(n403) );
  XOR2_X1 U459 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n401) );
  XNOR2_X1 U460 ( .A(KEYINPUT121), .B(n401), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n426) );
  XOR2_X1 U462 ( .A(G141GAT), .B(KEYINPUT86), .Z(n405) );
  XNOR2_X1 U463 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n431) );
  XOR2_X1 U465 ( .A(n431), .B(KEYINPUT91), .Z(n407) );
  NAND2_X1 U466 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U468 ( .A(G1GAT), .B(G57GAT), .Z(n409) );
  XNOR2_X1 U469 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U472 ( .A(KEYINPUT1), .B(G127GAT), .Z(n413) );
  XNOR2_X1 U473 ( .A(G155GAT), .B(G148GAT), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n420) );
  XOR2_X1 U476 ( .A(G134GAT), .B(G162GAT), .Z(n418) );
  XNOR2_X1 U477 ( .A(G85GAT), .B(n416), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U479 ( .A(n420), .B(n419), .Z(n425) );
  XOR2_X1 U480 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n422) );
  XNOR2_X1 U481 ( .A(KEYINPUT92), .B(KEYINPUT5), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U483 ( .A(G29GAT), .B(n423), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n514) );
  NAND2_X1 U485 ( .A1(n426), .A2(n514), .ZN(n566) );
  XOR2_X1 U486 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n428) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U489 ( .A(n429), .B(KEYINPUT24), .Z(n433) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n439) );
  XOR2_X1 U492 ( .A(G204GAT), .B(n434), .Z(n437) );
  XNOR2_X1 U493 ( .A(G218GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U495 ( .A(n439), .B(n438), .Z(n445) );
  XOR2_X1 U496 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n441) );
  XNOR2_X1 U497 ( .A(G211GAT), .B(KEYINPUT85), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U500 ( .A(n445), .B(n444), .Z(n457) );
  NOR2_X1 U501 ( .A1(n566), .A2(n457), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n446), .B(KEYINPUT55), .ZN(n447) );
  NOR2_X1 U503 ( .A1(n525), .A2(n447), .ZN(n560) );
  XOR2_X1 U504 ( .A(KEYINPUT107), .B(n546), .Z(n530) );
  NAND2_X1 U505 ( .A1(n560), .A2(n530), .ZN(n451) );
  XOR2_X1 U506 ( .A(G176GAT), .B(KEYINPUT123), .Z(n449) );
  XOR2_X1 U507 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n448) );
  NAND2_X1 U508 ( .A1(n568), .A2(n452), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n453), .B(KEYINPUT75), .ZN(n478) );
  XNOR2_X1 U510 ( .A(KEYINPUT27), .B(n516), .ZN(n459) );
  NOR2_X1 U511 ( .A1(n514), .A2(n459), .ZN(n542) );
  XOR2_X1 U512 ( .A(n457), .B(KEYINPUT28), .Z(n521) );
  NAND2_X1 U513 ( .A1(n542), .A2(n521), .ZN(n524) );
  XOR2_X1 U514 ( .A(KEYINPUT84), .B(n525), .Z(n454) );
  NOR2_X1 U515 ( .A1(n524), .A2(n454), .ZN(n467) );
  NOR2_X1 U516 ( .A1(n516), .A2(n525), .ZN(n455) );
  NOR2_X1 U517 ( .A1(n457), .A2(n455), .ZN(n456) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(n456), .Z(n462) );
  NAND2_X1 U519 ( .A1(n525), .A2(n457), .ZN(n458) );
  NOR2_X1 U520 ( .A1(n459), .A2(n567), .ZN(n460) );
  XNOR2_X1 U521 ( .A(KEYINPUT96), .B(n460), .ZN(n461) );
  XNOR2_X1 U522 ( .A(KEYINPUT97), .B(n463), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n464), .A2(n514), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT98), .B(n465), .Z(n466) );
  NOR2_X2 U525 ( .A1(n467), .A2(n466), .ZN(n477) );
  NOR2_X1 U526 ( .A1(n574), .A2(n477), .ZN(n468) );
  NAND2_X1 U527 ( .A1(n577), .A2(n468), .ZN(n469) );
  XNOR2_X1 U528 ( .A(KEYINPUT37), .B(n469), .ZN(n513) );
  NAND2_X1 U529 ( .A1(n478), .A2(n513), .ZN(n470) );
  NOR2_X1 U530 ( .A1(n494), .A2(n514), .ZN(n472) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n475) );
  NAND2_X1 U532 ( .A1(n574), .A2(n473), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n475), .B(n474), .ZN(n476) );
  NOR2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n501) );
  NAND2_X1 U535 ( .A1(n478), .A2(n501), .ZN(n488) );
  NOR2_X1 U536 ( .A1(n514), .A2(n488), .ZN(n480) );
  XNOR2_X1 U537 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NOR2_X1 U540 ( .A1(n516), .A2(n488), .ZN(n483) );
  XNOR2_X1 U541 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n484), .ZN(G1325GAT) );
  NOR2_X1 U544 ( .A1(n525), .A2(n488), .ZN(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n521), .A2(n488), .ZN(n489) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n489), .Z(G1327GAT) );
  NOR2_X1 U550 ( .A1(n494), .A2(n516), .ZN(n490) );
  XOR2_X1 U551 ( .A(G36GAT), .B(n490), .Z(G1329GAT) );
  NOR2_X1 U552 ( .A1(n494), .A2(n525), .ZN(n492) );
  XNOR2_X1 U553 ( .A(KEYINPUT103), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  NOR2_X1 U556 ( .A1(n494), .A2(n521), .ZN(n496) );
  XNOR2_X1 U557 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(n497), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n499) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT109), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(n503) );
  NAND2_X1 U563 ( .A1(n530), .A2(n543), .ZN(n500) );
  XOR2_X1 U564 ( .A(KEYINPUT108), .B(n500), .Z(n512) );
  NAND2_X1 U565 ( .A1(n501), .A2(n512), .ZN(n508) );
  NOR2_X1 U566 ( .A1(n514), .A2(n508), .ZN(n502) );
  XOR2_X1 U567 ( .A(n503), .B(n502), .Z(G1332GAT) );
  NOR2_X1 U568 ( .A1(n516), .A2(n508), .ZN(n505) );
  XNOR2_X1 U569 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  NOR2_X1 U572 ( .A1(n525), .A2(n508), .ZN(n507) );
  XOR2_X1 U573 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U574 ( .A1(n521), .A2(n508), .ZN(n510) );
  XNOR2_X1 U575 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n520) );
  NOR2_X1 U579 ( .A1(n514), .A2(n520), .ZN(n515) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n515), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n516), .A2(n520), .ZN(n518) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(KEYINPUT113), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(G1337GAT) );
  NOR2_X1 U584 ( .A1(n525), .A2(n520), .ZN(n519) );
  XOR2_X1 U585 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U587 ( .A(KEYINPUT44), .B(n522), .Z(n523) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n540), .ZN(n527) );
  INV_X1 U590 ( .A(n525), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(KEYINPUT116), .B(n528), .ZN(n533) );
  INV_X1 U593 ( .A(n533), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n536), .A2(n568), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n529), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U597 ( .A1(n536), .A2(n530), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U599 ( .A1(n558), .A2(n533), .ZN(n534) );
  XOR2_X1 U600 ( .A(KEYINPUT50), .B(n534), .Z(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U603 ( .A1(n536), .A2(n561), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U605 ( .A(G134GAT), .B(n539), .Z(G1343GAT) );
  NOR2_X1 U606 ( .A1(n567), .A2(n540), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n545) );
  NOR2_X1 U608 ( .A1(n543), .A2(n545), .ZN(n544) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  INV_X1 U611 ( .A(n545), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n553), .A2(n546), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n551) );
  NAND2_X1 U616 ( .A1(n553), .A2(n574), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G155GAT), .B(n552), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n561), .A2(n553), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n560), .A2(n568), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1348GAT) );
  INV_X1 U624 ( .A(n560), .ZN(n557) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(G183GAT), .B(n559), .Z(G1350GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(KEYINPUT124), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(n565), .Z(n570) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n578), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n578), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  XOR2_X1 U639 ( .A(G211GAT), .B(KEYINPUT125), .Z(n576) );
  NAND2_X1 U640 ( .A1(n578), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n580) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(G218GAT), .B(n581), .Z(G1355GAT) );
endmodule

